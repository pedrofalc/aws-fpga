`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YTVtN8QzWrYo1pFic/+Vul/WDqHelcX0ZKT5/4lDCe2h2pgu7WYqQ/lLOn9ykjcjgnJxfJGEPGpD
4edBRY29lA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eT9cdJs2jqwCov5MlLAVKkPTG1C/9KSX5UzxnfKuzHlqHICvdjqXrS56PTsCS3/OC0qpzmXmBIdI
5jXm6fWEYxndn4CvUXMAbZEvA4GVVifRiH1SkIqHaQGNseSc2Zw7znLTTO/vE6NZUQdfCqW68aLq
J3kIDJrB1WhdAW1AGEg=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
W2kLRKgikIYVbrbCUEOzZvj9sVTYc1XSCe2parkGOwIgZ/XryQvhmOLw9g47hOTmWd3I5J+vR6ff
N0SNxYHQNHTkdoqezxK5LlPCic5FrMwYwt3VA01kcjl95Hx2ywhuBQI7E+KHNmStIar5S1ZN/YIw
+tG3rjDnA+/uZo4r6MA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Pmt19WIAgtDUaBtpZNbJ7Lc1cxIhTjSp7+5D/N0tPhD6lSzmdzysgT+lKRPHLJBF3yupfRCu51Qe
3nR2Vxh75X5E50u15G6wUt9kQRGDuEPqL5oZwHBQZwiPDBh8sXONq5/zFHoJDpZylei2W7799CAP
whzsEFOuFxrdsds5DLuJ9f6DchdvGFoWhYjqEBLZZDFk3B1uQlaUaxYfL6hteOazoMHo9GuoB4xv
Z6VlTWdTmNdZmwbpxq0gWLWLaYvT+8lGBQJhRVLQwdVrNvieu7rW4zWvjyUcciLWwru8MbHzIEWz
iTdP6gJ1GQxM88v5Bz2ONgCqPWrKeSDknD0eAQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lIVh6WmUy/h9dIJL0bvhl87k7DaepshSP3bmQqWkcFvcKHa/1g1QiRA3e/hJsjjFQDn34pUe18x9
9m4V+k3kXtWkbbBszSjZ7SGcID4W9ikrmU+k1gGPlj/qmJ3uuN2+OWrsoqvRV3q49oOQ1t/gRZU/
yEqakLPUgTI+d2M0n4EeP+Ixkt55I576X9c9qjSOQVD7izTIHNSy7Ri7n7Aa2tFDVtHKujjZC0Rb
jy4zLGT8F8HCh+53/a5pE3pwhTcFQF5BWBzJkjhZ8EdcoOaCeimQFf3OVGJxKL+fmqHS8bVEJJwb
9uUcPm5ePAhDnDL85QhG48H6VoKv1wRaOGyftw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uVZP3fyoZWBGatgWLoQczDDlpyZf4yBvWNMZt0AryzY0se/585MwXMFzjglNp+BtbxwWMh3Gx3ze
MNcyo/doyzkkWE4Okk/uGSkOT2VGD5sgbnKLLqA8gGl9VFGgJnIa1YoVTHhEDRBjC2iGbL03bP9Z
HplCesExbsG7azRdHusKPaFBO60RtnkmVYx08xFTr+BgIcMBB0CjVHQ5IBNLZtb06ydf6R3MkE8z
pde2MOQ3qMl6Awo8aSNNEVujzrztyEzMT2acmi0v25iIsrZnjuHsmh+NcPTLaYW/foK9FGTQi3ZI
9+HAdzZmF7zpx5hU0EJ9Lf4tX2SfyDag5+APaQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432720)
`protect data_block
6t7yCo7+UAw1mvOoB0HH3wc3Hz2W6jELu51z4lPuYMggsPGDhiE+LynddfUyIbI3zCmzyyem0jJo
lAgi9M7PwLKhmEXPPNs8/0RIQqLUAx7qpnmwWsO5jIKvmbRTgolTjaYgMT+m5EIeWDPMIB8QlvqA
s40Um5eHkKZeZ3HLVhgDnYi05OMLl1B6Kp5p3fard8vk3Ilk+n8GAOmErLct88wzGNqhlfuXQ0xX
0IJOxtf6DsnOi0Q/KzwilB5cgPNSJcnBIBnbq7EC5V2dEWqSa8/gIIgpu9OrxNaKGrpF6Ca1O4ER
hvlT9FsuAjDHxaHSLtTm6Lv4ARHcpodeey+tZqXLMX5kIN8D0hAKcKM5fucG3ERfHnOEXODgU6Fw
ddyByxs1cLbvL/AXWvkfGzV/IpwhOKb4BtMsQGn7LmKRHHU/YzbKf432Q3IKWqxtRqbMPGNEUSZh
JOKdPo9vxiQEHlmK4YKGlKo8hpJbH0pLEIXmMESO4FT5kcdtKB65Xgv/aoSterOz39RLgbgDdDOQ
CNg57b1ZhDc+mgNTOLUgP9Nii8ij6nDoZjSSfu0KktY/jdbi2y2Wp5DJxNZqJ5yALtCpKU0NlrFU
sThhEomszFJGBeTn6S0FW9GN0/HBZGj+moR1aCCVC/0TRARosSK1FglByNpoa4lCgZwX4EiIuxL1
4nKrWA2GIbax9byMAq2y0ozkwQ+pZ28Ofwex7u1Dpis9s0O/5xym3pzCvala+mScLlqKOgMJ01yT
TSmCkdO2t3WIKY/oibUUFxy1Aj2i+jwdD4PYqEFH2Z7hxsDebM5SgpOBlqXNqPzCEQX/0d/PYVTQ
kFHIaiIdIN/289EzPWopC5ywuWQy8H05Tctx8oWP42Bj0CaZGiDoxQiFDZTmMkW5NEpdhzQElxRT
1mDZQgZZFaNrn9OxwwNisHpUR051/GeWh+XFJkV5dUGgtkKs6FSswpnA11oJkD1rZgXT9x23cdLt
/HDs5qRvSC9AfOdWJAHWuk5iJG2nIf7qhSsDJmAcX8L6pgKaLETaUJVi9erfCNLzMowtBr9hXUer
xhAd+YiurimfEvuz9xdZPuoJ1k8alyCKQxCjqhBIcEZMd5/upDcIuzv5yrjis1pwbRVG4r3rNFnG
C+/xHkMXmOOJPrWeiLx9SE+TPVs6+ASbhtZ5BoBHGfA3qANgS073hDszeHDxxDuJ7zfQ/bGqIkku
933d1cdrMmaDrwu+u5BkrtHz2mLqU8eBE/EOUgy7wE7Y1AhS9e/hCD+eYHmx0b+ATxhKbSWJWrIs
uYdyfV3kVJbPjPQmY1DvysVBMm3fU7WduHl9/85uRUpYZOvOhI5EcdbavdcDaq9YGqN2axyVYUbU
ZyLSlSVKlUjQQ5uEYV0ds2IgS+exU675Jw/rtd/W6Z9caxjvp6aLHoNYdl2mzISmpvPu4rVUmmJU
13xEru2PlWf032/XFLRhmykPByWauci6ZfeKKlIGup10EqjtTBo5SFbGlF0ZcYVUDzFG/7NUPf9J
ZbkbzVdNQWRTh2W0s5H8YLAikrlO+f2ch9cPOYsmHaiD9pbjY8qcf/+SVee5Bx7+Re3KXYLbHhyx
3um9F7uhFVva+iZnpypI1SjiVK7mR+UmcZmz7bZHIHHqf+AFhtBD9Tm5YZR3TrGnPh5Uvn7g4RuY
xrnL484CefKQ8LUkLiY/gLc7KYg+7RbBuOB1+T6HFnnTzYDCqbf4OoYb/jIAc0Tuj8oIKa3s7hrT
KmXrPTPIsNmfe3SsWLxydv81RR6nH8Yw6j2/muwcJRB4d2RLIUGZnNzzxkydrASFCZxCF8gCn6Ib
QiODwKzafeoYg9l8lRrYEHRyVrlCbyd7pAYNFSS2zPFCqTbbODhHMxF7kn1S1lLEJ3eAU7msSZUA
FnmwGvsbNipDPiI5OUASjvl7ynXFnzEJhb7j0lrVV4gV70na7Fz0OV3s9DOxWx8xiJKBLF3hz2P6
ybnHRvU0K9B0tBuDxyW3RdOQXd00O6zwp6xO+nOOWhvfr/XJ1NEZwW5pPGW4YvdHj7yaTGNR1bwc
TrWok5JJupQxJ19VNZqjJHLCmd/uf0PdJx/QDJcSuwTRh0079DIMeuozMxCoGy5uzs3eG6efkbuU
CdXvhKJq8/t1TQ0p1vwzRoZQkGrTlaBrfYpJj5EXRk9MUtqQ+Xg2r2t2zkQUJaPt9eKB8XTvUroO
SVHHrB8r9mXE+HYmR+kAn7N5nl7/Znry0+rZKuJklaO3mMarx441Jb/6Q0RAIFASz3RCQISFWA1f
K7E9iF2yPdPSITJQRvBbWwOEm/3+CBkhvW6XOeQdbqLTk6bjjK03pXnocq2pM2CIo+53hoYGUyBN
WgoqYNZdjOJiMAQsDnUTvo/LHblYSiNDPskr4+9M3UPDcnH2OTZKiA/diyQzCgtHN1WtBs91fpYw
4k2tjkG6U0XXjhgSkXJUbc2Dg1vDQtwOiUpY2WQRJUvjhBxHnoxGKidr8mDMFichY6eQo4EoUnn/
WV41wxABASYNxykoLoLq9T9Mdtewp8h9gmicmHzA+UjWU1xC5cO75412kTa8usftCd/nbLzqzaIC
JlrbmJacQI/6Ts++RMw1Ek0I/y4Fx8a7ej9DsVNUyGzK0Jc55JxQFULjH40Hwg3k7umN/JUnW5nL
XGVdCrrKFDujXbvqOotfujEhFAHTr9NrDFVhkbZ1TtNBXjT6wpa5LZqWG7BkzQe3+u23KRfxI07z
Frj585ztBe4dDjhk7p7moc98TX2LKQUm977AoXRNF6RAc1INcn36FZbbT1S0N4lo2tTr9kU+fxbd
XgJeZSKhz6GsAat4kFhoSBqsRTLQjaxZoNBi4kGZEO6w9IU6fBbCvtBmWorxBX+7RqaCZajiJEK3
aVERGjj19jw9jzjlKyRTFC1ymsRLpOda3TZPXR1rPDE3K5mgy5DLaqtXqww/h0cBnFR2dIBHt+DQ
C12sF5D4pwetYMDL/s7NFVNBKIafD3taVTKyi4pbZirzLiSMQ5qSp3R3wADQnJE9W3CYcKCURqph
qboLD/nHfnTHy7t47kklU3kf6IbwOM8BYug9B6S16ykNZNNUQFNKumA/kxms6Mao2iimbk14Qoyw
G0peQsc2Mf/G8ZMpebugyZ3cO+tB8e3qEOrLYdXspK0vRLOIdzxhk9m9mPNZGveL31TBb5ndisgT
1z9RlV9XM8TNSZ7SXL99W8OaXX8aOrT2cIfrZEJguZ7UeGTCTZaCyyN3V8zLrGtoG+B25uYCiE3S
tCGcle0EgsCGPeshPrlZlxK11c23zQ0N9A9bjWt73uoXkvchv8NIzQa2xsV78a0NvNg1iDKcJ6H1
aaNrCYK3FwxAAbf6EVuLrOW4Obq3iZ4fb8BYs3lajGpeJmKYtedFlex1zEOzfMP0WKBImPxjdAof
Fzpf/b6go9bFgGM14aBwX0UNU5/FxiJ105XpaUjnezBR2BxYQ7SY1CRG8RFw2CVMxFtljctWC2ss
qm/zVuWqPpHS06nZ1HXPdT6FbWSUCnXtCrzh6jXxyOVLiXgG/FXcCBN7jmHSHBnDDQ2HJJBlXTsQ
ym9t9ozKasDhsS95cYlNtDJ1ZXAd/d57fNzeGcD3P+Y1qi+KcKqGsXSUPJpEq0Vl0rgJTMaGyygz
71YiK4xZb7Ak+5cswDLQk3sajowS+LnaUwzhWld/r1uRuUJYBGxbvLtp+hUXw+qSyA1As6cCL4za
7/YDVIfO7y/oIf4tvADu2CWTNgbujmtY/X/FaL9FTkBYt4VoelOfZrdKCvk8YlnycYhXeTWenSnu
I0nGmMkb6gH+6WIwaay8ncOoWLOP/e5RnpU7x27XoyfE6B6Cwvp9Yp+jk0BelfVG32dX+T9VEsaj
OlyGbuj5X0KxOqjfdspptWW4PAw7DUSyAZZbcSXcaUxo1zGhljuuE8kgEIOUWSsELFFbnp9z4Bw/
v/vgOsPD7S3E+iOx3LZnBrPKpS0SyUWrrgO7a2Oo3SzKBrpR4a7cPiZqZWMFpnh0BsVm3LVEkzva
PGs2t2uAf7ZlTA8okFSw8d8QCkvSNgKJYMu8ODgZ+bahDZp8L96NH8huKRFsPaOtIegYSpW654eP
waidxqLhvrjfUpufyxosOP408tKguALccADuR/w/z+48VUy9pe4j1/2QLryuV/fDB/qk5yoVg3Mm
OMyFY/Eu3q4fwEGSMegebS9uPAa+Z/0ao6HYyMYWBd7chOFDIgcUjwDGEaiXmSK1byskkb7Ln4j/
aYm0yhBrfAmIC2VnY9K/0p8yPyqrMoS/V/pk6Nwl84lkDcZhkyvlrK+TRkNexrsxPs/JhqY4kuj8
yN7pVpZlkM9HBdKpyCPJmu1tk0KGl9dOeWYUdQo0qYXA2yfbexCj4CjPGPMc4UU21pwXBE9hAMN6
uVRAkkPhLhTqGYTXlKFgQkSxq6zwcyWFQBgYTmy/NRA6F0GAS+/ji7LYmx5Ll2+kKKdJ0u7xIwfP
JqsCpeNrT8/o1RsL/QSqoZ1mCnhLzABciCr9X+UWXRfnqGXuh+4Mdhy7Prrli7puWDr7uTkxhFGl
rn/NlgHdw++LZ6+pwh08G5jkMwBYW7NEaEntgUtrEFApPSTjBzPlXBKVxXfGxbap90dS2ON6xdAo
HMbpThkcVTypwu1XIU9/j5IhuNqig6NV5tNKOyQ9dXAyjJ89+gHhy8HfZXouQ++P4quJtqJozQPs
3pXWwS1U7PXkJKtN66805BpjwPXuztNexvTYDPBUBAtAFX9pOZjbXbCLqxN7hKNKZdRUJr01Vu8n
cMVF92FbsvnSvr7X4ahatZaF/C74ndLyIWo06/PKg08ytgmhfe5fBxdW2zooT4+RqMMbIOfKduR8
jXQgjDD/wuVm5Zg1dch1wlc35ie3+gKe+lymYjfiEwtUKnu2xdLjFh07WPLyKqfgRW3kdCz2IdVi
Vei8BxTgkAgBouUADUQT4wOJmU0NJpw/9fGaLFa5+0a8HgY3vGRPaP89+VrJGUZLODhjzmVYsHOi
RJ5amuHK9mODDrXBmfmrp3EBuxj8IoFeLiomTLUoE+VEMS8IXxPEDLIEDk0pUzrVrI9ra6T2sJU2
q2ORksMUHilrauoxqGOadg3T8NN6Zz7dv8SQVZeKh8YEoTnjznXUpGK2KmwGtGV/5WBc0RTChIFm
Onz3T2PUcJD4Fhh3uIGqFjtRwTFs7WLqrjSi3gqHqsU/JUBas1o/nihKbrmNVQRLwhHi0PfziEu9
pB4OssbAwTvxA+WYmgTn+LhybE7ncjVEU+spDVYUXN5S0wtYiVPHK9hOnsX/yoZ3CrQeR14AraOs
7qYCEwQ2AqvROsBuxp0WkAtLJDHyVWULgh2IWEB+NB4aeN8F1FbctML7MPI/E03R1/y+7BMZfi1+
A+rcgLIKBp91gtMFeDqbaBpQJsvq5+zBFj2cW+Y9HOhjkNgC3CzpdhsJDOPg793DZs0qTAIyBy6u
vZh7UeaJs6eBgZiNhSFUoLIugn3weHuajc5NRERzLidUiOKA2upjGA9k9MDZ4lNfaa/D1uY4z+et
0iY7btWiEGICNqQ5WXWk0VBmfSRGoEz8C0+xTAU4PuoqIrACtMMyenVAwoefuE7eiEb98rqkDGEd
9qgtMoRlcDajdrx5R92HM/umWIfukGRaGqjE4u1FAyb32FHzDMlJTERT4WzWA6dNxt6Iw9hE4HA1
fG6q1gQ/lz3N3JxGnTcMsnZL28FH1rYqZSiRRcFCCyGOX/VOwd7Fb/0VOgNQhNchN9oV3rluI8nS
0IbLB3Ox5vj+/D9OavOPjFm/H6T+mac/la5hVgnv7moAdmNYGEPoKH02C6ffYsEsRajGUInhNCMS
+gSl/kzmmBwPxKxpmP9uXvov6RLXc8Rl1HW87tqK1rKK8yQ8P8X8lWFYt98hzr3Ci2Fm8rNJzLKd
zT543XjOgnW27yxnPXuUYGpZHO8wIkigthGWuaENndXiaB53rQryAeT3noYOOqTipsF7909kN2YQ
NmCZmOg61dbuFibjng3Aou4Lfc26HdJqRZl1IAtXBH8U14IJdMY8GkzoMfLe5JT53HZxIK0hMFAf
+CfjqG1zWpsS0s4al5fRIOxrQGjxscH0aQnzZaoj7aqEtSuIDTg+3G7Rhoby0h0gucygon9GiTSk
8rd231LvXKPDt9XDxPqb99PCra1+ldewGvk5jACJp/zlKWvfzK7M65611rqdkZJhp6bmPyV+yh78
cH/RvtnbMGEgQA5T5jdJKxxe6pL1FRLSkC+czwXsfHGF1LuINVavC7tfZ9wo8dQ/qD7ZQN7lEBCk
DVSUydrHsFVY2EmTjsu6FiJ3en/ku5PlKt9pjfto6ReRiUpYXDL9yOuFqlwzq1LevStBpGsyWlsf
To2JgZu0PmbHAEScFFHz45oB9ra38MlyI/RSNP/lpRSazmLfY7J9Bi7Z3yUzZBB09JfQBH7qDxN4
dGt8jNaJfKToC2Zsj9J3NfHHcQ7RwTbOmmR5ffe7X9zbERR7aPQ/Kzq/SoFz+OtIQqQySds9IRDX
H/yPWvZcUNpw+X0gFvB12q+RQEBLQmSR2v87ZFR5Fd54Z+ACMg1pjwFIB0V4IznvGIpFk/MvWgpX
gjtrqiNDCoTWiQGn566qec8PSF+0YT8N9bBfy7O4qEEFjfe1mgokfvBcglknl2A7nyYbBXbq4kEP
+iJYZE9h+pQkyYJdENRAn4wHe9KNloAkFIpC8cLkkCMZh81gb5UQLtc/tkJ/8CTTumEtjp3qz/jb
a0jiy1OMMj2T4fbWBTle2NEuS6kcGa7WVLb9HSbdolhiB/ZYZ/+dWM3x4+TnLCKbz2OMCTySAGb4
SdX4u1S1AZTP8Z8zcdxAGIj9WqMMOypOBvolAxmrKrPYKvTctVJ7P/WgO3R4V7eMJ0mSZuMSZ4XR
Z3olkl4BnVS3eE8zGoBm0DSlqBPTO27qutZdTBwZ4V0yDHHu3eiHSZEjKfjcJdc8E3pfr9eaUqIO
0YNO5wn3/ICT9J21u3tG1814BCCyENsVcmciMXv/hgS+8o42Cdp013NKru/AVZkUeboqx5nV3m7Q
t8Oq7jpHvE+msqoPk3BKVeLi9fyxKA3MEpmhSibqkDXk3dPTBJZoo/JIQ2dyzNQ/Ab/qNnGIhWUo
gbTqaILP2nuLYfSJX9O9tPDCDhadJmV2dc/tpjr9rVKm4pdTK7OJj1mRLRb3sDhlpsXZcfpSS1xr
eFJEXGAXg1xqY4GWcKvfrUmKICCBnssFHCrH3lK18A1IHDSeG1A8ROc4lor508OF5fkRObok/3Ph
4+wI0oFcZZxG9l5VPzp7xXIFZaXt+U4/BaCCPMNO2+oYJOqAnUfWVPaG3JZbd7NsSFdC/n7xx/S1
Z9mH0Bi1OsvK8dHwx66064DGiilO8PUtL8HiOQtz2H3Izm4BjU2RGfRdq783TxKkbWH+q7ntLaTY
I+LxR79rEae7DRHsXHCQbLpwhXbDIHNVfNMLEDikwJ33m8a2A+9idv2BhFXG3ha4JXIldO9hYvAm
NYOkNWGHPIYXaRz747qf8tgq3LMxpy51BFy+iFfir9zspjBFQwL5qoGTZCziZFrJbE4D+WzoRXc0
OAz+Y1rAjq0dt59gqJuPrLZa+AIaH5ZluWdiczmzPcAP9WShoruYUQOhsrb6m5Plt+mw3XV7yRJy
fPCQh5O+CiPq7bLuSfcNqtg0vcJcfX+eh0BSrYrQ4Zo87hoBRbapJJMfV5FybMwuhTIoksNUL97Q
ObsHsj1m9lFCxPGyWD4dgP5rcrYxGp3LiBaEws8I/xubYxsix8geWNtKjXtfNQ1+u2hyZC5GeyqE
TD6VQLa8828E3VQaFg5nZ8AUyf/0i2kpPm28bKcMt/n9p39HDHADvczz0XUg22dxmIZB2WvXCkDu
gJtCCE+l4yxMGQc5lEx7V2HBujCbJzOkofWfCn+HQ2oHFkjJ9DFQsQ34Hn+6dRpuTCzFA66Uy56Y
aZsDBK+2g4Tmzx8B7kLeXeH5SQTP3pJXY4axPOmgAjHnM5do2xFpOP07T7C9JCaOi4nWM9qrqSH3
NWApcQo54K1ZO9rx8vdRz0GaGVrU6wGJwi+TJTfqQj3Thr/92LsM81kwRKonMpacYe8bI9e8ZSXr
wamdj2asL8UzrcYyP5KiC4Di333ARb6gc86/6V1Oo13G36poVpaayTK3+cIB6f16E4j8gOZEhxnm
gR5m0jsD05qbroq3ZCzcixkIM6pEeYsGXTDSUXjzxqo8RWUoO+01CtMHs665r1Xf8KXgUxV9lTdX
VuKNkZS2+K7IVUJ6yijfRyi5CuKSEvutxPhx38wfpOFzfPL17jggkih+dwNlOhP9B64LF6lAVCPH
+56gsOXMKB6cCTWROIZvH0PI0llnWNFeMP3QScgam3jgGLUU7Q1XhsprCfba4ZluW1FNJ5aoFmDu
VJrmz3QR1N312xChPcWiyf6ojhAK+9Pn8L5kkRTjWmzwwD/3vj3OgH6Gi7EifWwTCODOBoSX2q7k
HFMVph0464Padc2Hx/6RA3mdLeZ4XIigNnGcrzuK+HxWP7kTQWPfoW0w47w8ZLvzb36tj2YcWxi9
kgr8AFB4EBp3R4lcs74vpR+HpVijRcfidJ9NWK292NiPy0BIKYW/KL32pr9Y5Neh6jIVSucgTtb7
5jC0peTNT40l0VXVtlN73yig3u1fkacs8fPGCvRnyB+KxIBAwAJ/gSxibCT/QBMIWUXawi8OlKHM
tq4XGyIQToxsgrJbrHqS3J+o1pVvg2q+n9jnYlSpxp0/k4dOToOo8Ql2Gt/0gan1llXQpKfsEBNm
/hQaz8BAMObsir+JMg+i/SlscXm4+QFnU4ge4qIY1Kc+RYfKtWOgS0JQRtTMCPzqRKq5rJ3F4Ol7
iKahq0CHo3eMf1QmjenFgCxK/AyK5URh52YnP+GKRdurjHyjBpfGu+y3ZHt9o6apgtvhJQLaLLW2
L9n+0XGdbmmsheBnEL1sD8ZNKYLLe0oR67/RbEayxtxRj40QPYqic0bkfFu+dpSTNwv0DsDvE+q+
oBs6xvbn9BluZbZOzHoqUPxQw0YgyVx0nEitJ4ouds+fj0YUb/d2BImWDVxNYMzBWayH6YLYTlj0
cf022roW53zG07vnhCO65AAWt4DW1oEPYEp/85LLrE4XGe1oLCXmTY9LpXxvlMgZWRMUUv0J1gEA
aCIznv1NTG9QD4qbowqpchUpeW4WlcA6hEflHyWNbIkB8MSD2Ur0uJyKMCBDeFqlye8SgF5tdgyL
J7v6JjstziWbTVFsyxK8KuiMTvkjudeou4IZBwlRq6y648SazIJVNJ6CxzS1W3ij81qjf8eM/3nh
H2aqrVSbAtDseMMtPxnuoHYVnpyfJCb7YdAvK2iWxcpqVObQFzrqgxnht7zn0Bfp+jlANSGq0zR0
Lo6C72SpfIWLieF8FHfpfyqs4kVMLSwzqMaySJu1OLqgPYjHA+LdmPvDQh8pyQzXDRxpTWS8cqnP
Ur2C9Nfx15sKSGbHB1Cqpt7WLi2iHhHB8hOMfvoHSvYprv2ac65x2Thh/VkccY5+S4asbHbRQulA
Dpy/DzuI6wUnNCiJ8NO/DgTCCZOMOLj76t1xopTEDHaAugeWKyiEXHKhn1GPlIIN+0dJiiFiZNOZ
V2dtgY/JYhgosiZYhorRZVkj1+oxW0LJCrqgvJ2TqroxgoTUmcpnLs4LSsHrByFUSI88xpDeKFJf
/q+B+hxnd8neoc/aajRxWXH1A4OGGceAc5NkrBjVqUmAkURucECe6mXJTmhNHMWHIfk6Un80DBda
XGL60bFToYXgV0YNtCnXRIZvLp8i/qyU/VvFYvjeyGscowMIRlP0/x7C9P8OExfwZSwxavx4/g+l
ViKvVSWAspP8qHBEqs/BDzk/YeJfApK560pAThpDpUx8SWd24Fnu7KgYia1sDTKjFKOkVx+XM5L0
9ZFJdS7JiYSinaZiG8ZTCxRhzbq0KWcnUdpxPzUX6Y19vVDpOeyJWI0XRKAc5r2Xatr036Bfcxfk
jrsmkGZUu5BRIMPaUUVaZzQZv9k95tTkAtmDZr4tlKXJeXTo9mf4W42Y3bmxhYwv+9A0mwrL2tn2
uXxauuIqT4UYo1ZRQvwSvvjIcABw9p+daG9524F4L5q8bJ0yRTK9M0Vwozb0ddo9063gjULP/XnZ
kSncKKJXG+PMxIAZPI7VAUt7gVmXHB4xQxzpcQ6/Vjt/nGIO7MOJnKpzLKhKCb1M8oy0tD/PyKJm
U6axVW/g0+w/STFhzzoKrpcdCf71+vleB/C3lMAnceJpwMb9JplRRNAX3mXAP1B6YRTg+x7derVL
siIgqCMdamiY4BkMj68cGWoEkPKU3wErL2odyC/9TrMakGFmHwjNauEnGismoCXEXi8DsSLDDhQM
R5DClXLPZBf+ZXIosygos4BhWKVQLmcVvFlRii6nL4nerH8drutL1TnFcxC6O8Hwwz2q1fGjisd7
zq/bMLQPGeK5JO8bHf4sJcRi77RajKKdE9eD7LX+WPTQfS9gK/EQsk5dvMiJadNmohg4Z5XqloKL
ZtztIrBsLb4cZ4/5UsaM7J+oFNSM61c6+XggvDdegQJV8vF/Qi3dd9vSP/KlRndJWOXlrMJT1gNu
GhmqlRj31IbISwZ3iHNSOh0daE/Kg1IezJQE1gtQlcsxRrqTs3AozfZ2uZVkh7PxFnG7LPH1WOjE
bU9a7j6vHtXLmoqvgCipIrOWmGTwLLvEV+a5FYBImuIWaeiJRpGP+ZbH6i5j6/bs2aAGSju6H2mS
L81H3AoswEg/YvuOSgfDET7UEm4y+lBPJMcESedy1lqLhTnc9IFEUS2/D6V+zscPdXY4wBmboaGR
D9iBEKoiLfQLyFXpcNoAHC+CUXrZ6SeyE+p6k5Sjv4D1Sdf1v0RxiC8k9SRVXaLPYIo4bSUfHuWR
Tv9okj7JDn2iQL1L/djlS3J6L/rnTYH/D6x4G5JBdNum8DLR9EHeeKzBsL9rOtvgYm6D4SLGDa9R
SujD7VufYmxL0RY04roTjDG+ysA5V2jipc0DqJWNxG/E6/g+9MqEaMTW0O0gAZuC/W9Q+4YuFZZv
O6vQ9QIh7jdVNVVVrr5SHYdZFYuYeqj1XDCZOKvamMFuS+hmmjkqEM3qupK8CVUTKl+aK5rJ8mPb
f4pZdQ7QbUUSXlq0qqUH0YTyXWBI4vBgrtx6vxZCerLbCbYpF80V5hhYgulndzUTlpJbMnD8zyoG
GjxKeyTzbemPsXrWueuq15Z5a7zDFFJZ3Mx+QRLIBr3S+ItA2wa1iTn4GWB1xfT78I9Tjg6SchJc
hpfhkwIwg283uxAhDtxKefJd+dlC7wy2fJlVlPlhtSxlt0clmxWTPQd27Jzdf1AHiXwPhw7LXKzP
w9tSzKrk90gAtvwZtDC5vIGqH34vVihpuoHhmGe+RL45zLPMKmNyII6/Ppnl6gc7RfuaoqIb9eaZ
pPxvZvMHMD5uERcjHDymF8HhuBGZNk4hHz/zn+iD39nJI0FwYVz6QEre7Xbq0TSR2j3+jHVGnuPX
0SuXUHqdqmz82oeG1YlabH5YzDpNnR0k+1BN5pFFK76v+yIAhV1/qB2bKRjspY920tddJjEON/v0
3UpDK6cbGpbnwI0oJSCbGw74kAJKXcK9ml9CMh2SoH5WCTDzYE0VvuxY71uFUef1jfWksgRo4PhN
Wdg2uU68B32X5o+bynnaVOTFbRlOMEwPJjJRUt3HzgWhwl+y4/99pIDqLoDSY6wtd2fQ87CbIf7K
pSW5snwYqjGHipzYt+xNLLH5U053587VcNwb2cyT48wf7RztAZ0uaMLPwFAtaA1KqmqYTdVVYz8M
XGafKPnrzG0OEwizyvuOZroFyt82bYuXw0gqWV5yFs4N4a/oNKigxjz7XZmJitTIO9jyGkOvHX++
QkuBNd3ankPTWnXaxzqytLPmiefyLl5wk3Gslpq+ee0sfzrqFX0OCXTn9pMyc7p2jbSZxQlQowLG
uDhtj3ikTKCYnLRUeqJJt9qloVt0u2W4wEF7tv5AFoXqrY2k6MeJtRmtr7f/tb1LXTc6Bu9nVEbk
5le57dEyF7DiXSJK/JM/G4P/dsiN9sT9yV60djt3F25cy7R1jJilp3gGHjVY/xrq/cxUJNzp/BZd
JiZoEIiucjIqPmJ97zLHSrLN+6rmN8LKhpseih4Fq+5mq4NvLL7T2zDzR8NHk559Fc//vP0LYJWi
iG9HngW6lP8j2IPB6BMceqodxKZoz4Dm5yLZPClhZqPHgqv0pcaZayhqVDyXeUWoNNOMrfaXdZCM
XHWfUA+bgYglH76UUInX8fytbsJosK93BOsJbp+to19O23unkbjBuyOmoOBJmCUyWeBlm1FBfvET
aEcyfHuhNY8fDt1BEJEw5uHrP+9AnC69ynVA+JDsFMTzMxQrffSTTOIsL+D/m9GT8b+v9/ZXPcRy
EaF6BF1CE0GSjbMA4JWMpqsEv7UmO4YIFU+lP0JX4dcs/+RQpEacQon/DaSVxX1OZBhv6sfz6y5B
IVOnpjBgpNvFdUX/vq3kK10fT3tnOGjWBUeyJVO948BzY1WVm0heVOMLcK77Shh5nSZJKcDb7HDF
mQ5cvlFb/L+aOb1g+M2jeiIPJSfNJFJKGJXhcvnDwWYR4g7ABdyNnmZGgSqMx/pLRSzK13vPTBMm
LeKjUfvmEvjDxsqgn8dfqWu5EJ0VXO3Qh69QzZLOwxdWFkmX7yvbiQ9X/pecwQA1rbUS4JMDqNRy
J6Qy4z2i5LXbGhCEeHJacBtMN1wiU10gaRXUT3F2yRqqpsfV4xtWUiTz6N7TurgC9M2exJ+Az0rc
/60OZKgy+H5/cuTRs7rBsL0AERwnApKNDPNt0GYhY3TB0J6vdWLoZ0S2Zbv4rK5qyYeHlqan/dem
5KdlTF8B8mHsn4+IquRIXaZBujSEnFoV/VGniDWK2qoBzxzBGh+3PpJGRdbLyqxAtOg2kU/qxN+n
iCvOuUQBRGq7wlF6H5Qiy5G9kURKboGcE85tVy1S9eGTNNkyTmJvBvl3CPT39vg0iIEdLi8P98/f
ctHVBamxdc4tc7rPY2ONVZKYZU+n3ZqyZbWatmT/bnwXO8exvogXdCvzhYyPe2ia16Jt9chBp4iD
M5RCZQvm52D23JELyzjUMRc1C7fE1RbKkjOCY7k7f40J/eFUtA2LXKPNrzk5SQXywOgY1LW/AdOI
4LtCGjnfEVXOCLQp10H6omaqt4DiTuzE2pJSoNbK/gOJVsxIGDLKW3BcvuCVnrDCUmuMNA4qxHgD
DUEq3mYkPHyazL9mUqKVl5ugxEReE8rVccPzxrZ96uvK+iCMPdj2bgZB8DjMxxp/wvB4BQAzrC7L
8Y1HvMbF/M9hkQhRtBVeLBZ/7yap91PLYi00nal0PIWrFJHdhY+M3IFNxfQPWV6z+ocULzcs0lv4
O/q/mRCykQ2oIVwrSHkMKufnT1EgqlZcBvmBuDAtumvZaP4YcXVWbnjSbosjBq3oKL1KbZP0VZcM
kUhQkrIfzpH1dWmGuZelgyLE87r2OO8JQW6rCQgSL60g1LtPmyjQI5XGke/4I4c99TmCJDGCdMlj
CgHDup0oNSTmlXPpuGH202hlRorNPXdN+klyRyijSWd19baH2zJH02D7zVSPPJbCgkX82EVPdywu
IwGD91oFpo5ZHQTP14a7fb/WMKZpq4fiCC6R4CTuMdUxAHCN3X9Ssrg1D2c7mmW0cqnqmxGOzBIr
TzmEb+ZPPJOOyg90mQA90lD1zOaf4zIMlOcP8au4SG4VS18yjPemV6IMOyAoV8vuFsYBU80zLRK4
fzTMH+8i7jolFHUy4vgmMQzECi7R4nMf6H8xQfIrewtlqUb+IyhzStVB5UoKLoVtUSpXnICFhhOA
WM2E77DIlDHNJnZFB3kqBrqNEk7wFy7g/jCA4PQKuEQcvUIjM1R/Ow+d9ZDGYIyzdDTwRN3FkWv5
Lc1ieDWVnP5w2HIOw/wpcEi63435ke3lhREOYKOUsr7lR+NeDq4QJUWJMphrjepXclqk0IYC325m
/4Fp4H+d05u1mvCtx7wlSUbVpjeoTzoyLPbKwntCpjzvWKovgntk7FC0M9jOlqqDJp4C7gdkoUus
pW+5sgkOa2Bwk1L2JajpM4W+4dZ/2HlTb6g9/V5TKR34vKDkRhmwGWXmvqe8vYWy84zKXjEAcBSh
FSOLZDr82zYE6TPLJZFyA/Ax2b++uLLbBjD/0ffaRhsbCW1vwhodAd52qnkwFgUdFecHWty4mPO1
KVA7MWBxOA8SyJZScMbk3TbeVtjQ3Ws73c3Xg4inWEFP2JQILcpYoY4m/zjaCTP5wGjWHZ1fR3fy
HYQ3MxJP1YHHLWxZnrBLbD55IX3UNBZdCpXt7S5bFbhhp+WpbvKWtZFJLJI/Ood5x4jmEHfUl8Z4
47ZTrUYt0s1UwLHReWqIiO2Vt+XGd4dSgeh1xN2wnWcoHE1Hp56COQo9ANJMoQ5bcaVZvVmtGlZc
pF7RsfK0Hg9YMrLiRvTr25zV9+xgtnMMOWgIQNbubVdDZZyRWrKZEksPwjRMnfWHYLUgeJ0/YOoc
lwq3DHGuZVLB1eRL1xlbygvsMCcnMdZcfSfWoMH2yhumwBBDqauQrVCV6A4Dx5WIYGYiAcYOLAyh
aK7G/P7w+aA7cuAH+OpcmURv6fyOhupAfMESXbJ5wWDzqHY/Py2R6DSnmdGzFeM+isSfJAUa1A/U
fv+7g09bt0dvnXPqTEG0HxIb1Zn6jDbLn2Cy4YomWbjy3cXxAFg7FSLE9hsnBViO86UNR/PHDkzT
cvnndB6O/WEDuPhOtNFQYBJ5Fy6hhkjwpZhNBYYoJEf3xSteL1r7TpzGBNzW7rhYcMGPi+1QdvG6
IkSTbCTn7XM3Uncspk7F5bvi/Xbc1bj51bXHCdFOPYP3CouaKqQcau8ZNaoJ/IqPa7+LJUJ1BvUj
Yy0kgpupje8tnj1wcjudwlsJuoKvj1Mp9TJntXs5XR0qMUrtkFxPoX9Wf2Xg/ZORnWtaG8IQ4VRq
QfAx72n/P81H3GexJFKmtwu+sU21r9ZP28jtsVvx6WkuU8uFPQAZ+pZYumOdoGySxDRlgtcDhdC7
1k05PwhCYDR8UzRBmbCLxRvUt5WCsOdvxFLwB8Tq+UrCuTOaS7+XilNSWSJ4Z+SF+7vtvkHHnM/n
aKXkAg1bvWqr1CyF8rL57qsuVEpjIzQwMvS1NVKr6b2gP+c5TnqBCTH1UqxLGBBa1voVkkQHJEoF
Ir4v9KDx2ObbAs/alvLXtduZUGipnHwXuln4Le3GhpxwjS/itciSmxvOq7Q8cGNMQvfQAjuB6LCm
PS8MhYDJXclzpfsXmrGUX2GcGqDsGxmn3xfvhxU3mJh4ZPzcfebrvAvL55IZzNOGRUnJ4G3mEF+m
kQwmyapLk4fQu3A1L5XE+h07fOxUN8UXEuKz7OzrNWoR7092mV89hPa/81exiJNog0+Jq8CZtenb
mRT0D5bHgPsLYcOkMhTH6gL179JlW8zOG4VAGP9HXPnzNRF3Lmw3Y0S4obKdzKIYKOZMDoEEfKWj
96xjb7jErK37B4L4X17nMNDPLYN4WDw+gwpS33/K4WGW67Z1bg+NCultdrr3UmovU66LNiX0Gw7U
awgvlYxYkxWktb5r4YFVLQeMGvNjxl3qah+DhKZcbtQWUrh6ASUMoctHJw09fzSpMTGPkCiqF0KB
WhxUkVA2y9T6t0HuLd+ZkvViTzcE/TB6kfCAw70Ff0+F5IMIp8AdWxIh3fuDLWkqvslQKKies2Yr
ma6L4ZpD3FlmWtG8gjv45U/cdnmOR+5H1b6LfGWU9hJvNI5R+e+i78JByabxgDzVU6K4mEANeFm/
esyV+PQv96Al4akGSISlLrCaR/2sf6tk4lu66QuhwVcByxi8EJWsPVDpabfAkV6JetgRds7J7QnW
Id1Sl7hPwd/XvfgN5YA0WPCrVdhHwNS42ho/XLhHLBpgCufwBVi8uqv1VHJrptM7Gi9pVjkJqES2
r0HdEXTgAcWRym17YN/1EC9pW2LQWGDlLoeBvQgHdy0OdU6tbkRRtLiQzpRICi54XYW8EZ0ilm6O
8swioKKKbGsNS/GNEoxzNl/YVrQZ/BAY+kIY8Lja1DkXPhhU1HxWrb5Ldl8Lp4G4AvrynMxejr57
1qggdkmrfLSANVRg1Ls7E2jNVg/zPPRoHmuI9mLQAu8d8Ez2UD1c6L47a3Gz/pEIdMXzsssWZJa+
45j8exfk2fREFiPg113oKR7f9z5QziYi3Kv/oIvArByJfNEyXGQnknJVM5PsA0D4h5lwNFMfzbXi
EUv72963w5Z8gqx3ilZaAlRzQkFPt0cTF8yGCfeJWxDoJmoUgAsF17lvTsldzlhWL/dJvi6mT3A2
ehq3pPGpjvosJuTugM6RaTzSdyFykfhERfellbP1WVxrsTPo7d8AhBuxMr9N7f4350AYRywdlKWA
gOcXNr4uVJepqXDNLlfc39KTXg9T1rmNmUKXT2ELIgwGrFP2TNj97E7+iA7gdeQQcHXLwNv8+HvL
GLJDlBpFPN+Rwru8LXngJfyUTLgz+bEiA30LbsKhBpXFVYQVAe/EUfg3v0dl2DIwHdBDXRFH2l9R
R1wQfqF76iMKmV/LFf6HH6ZriIsr/m9Rla0r+89svFq6EjtVjieyUEysQcDJkdBLdfodgRCUWqZ7
DEFC6a0edhePwb77j45eWoDIz5fmWXYRXOkAO9mmxO+Cs5sS/Pl7k6u1sd4WHlaTs1PdBNHMqvUN
CxyB+GyEgGxok4uJTXdMtLuu3Jlt8cH6lzIDFh+pGQ43nHgmlG9dJcP3AvqC7DQ6UBuBBBSpFZSU
aZK38OlYuqJ7BVohgrPhHDwY3eZ6xv6Y7N7CbNceLLbgy9bBVJ0LatwRaWWyTYm/6FlHUnLBPNwN
0fqgaTYM4ZdQs6vsnc5rULJSfaF74RdxtxCnkcHRhoTMvJgSAbOOQ4dYJ9U55eCeRQO7hSsudR0v
DXKndZDr/6gIvM9F6d23sTdVGtIpZU4DVljE2icS+5qwn3Q1zOjxW6hFw9nASZH6S1yih1PKs/di
oeXPG+Pu4deHAeivkWAvUtMPvpm0jNNWAxE7PiNyotxBHYM+HWXmZZo76Rl9legNUpjw8CSLrc0o
QlgGULnBfH/+2BXGwEQ+gfJ8sUyQJC8/+zXNKm2Sn/EZS8M9wk1ccjJWEeihd7R3tXzoM6Bk+pWM
njZ8LAlh7LtjhFfYPMsgMtfVlW7jZiGAZG7R0/nLgXzCha85L7KN3P+hWYCm7Xr1uFl/w+lUrYOz
8RxCdHxOARnJtDGbr7a4bB0IrgCXJ7Hg5x1KwuUtM8Ii5griTPrPq9q9/PZ5eBLEqUfWK0IzIKQh
uzwn4YYr3H/Gwr4o2V207YC8TyEAPvrQ/KmhWvzN6+MzKN6AckhN7Ac6iQ6wkX/3AdSRWLSsM82B
V+4bJ71FiEgaTx3GQPu3bB5YdSIQzurKI8TU6/smRLOjuxiDJ5HlOtCZRCzHL0NWD00TVuEOBGaz
fw03ktLeLOFbWjwQf573Q4fp+tdcuuwWcG2ma8qDxGmXeSb95MClVyjr9zvHn/eMRcLEl9cmkzr4
cwBnxbL2SvghKHRaELnt9vkdgBMqdVe7gKhJNqSP9j2hvJlhvy2EisD3mXFHIZ/GoZoZOV1CPVjr
qjSw07+NVfLXHm8TsLue+0BZ2DFs+iWT7jQBN2o3QuVWv2hgVl/Om+dk9jmfSSM9RbPr/s84WNf6
g+yYfP/xK87Rk4oy9uOxOgVrbV/Y2q06AmnwCXtNqxbYsR8zyW1ojuOmAGXNuTiBlL9KqsbN+9jW
Pf/aN9q2SsLgpwgndUBrsMX7Vf6W6WCRQIkp9bcicGp9XnZ5IireC7q1HBNioYijpwuw2clfeoev
I3SJ7gb2+9mPmAlm/K9JCLLVZYuMw0D8tj0Xw4uiOpnr0BjZPxrd7t2pFtKc0d+pJBU69IQxCgSW
g9aGsE1jXAeRcz1B7V1TMel3KvfXsV14s+FzKXrWBkFS9CCUnNovZgomX9Npu1DMcNQNjFo3lRC0
DFjdY4D7+TAJabL4hSI/SSkFxkvClLNhHeGzCS54HKRKHJ9LHfd8xgEOsdnUZQYPuI0UMOXLk7Xh
gf0e7kWie3RH/uEEj3nLTcS/KmkVVQ75wP1Jh5jGvrHCmjkgF8NCsIACiVEScSdQT0r5lrZuIRQ1
2BmSd/pCUKAyEnkbrBDR7t+mASnFh3pSecUkVwV2vFAMgYTMnu5r9FXv7lbve1ZNsJ+mtmk6JmuE
YA5EJPOd6dWhEnKFooRhpIdtwmD9YKNFAv+Liht4T5jfjbD1h4CYoyYpB8kYq1RcvuowxcmJYW1p
bbmbZSlvt3IeA+YeYlcgL6dJnBIwvGluDB6xfnJ0Z+mAm7CUlcCut/BKSex91Qvet7ddp6i3lGUW
FBGc2mQ2qF8G3TCFM45oXsLa38ePmIS7FhOeh7b7CML5mvIJbqLlFpWIDe2ERP54MZC5hIgShryu
J1zgv00AG/8mOrR6XKeOERZ+ubyrX3p59yBhZaF2Kf71T3/2SJtlGlh6mG+6k18XluqPHFJjIvNo
zpWFh/mZANtzZRM5vfooWE0ewcJuPORPJb8r+HwbYx+jefeD20FMdRXOKgw0WOWMqUGRJussEh1m
g6mqyxd1qB91UJg4r44/kcBomIQ1i0hOJRpw/dQvXaufdE508vO1h1Txy7omD9y8Fo28vRWxNFIU
nwt+hRt+nbAxkosN52+Im9hI9dIKtachN9H91JXXUNg2BgOUeXSy+1QS4EDepjA5W7CE0xqRIWhm
S1qJ8UhUVt63+OVfZqns1U+fK4TbGGMO0IbmhghjFMnZ0wOlpW5ILS7+SbejBlXEfCTI8VxX1s0b
6P+eeefy2Ab7CFhDcEvcTYXp7dtx9HibOn0tVnohJn9t6kPn5cCKU1mwDJoSUSvWwCAGe1CufgDQ
bjuNIL2BcI8ucY4rSrM5NnAoFqAlwvRIfZj5pFGhr4cRsuXqyLuh1NMf09c9omIsYPUmrBQYOBrv
CkWSkFjlBIq09iCrHAho1tIt0vabBY3uEhstfLT6dbfOsA5V/eak1+Hiv+CDCXI8Zap+XeI8AOqV
3x2mQIPp8Lw9RIODQE4xpOhnGNybdYhSjch9UdbGXWyLCkxplDw0aJ7sAKp7ykN0IpJUaAvwUvJK
uYuYUlCFxffIKmsbxqjzqImibg6XsxCEpXS83z8A1jA5Wy9fRFS6TEUgoD6LtiHdFD3gTufk/k5I
MJivAiMrIwTgVV0jgHId8nzD31DGgjDDaElVg43fdGRwVH6MZCFIrJT+82XiXJ/LuRKKLgEad/z8
Y/sJaQHF65vKLqMSzdQwTGPcCKeSS4PxKTmmoxGsuw/8PqbajuWLN+M6GQk53+liA5Q/001OUzUQ
t3z7XwBWnEEoojoTWvJFDX1XMbJrJB96pJmZ9n0xYN5c9rlXpoa6nJQjsdLiLq6uxAf4JhOzEFDW
TSFenQFGYFHOcbCrePtk+cbh3eN38dFhMtojtqozUbOgJWX2qVVNsuN+U4PrNyHvBUwofJndbee0
Ne3fIqr5V1SL4yAq1aRSzAp7LR5kJ6BHL7erC4uq6mgRtdDHKBjO8P8lZsXzJa3OqXPLfPtJQBNV
BO1pAemdqpmJfZ+jqjgFIULw9A7CFnki8IiJNg4i3OlGyR+Vh1OhhsbEmJVzAr8db0gLBFM2frnX
IIoLABRZZlj5yAHp6yj4+JmxDv54joryhhg81hVYjT7wlRlP6Qt27D9qGdgfMvZ1qEyOxHxuEbpX
nYCLvradAIgQq6Vn89lswDJzk31Veov46ifkIbmVRX1XIk7LBai9Sd5sUqpzuaO6rXCj8QXeK8GH
dhFf7lYLzamUOWte9t3aS66yuD+pm1pMyy1YaRV3hPosZDaln3VwrntAE8O4Nt2uIRpD6LyJkekO
xlduz+8Y6n3rVHf3Z+xKhS13sG3PRKVsSbnIWXJLRQ5hIeRJ2McfZSJTEWgBVySg9gsuBhPFkK3o
nBWc1Zpw7CfvhiuB8/EOLMxLIM8vNhBGcZKt/HTWe6qaht/b4uTy/ggFbrj2XVY9QMMLvWAI/jBv
EYJdXd1rcJEw7CtO+pO8AK5WvconJO12MYrbkJVkixECsGpPbo8+UsqHzA4ZQAwnoKqq4suv09mx
3bHWQiRkbeENZxymZGII01siO+itXTzuO0d7qyAFCCQDmh/Qa8Yl01rezDJzRylNbKhLBCgSLird
wwe9lysER/m5qiqDlBDh3tAbPxN/c5D2c0WaGVp//0kmWk29ly0SSkXyRO5GigRFiZQyNe6KyPfg
y7+laK9XCwyq0Bxo+F52Z7FLgaB5M+3tIOgVYiaQWcR2ifEBoQmvk3OGkFjkp3RN6QZtNuyc2b8e
U5RWlVYxO6DVXt3HJTPGTQSZJrI+PnO6uR7cikH+O7U+WOVC7Ms0nfWVr/1YXBCGzzFRS3KEl3Wc
bCScEp/DTK2m7plQ7zfB67YjSUPtxefeXujBv6G9kKEmOzWaAnq0nVynoj5UKJnrMp8ok5UVEf90
FKvqG59FkCxaKp7X5f84EgySqZMxUC56LzmQpvlLJqr8H3VU/b0xOND/2WjwQ7jKCT6o9QTmco0B
0ovD8okT0iWBKnSzpcxHXC4FjOdtuje2z5ETih7lY2O+1pFocjfaP1irbKPB19mAJO+DgakspYht
5tQd16q5+YWrNzmBrSVZl3yis9fXYpFYeOGgA2nWjYy0DOYSP970xQuvRCzuMVi7D9Yp12dG74Pl
dJyR7TjLo/sHSMP4N6TrVp61kG2N5LatAtDbHvA46JwyC1rOhz4CHlf+6P5BetHGoxr0OXPHxptX
pw9YmjFpwZUvQkcja5M5wPllO/zqzooFCdebk8LwvdA1sKpRXcI1mdk2gQnUnzkzcPj0VOKZICfu
63UYRXGLIn4/bCRdHN9fnb/QjKwH9kiW3Xht4PCVaGVgRPHfYMLy8/KWFNRZ/yi/Fw4lZ/uafD+K
+dvrFfSLjcGDNhRP1hG38G2EvIhZyLE1zpQM6eXmpZH/5C7tSLQnVPXYBYxEFJW9tDsk3lzbS7H7
YFZn1CK1SOIpjBwESSohYu1191xNqjK9A1rVltmENUuI0Qwa+/+YGBupvs/lksnzk21GliynkS24
L0Cn2mrpmYJ8BE+rAVyMbIcCYbQDITfeDr6E1xp8yxnHG7S6RCBZyLBwJW/gq+9VE6RAXTXG0yn2
Vo/+w059//2pvrfI1RNCEwIrFD/8mfQ1cs2x5NsPuTS+OgUvbz6QxtjIZLQOp40vCKP9xdGC95et
PSf8uCkNxV8cAlW9u2REUIll+SV6KZBH5Nk70zv7Os8iifi3TClOu+zdOXjdBTuh6Pf6Ii1vDCPK
tOXi0OQPPzlOilM4IJX2Q0XpoYx4OAR7zBY7PtSsBSkvzRrxSkmjkh1CCe2RFrsxtk0rcYCQo9TW
GvhFgrA6EpnuGOmt1+LbFsdkIQ/7+GonWgvpFAKmRiNJEGtLM+G70hM0qW/veTSQZZbfxsDUlzlP
JHoDHEOpzifRAzeORk/c+kzzokdfjVF0MobagPLKWgAXDODsBYZsSsTBT6MdAb0Cqu+0Ls7MV/Hy
C8nss8hGdfO+Cqe7p5/aOUkFzz3lXuT3rpPb39LpusCr3W+qQHSW9JT89BAXIVb0V75or8nuOqhz
52zgfGWtdlFLQT5/YW2W1v1JDEujPMMXa1f3QIw/E5S4uJqKRuw5OJzdUBj5ijRugWC9W2g3UfPC
P65DcUNBn2IVOjIqasBdS7aCOdkscbQsEcBrq347fQnSB5KSapKa6T8FN3zypgiAbXEbKs4YV898
BJvQetV9UkxqKcvy7cDFG9D1JRcfQFJx5ovJNLgpvEJPBw1Cm+45dsH0DiJT6Jdb3SP79l7mBxI5
d0iA/ohnI8b7am8t51yWfFx7ofANt92YSehZKGJX+s8ztK/It2v7mUr8Edeu+7fRqqFRFpcKKn4B
tVzVZ/f1jpDsddpru/iBt3D/xwrdq2588qlAd98YcRudwQ6bNtrMOo6mBlFyM/Y2AlIefCN46fXn
zxrDvXyoZclYlziEYNhvgzIYLtaA3E79deDYDyAy7K7tEFlCKdBTuaXZ9Gbwueun+KB7D/9z4sMj
gKrS3KKmB79f9uNM8t64+n4a790r+GDfuBxkOqXYZoGqtOHsJebcQNxuylE8LT1GwkBs+MOJRmV1
uBkh1EgFQ/qFjZVyDuowEszBajHuTK+ZxrdmyMNN0QUqwMhNlr0Jch6rBKC9PwHhpQeRmy7dkz/J
eNr0xBt0wJwOrCr9UW8whhN8fbWEAJHfzrAj8j5HOATPJpDk3x8jv99PAQfdlS6stMI5ZE1A2c3a
hUv/rbCOEvCSdm6D/iiO54vt5H6rTAdEYTZfSaEexUvXn70oLLclznvGKdNu37QItxcuLvgX1vr9
/hwPwCwMH0uMCixMn7hYWUmteEBZq/EKF5D/BBIIKt8f7Qj1ynbc5UjZy/GvfOXKJVT6AQABhyzM
eOIKbgnMCVmwCNqQWjEVCtABXTFHybN9zpW0dsBjYSuzMV1gZ3J+u3ySffilL+8lVUGJ+gU0tlfH
BWwjQWI7JDmNnB+EEQvYgAyeoUEXKCSNG2+qAy9Sq5+QVuzVKP8uVjkaWtnYI43Ns7ub2sucZsSs
lry6iqflqbzgBn4QY1vAALJgKkQIb+CcpNlkox8fVxWmzCNZysXF+VluIvRJ571foNzOx79rXoTc
i3yI1zVvpMUdfxDh96MT0Uy9xNHOKvsMPSKqM4DRSTk3DcJ9ggzMFbqq2dFCWn/tvJi9zs5WiI1h
2zSqap/Phhg5xVNTDmTXukPA2bPYnAsuKNI90pAWDUMYz5DBaKSpo7WKjv7OVaNGhrRe+7kQkhRh
dQhuOJhO5SQZOVBlbuofjvvnil83U9JRsT8ysfGc4PkXW6eS6nQmGiAOJJlqz0ejuUK1P+oCXY+3
c7U8mtbv/pHuzrxtTyOptp15BZGMFAGJbZcQsCpcjgOQ6nanSPrkCBq0JM5dhPDYe1drQj9TNfvg
3CltM2BbmD2InlCWGyPhPr0UZEVzDoXxjNdEbxiXKgE7yE6Xa4NIiGj/Dy2kzKfRy1eGmoy8/4DH
kxNxs9NDhtSPqyLnQMtUHnQ287aSYCrYIki8Ye1H+6SUGER/YWxeBf/je3pMMT4r09q0UeIoBafn
k3/IusyCW+OdrJfI1I68WPLHt1DGT9YzXEusx6yWREkfjwyim+ybCi89xUcTRvqDUEwEblSUNbaE
jaAzlEGVjq+O8OQF2hVWgb/TvZ2RmDatcYuR5FFkACLTDIjZqNHocxwMLaXZkeA0WNrTCpaV1w4T
YwrHVO4psim5UnDAAu+ui9lgpiN5uHuFQLv9+ESUbtxyX0+qhrTOc+d+Q21Br/+IULaq5UuurcPl
VebWzN3P1z9hNbuG1OARqfFYajcvexh9fVkUFlX+P3v8epAP4wuUhKtDWrQDQTgumlwwWwwxseRB
mIdEW0Lry2YMb3n9qpVzHxTx98kseZ3CmBSAuoowUmznl9Sz6UMyBg2KJl3CAG+CkWZvSe6MaXHI
Ic1RqxCXDtp3KnZlqseDe+3+6wC/5FGpyjtsFPYbJd7WUPtuKIMjnpJuRc7l0ujDIc8Fn+u9g2X5
DeV45WizogU3mooF9Kp0RGY/YkuXFOXlgRMFkq9Eu9dmsCwbIN96mzSuL+QyX95ZpDD2ckzCI/j6
KQOBjGcLsik/gok6av4t5OCPdBzs2W5kBP0LBnDUyjdbSokvL1OxiJffjSZ+hTsCPOYB08ckUFDO
f83QZftiU9lDVlQRjyi2AOWGLaomXLwkR1LevnMl/7rldG5NplSNYOVQgUhlsn+7F4gx1MwV2IU8
FrgWcs/yyVoFkkxI52jwW1ONj4FHCL5YqRk7tBAbCI2xKCNpyUaoLch6M9SN0rEtLC4j/bp0yByQ
xZZdydyhqQBXhe5hS+GekxHTcrjQQ8kyakkq2V6hW2B/QwdjutJ7+taCqf1bv6yUPOyWA1IL9+mf
NaqzgOftQQqaccEiZpRj4znFPV8ZHtI6ZJ+DfgjbwRBHNSdea8aaJD4z8wknyTGvGxNeVhEHMyRo
GhAY3aNHusJnFngp2EaHGDZZnmnL4uAsvj+q0F9puCoxUAjeHhU9PmRaJgk/hhOUsdhV3QdtQYg5
sMIQ11DYxpp9qkwPwculJJEggsBdoUEgIkkuBitZzJM36SuRt9YF9nUO53+aK9HANCGPOMVMe1pz
OmQ4lkJN7wxjRPzralGBap9X4qwQLv5/V3aLoRxzOUaTM9t3hjXTtcqmDW3ZEnfnvDlcHJw4auY4
8yYrnOOjzLS22UrEQdraqrQ+m8JPb+XknqM6JPvVvmML52jVJc3g1svQkLRRdgU/rZNBzRpESxh3
I6ivlVxwiv+caV7YjaRcqd6yaCf2tdqdWqG0OFg1cwKA18ytGijYUB1Kp/9OFKLWVEsUt68fQxlQ
6vQeu8RydPBgY7XCLmO57OPbjIKCh03F50GgWhvFQyS2gn+3Y3uAJEV2W2tnb+Gr6GQMdFcUI2Ho
knb5gemW+OVyli3HE6ylrG9KYxL5WE+w5sj4YdGVVaaJmefrjO2Av5qcXR9VjOJCyXGf1DhlTxia
ztSmbooi9cgz6hY/7L2nphh835GQNZOo9N0cCTlUP86DRLu2U8keJfNiSggD8+vxlAeCfImVBwnr
d72RoEQzaYhgmfT+6JNmluX+uK1mdwZ7v4mJrgBM6zsZNcpRqf6Gjz0U16Gd/OvoTAdi3yxRYhpZ
CK5kzBPjLp6lqBE4N2MqzGuI+R4idOSeWfvKqviWKKmOc9Y6+u0rFUqdmfAmm+dqe47toyPDXkRx
setA5S/oEOyyoBFQ30274Pdhpj88Zj0FfUzqlfWM9bue9qhHvb0UoT1SLdk1lfxUxXfc6bHto1M8
eTV9GW8w4Bgl7Id9o+BuVOdqtyl7CHpGJ6Rta+fLzCBX12e1P2csGWXxPexp8hffnKwbJxj59D7Z
/GKoKXAYuV5qJnF7PS4Dwq6k44Bb1A2onNqNMfxzjHNWLn9sZ5xUuxRkTeRrAoqU0IdXuWyMYTXb
kbPujCXtOtY4IcK05YeX5DCuC/aprPIXU18q279EJUKAX8/Me2TvC4TBv+Ox7ac8X7daj7HeLLLt
sb6XAXrAHLDx+xJ5CfpXw39E3Pz6XRT/lM7j3nruXVtnHn3So86lrBcW+YbMLfCE9aby4M2idqCk
DC6kKDjeWUZVuf0//f/bENZerLAbuXJQYsy5cugbrHSiHRpo592uhmXpRN46IE5Z6lDIMobPbv72
YNsO1hdwPkLuFp/kf9OscAjAmxnrUVfsQTA6icBM9jvxXuUpBmVhSPVxyWZkEngm76hhr2SjKCNh
9wettmIkDBNL4ohsC6nS3zynuaajkz82+t3+NY4YdWIe9bJI3L5oei0deAR4M3v3V6uxIXIQdAwN
wkaXXb+ET1aj5tI++Om2qP/JLIuNicgsWNj/B+Xhsgjvnltn9pZoYS0iVlnUn7VTi6HeIfYmPbl9
Zx5WDYcIji6NGkKhuxBQWZ7+kW6TkYXRBb5MT9tSxetN8A5ujkmuGONhVi+aIAVwQ7li0GT2zJee
EwoLVHGpKI9W86Db1zEGGSNCs2AumgX1eZ6Wr6CYsPE9UqXXjHu432EBC9v9TtKXh7s5HU3UOkb+
N1+0Wr/SKuits24NWMxIJYMSxFxJHQxJbq1jr51hotiEdWg6ThAUpdBYrtg/qBzi2uKvGVX0RLW+
j7NHw1bDNSs3S9FOx3meZ5lR7XuQkptXo2iS3/01iZxMCsQTUwXmauXENCNwWtS4fI6n11WlRDUE
dVwxez0W2JA+4gFxkrffJFC8wrsW3wpsTxGwhe3poydegZJX4CBPNTwPO4j2wOjwVtnSR9+vAfhH
s4y4QXVYItD6tqCZ6HMhtlTyGJzGYGI/VhsTmABeaFv1zLm58AX9GOvUt7OdP/Jw3LXUL1LSEvv1
bonI35gDwFEtbhb6q2qU8tk5PUDEPTj0PicAv5vbWPifOsmYuU4W/Zt5E1bsbsj4hokaMPd3MtAe
YFr+DE8O2JySowazN0sTV5g10zztFYJTyXvR8AFPRIxo52OQHBLDnPN3q6zsqbHD+ZSPUPqKmj43
nYTi9/lEJR+knfvBm5elR+g5jbo0adiM86qXEP7oO9lsJ/6DZ+zZQqsytu7pXIHygsy/Ua6O0iUj
BrpwpL9UokfnF95VtpNZqakSKMah6jRbsTE3kWyTyVVjrqr1xxmM2Nw2/06sosmRTR8hBeOdIX+h
piKZjJqbMmSj9yxgwJTZx3+cVgtjK1f/LsNTHqcvdgwuynbGXV6e0q+MKGjlHv2QoynS2uuI+eSV
rZZm9PsliAsEA5qdNYAQTG3TdleivBb4NpYEtVjrPs67oC/AIev7P9W31Gdk2ZvuF+XRDcjnILG5
+PD9M3xGrZwCKtTIzkGH/lZZAGxcQIfGfB53FYdGH5T5FzI/TLeM1AyqpZGRMDGrpzaCI+Y0z/R4
zzhKVJmUSS+X73/4qnhKARWRMUhtRRBjGeNMrQRvgvACF0cGi7obayZYk6o/nE6Tv6p30VCynOZP
Xy9pmjo4vj32R+fxXpYouerJSwYYAgHFt+sHiryz1GbWrX3wMBCcB319DIp6Jp/xNPRSx8fdszJz
gSlZahdYyHWK+GO/OA0QFENC6t67rs4acOWbICczB/f2trCt1FL+qCqk5qGKd9vbGa0v6cEaamoP
XFHKWyuSJcBUvDKCuH3vq/IC7bg4gTSDff3OjHTlxhL4r7hz0PtDstIZ4x9i0s85KWtmRmMxl01c
1DCSF4Mnj6sr8InYb+pYnH4d5/HP5kk+EDWqYX3BCpryM1DDAP2NGNPvbDH6seixM9dsK4Lax2vg
xFcQNgSHgkTz4DtajqQTLzKQHvwyNwnUZ3RbswPImDJyfpxETffEn0RvVdHGDUp0iw163zMfulcn
EQZGTn359mReL74/QV450l58vw+zYmk7U+VJK6/mlZKgzEy6jo+ZS1DFTPkwTO1LdNOMxDUJqzei
YxgU0Pyhil/0t35Oo878qjCPwhJf+xt5/IBY0TlJbOU4xJnmxETQiBUNrfMKFMDD1S9p2USjwpBd
8ZGWKbUQv29ah84OMb0foHIiSa9HMy2SscxxGH19SwK38cEp9zQKwhHNwdasQ3lyW1/EXPs0uLDP
sSD4G2o6L7tFEm6+ITH1VDR6j0hwAVwr08tfYfkP0PoBuYlSpgn41W+JDgmMncLIMBWoe99Pr5oO
W5v38KmbVIJmPOjcBZ1d0wlecg/AoaEfQO6PpsxW9A/dSiVg/YIEsvBK4lVn337TX4wehAJsBeuR
PdZu3sdg4fdWnsWh0z18efxaEYccZ8fFUHlir+kJKMm7Y5ihmITv+GWsNYmSCV/4kjrxR07af3G8
7nBeiMAeyk4IjBEo+NCqmLUfJwtRGYR1WDhckjXBj81gQfXOG+B4SnnF0hB28wGdadiWKdxkio7l
wEo0KD7YvCaSs/BXRDCxLRFbLWicGEhoP42nKJIWY81NE6tRflomHjVPQsirVh490LLtvZfTUg8V
SvqURmXTDZTpV26YEMnizcbzkCfVOiqYqHvetWtFHzr1thsSO84eEWQGhURc/Hs3qQ2YR1opJXQs
jhxOwQ1XO6EvOV6c9EA5jP6RzFry2qQwoXRDDaAx5nstIN5uSn7udRQpwq/hBF039W54KoV0Z30d
Ip43X5kYl396s5k6XmH2slZUuSpgkBIu+b6lVyRGS4qKk1aCUREIm1UmBK1GMEKlZefe1uyXGaRi
6A1nQSKQ2ZIdkBit3qr1BHeFnGf0mqRtZrZrQ7H89o2PnGPxCw6CwKvRXu0ZMJNMpsae3M0Sapo+
4kVdu5UVnSzOIKGgEkGQsnZMUJapz1lAGG42X36M5LCk/ZbMt8t+AmuILDXpNbKCgkdilxwA35lZ
upyTqUTe4C57L56MLOd9CU2plmtzXOaadywahFOTNqJquYVePthN55xLEryAsDYfzSdg+ljo+tim
0xK75T8baQY7KwvXj0B/EjJxDqVLv1R2nWykzMNv1um5QiMVRGxRGIp5F3aYMiQdPWiOzyRHHpv8
lHryhtQEl+6whVh1q9q9AAwkvd1ClRz77kMFfbi3NqDJ1XhnQboB08vVNNnaie7Vu44+3JxqKLl5
bRwNilRCBEgGTHesfomrrMy+StKwoKhb1BT3FKMATq13WtFfUWE29qZIFdNh1/27uKgB/XElEF6c
KR8IG+h3As/lKdcI5ktILMMjDBuAYUpBtkGjnE86b3Er/QXJdNas2Yv7kQcBz8V4DB3zSKvz+IRj
H/MThyTbE2MIbN0PaoItrieqpl3FMlJmSlcwBnbU57CAzbzSHhUI5EUANQ5cbTJT5RM9ic3IQhZY
XFCgDqIeu1wGFNndlccd1DXID7FblF8OXqApg+iblS2IRlY5bECA5jiCu9U+NDjjGoekBVKzaQ8K
gPtZdA9VDI5qUo4Qrkb/19EAM3U7fE0eNVaJe+G1ncV4J4QpfwgEvEb2AK6fs0KMYb1fCfz0ZsJU
Au9ItFmDUYcUxCzS33PtxcQS5/bdXtxwU0RJyggbFvfqVhxPr9lK04Y1g98mfORS11B1xPz3H814
ydx1h/ETaU75w9HzU45Vo5dWMBR+WXGLJACz7Aoq12d6cTDAz8nkumoSA0vS/5dD1eCt/DHDOBSw
XwT6k6JytjlahP5PUYW1VWVZtD7YA1lM1fE2x2guAY+FllxTOzTrIlEdbBqefTMuV7V5K+3v9yjf
Sm2X43uuuycfvTngLySiCfUFFO3Sl8nCbPKKdIhu7EgTRtRur0zToHYB3WDYrkFuYIJiVNViMb58
N1ZZh9I8nWGaM5uY9n5qiBRl/68tEbOyoDunWyMBniFq5tQ8LJ7zqwVzhgfRE0X/JhnQsWFvrFA7
LNb28reJjHopEhF28EteYHVs+yQgMaxEfOBixmfdV05FnSvcaiycCLIKhlvRaeA4MnIUkgO4HwJs
THAQKlyTL131gl8o5pl9aBNBLXgsjzDRfkn39aFxlCkhEFAQxlKTgv619mY5B9mBBGCEXleA6W8S
tjpeQk/6/5Ou0wCEM56mbTkzr4uTeXCipgdZwpPo+ydxEmFSIDRZeLOvtaJ/ypNNzOTL8v/RM2AH
OvtmUex5OjzTPUjYbrB4ptOyAjdpOQCReg1LygcPVWKpesqAG8NE0kIyqxU1DASFnaPbK7ZRIoTu
7dkFjV7Gj3BVVFslFqJQlqKufeF0h68tqjmoizVcMXB8ZoKestAycgBhXqfDkpWNg2kLEjHGJDo7
vhIUc3HOtCrnNFEXrKboWJaRAsyiscL+rQbZS7hBy28t5b+vCbIc+0Dbla3iuskLHb7tYyzVgFAN
KZkVp9bZR2SO+LkMCnCExl6wp7EOK7sZvZ5dQfm8C9SLQfczW2MJ0Qcd1FEwaNvcYFp04Z2i5e/5
EcLL/8nLRLn952rLf/UamoeeS23N8A7AL0oS5SbZXQYzDtmvdE5nFIZjkkteED+bqqJfgB+4szV0
/SPEwJkaRpf0/Azbc9Zt61LuqF/HtcIihoxKHoE0y/T2dnjH3xaqV/uK5RVwq5VOmlJO6hs3mqbi
lpiB2SKsfCG0ywY3jrJv51xZG8gD4mpF+PgNq/tuxA4q3kgwql2zfPC7htN+fy0wo3WwfEEXGnh+
zg6v1afXwwz37iXZGTfVzr10cn9G+A16MNHVAV5OiV5NsW6q2N5Wk3cIELRUo0lnUxEHV9Ahr0Ku
CIfL1PTuTZmVyqATHPtK64wfC9r4skc+/mUOehcVM52LUMxdZhzoMoOR+IjRwEBrriHsDSy3WCXm
TdFhPycLPLRZf6L14lvJDc5qi8mgj86GNLvsXCqfAUVrtwPYazRELtPGujxfXeph0t0z3CHgKIzb
ufdP+y7nWBwbtYEQcVC/6rfjgY5NHWbe7J3tKy6eTwtC1zjtgWybSJysQxbYWrY+OwHeQ7g1mnYK
YA9i5fDyXz7TZxxBBwujHvINrqEURlyD1fXMeE7F7whCqO1qRx88lAMjSOOokkI9JfDmEXyX8qoC
gzsNcKbiEJl9naj6sD49zBlaqWbb5zg2q7nn4vsSIIt6ZXoV2KE3fWC9J3LFJt2e5sLapcOhDFju
C35lSNn1p0yJkLrThdVa3+4CRZlebw2+VeRHV14DhvTa1wyAERotG3mwtxCSodWxCBp3NdOGWkUY
IplH+W3sAKGOxmduEI7lD/j7Tx8cTK4o/kytLyJWgM6Omf+7DkTQYPOFoFN9CibAOZG05Nawmqps
69/HDKhZK2ua8ieKt/3WBFNBkGm8S3SXB3BWGoueU7vMdwgh2pEkcCoMFXBo5kbRczKT7JQZMrxn
bohMNKVRT1zVpuc2uId6MTs1CNhtrR0RX4dsxYBXHOr4TSjI2sVc1Li4R+EyUfWwfkhRk83dMeZw
7t4xzjqWNqwvDzkjMjOhnNi9ZWhk/ssYvcBzSm8boVK7TjIgN5HVKt5eszFpRGXGj7AU3eczeaIA
tf4MkxkXcqod+Pl/sFkg/2dPmb+YBpZxZvER42zz+9ssOt7R9XRm57JINH8RWKNraIAJRk5F1lwC
WMT2+dR96h7g9dp7gxZOJo7JHxVGSVuNhSZAB0Qy/b45rBaRDABQQJBY2y2pdmRRQCrs3zH16SfX
ROOafXAKE5yGl+QAWKbzwvXRlZmWuDm+0Dp4dXDtWcoaXi8IynN1TNWUbM/kkcLzuw4BraIJKr4p
pubmB0P4zVvRFjYj0OiAdTW48yWiaRjYvJU72AVfXxcKVlCALjphCdMwFq2XN3q6EuYuq1vX0BbM
9kH1mrP8hCCQpsjYA8fSKrM0RxWhe5hnlLxjuvezX5kZyd+9W5hc1j0B+mDJBYAu6x+IvzrWx77V
kuFNcGUJ2eNoMr+Nr+kT0tq/PH7MMBlkMN+LdrF1gPszpWxyhRvL+A4hFN1MTUX6d3AB2rDU3gz+
Cg3zvZS36BNlwal+CO5JVuoAFkNtFLOAHrrtG3LPcZKkta1Lbb7Fl8reWFxUcQoQVTvufGSUoifV
6DEBB2ZRNsVScMBHeFTgoxAa8S6Rb9nF7ojdlKWbbkNRWEeJUH6A3txZogCqBtvL693p6AqsulFa
4TY5kRbuKdJ3bQoA+LOQsuKlJtj7xWOMCSQWY8C65TpM0km27uDh82ik9nmXFo9r3dT04bVf3WZt
o0gn46YdB+q9aXgglkMkMP7buwx/Cjr3/mTCePJWL2m69e1H/3A5Dd5akQZMqs9aWxTU+3BVCN/n
6FSjet+AqJkihtvu+WDjNH0CD2iGKpCNWlr3sQSQYwAsu/Imck2CyZRyUqFa1IxXus9sMhyxg0+h
TA0BAcr2k/y6Y/GHiHcR9fQNEqtiPHFKbZQXSwzcyNoqzu9OIXEP8DKelfR69xIoEU8DmX4BLTCk
rfSF2KWb3KIjGZh36TNt8aAN47+HPpHg+gPlj7nRAcHjISArPmClv4EXsiVkulGaT0wtWZVsjEi1
zBrnfRdZnDxoiTKWPyaTQMgHEsWLBx1pzNi+LdU9rni7vu2lRo90nGzTIVBlzqED3Afe1DsYgDyv
KFM4LTFlzN/BJYk7kJL2zGdvv6W1cCWczIS2JxINjrMwr/X2JwLUg/vmK5EXO0wgx0M5GFXGJqIC
I/Dx2F1+betB0yHn138GpUlB1lUqw7g2G+Q31NT48llPsiGQxEiU2bTBLdfrVkOo5eDSOtKOwR90
42MJgV4OQCAVtjjgWU/rU2qqtmmsNp7bIUlIJKOvF0jq7mdC69jRV+aRqJzwR8VeyXkeDbFJoUMj
J28TJ5QSh9wrfkQrW3LUE27l1MZLwSA+ZVS7cO8Hembygq8tmzWvJ3CTs0SDTluF1WvQmJWpryBW
GBrSIlcGWHx1/ui4eIeI6nAru9LOEvfQtVAoIo4/fRMIUajWhEk7Yz/SLYvJ6wuR7gC9pWK7XM9n
oGck+0NPqSUAPcywS676shT/ATCyBVYsibESOmFXVOxlHqgakG/xx4u3EdxieUEXzUcb72SZ2LgF
u1WGZ3daucqyoSZxDA2UhEmBlfNlfQQsiO8GHwkwiQNHHNqPN/IOyk0tyhOnsZp1jFBSWhC3jsZ2
uRnk3MEpZ7BI6V0sVd9wAM3932aNR4OjDB5zRCjGTsQ7HhDCcKDPBooOed5Ki3n0cm6mob9BFg3d
DBoIWL28mFRa47fNHzMXHCsdimIpueTGOoCdWZQ/bWo12Y06cn8z89Mw6Z11zfTvRoYizqNm+wCO
3TRTAAk8UN/HN2JX/Fkt/79M9NOvE6VxiLWpcYe1MnEow2feLd6zbrmfyHnoFY5/YgLnRjY3kGvJ
lN4jrnpBLRwySASFQoBBmQyi83tn8Ems0UDU6RQ6fXYmIKasLyrCanoO/8EsS2Dlgv9rYAkOjTRE
TLkCURh8ucDxGgbN2wvKWrSewVLMowzsSEN7uTESdDKLEbJnispQyYxhbBHTgRmwBUSpBY98M61A
9YPOeqBxrEsMfXEzBWhRS5kW0IeCwd2B1nNOQTYFKqW/cdpamMnGiZbsYfXf2X21MG2guqEW1vxS
C6DOLxro+HvN4Vtg2WvjeNFgEtOEMPW6/t8lJyCPCmhB/eG3N7cGEa91E4XBG6eX+7dLm5q3c1vk
HjRIxageNhCdhnKhScOOX9uM5GJslr+UQ33UAHXTABYlW/6zM+S+OtjYCCESbXSkVNUbd+NRHKdZ
Q8vbA6SKPKPOhNia74R7BJ0/sxLZ54nqD2UIEKCN/ShcT+Oa4zEglZf/yxnarGbqh6h4eO1cTVbV
NJBcFyDZ76Aa5Jj5a48TsG0frCtp5ru9/mrA70abbEvPWFeVH3w6srRGjSw0QIlJN8haXSOqSaTF
JhFWIEI3ZNiy7gloN23Yr0gN4+Sf9Pg3BDK/j5VpApm+nTIU3xwKoK8wHvi4MDFLDCTqeiLJZz+p
WPZoFhND//AZAmeCeINZ661/bs/cbZkBxdol8mHXSnYpyfaO5S2RJ0dLXMRWdyy0ephnDeURZjDD
b3SYD+bYc0k17QG2rSkCMXwBqjlpg6z/uO/m4RKBcsGHMFuPtBU3DoLbyCmxIeyat8QzqSJ8BayL
ttC/2raHxTpwoWFvHFcrCFcN4Z7d0N9vUcyJBF5FNXAeWxuZ8IeLhYUZ6AeSDcQerrdzArt806by
3XI6n/TT6jySUSD2YnizYByQAsBp7oi1IMmveWs6DkFV8ir91nmNYHa5AgwvR7xuMnBNBCpgFOaz
KHNDmpghr8eZeBR0DCDOwcXmPdjLFyZKPSCLNAG9URzbDZwGn72h9jt3scKukRgRO6jk5yKxcFFq
pzeYHkT1MF+oVstLZ9Nan7zl+72O1ciAJ3q0GSFAUqut9q9AB3C7VsvSw3V9vTL6iaYngx6HHArA
jYPSRsVsD1iB/0+wLhOLB2NTyuNDRC2Yil79wDCTK30OVBBs9xFWzpUqJMDCOaxP07dWYyisJhDk
9dmDRFfxuYPzR0xxb5H4HddLlW+2KsWIC73X0ANG9wHMfB82eGWIeAnjrI0MKNhp0sNwDjPuGUs1
d8bCudMX7w9fJKP6Nrpdwd/HtrGxHxvsQgNPha45SiHnh+ku73h4JQ0BEt3YQ9hsC/V+OHEl1hfQ
aO26bXL9VlVpObTU5oFjv9dpv4AvcSUVvWL1csoWO9LYZ1WgmKulAyJ/Y5BfBY5ppXgGOBRAINDg
/Ol1yGFKTExFGt7HMz5QUWFtQF84EaD80zx0ze52nzAwihxBcnVqbFKQmP13g+9JllesHo/TiHiu
0Owry9ytCrz06tOtfC/noIaoUebm149euR7masUMNgipilsJ1M36KPbIbQuV0MJOURZ6eUQEUUB8
qwak/nk87GKh1VIYCBDVO2VrYFenw/MzDkNgGOKYYRGyCwdiNCHEKVsoLexRZFQBro/ZqEiN1svH
Z9lVBhQuo7IQpcX0IkS3p5Mc64oNotZl4H3K1opG+dEGmW0ycEiqEISivoU8CwJYfPrLOD2LdR39
LTzUNnHhj3I2TTqHD6u48bYErkF755luMggFkMP1Vasr374qjFfoHWkbXk9zh5/p0JYEsdoKRLzN
7pRelE7nijcId/ucGgdKnY4S8HAvOhlPt3XkPoKJXNvKSmUcFgRlS7E/8wS7z41sAq8uj6I24aUS
tGiOiQX7vpoSYuEsvWvQ5ZX84GBiSRPH/GV3XhAahqjcS8bE1IxtbIvHDx5QBM+ODKVGxi96CxKL
NMreSSw5vjtDu8iBSCRzNAW89tW2V6E9PFPHZdkH4MvI1V2R0hGN3S4kgD8PA7Vu0aAjSD5CscRP
5Efd+rRtmRg7aryup9hHjwYQ46b9+hyGfkh6FVPiEctSF539RBZAITR3EpAnHFzeK7eNfExiYft8
Kr+QyAtxxSowrLyeZ46tOOk5mFm5GK8Xca2EP4RbhwwPJvwutTMuNSHKwJ1xlAuKo4f3MbUYIN5B
jbAYS2LqeAbVeMJbH3fz9UTKlZwZWmP8VIOf/Q4xl9w5uO+gBRIZmXIOzbfnhnhq2a4OxE58js1G
SlYZZYv6lP4pF5QnWV+UgU+xv1yb6iGJgwbWUafn528/JgCiSOKBWBRKoFgCU9ixoFGqu1gcPCNo
jukm/nkxG1IwjEY8rtffvGAmptgWzd299U7IG/YdPlGt7ugtl6d8XeDbmH1ALZX84mJYUG5N2R8b
YRZ9WUdvkg49Xkgdrg/uQ90jl2oALJHLRDYA7lh79+ae1yMfHY8uv6AESD7H6NGDdH4RY+Y54p6m
ZSd3x1VmBHsQvqay4p+LjbQ3eLl/HX3HS/61muzjl5clIfQxv1sw84CJNc7J7g/uPu11sMqEUn9i
NcAbSnjqWWmvRF78s/PgvxpfGaZzjnaWq3g6yFtm0Hpj2F45RUzPXs/IwnhQOA8IsxkgnYAORLeV
pCX7Z0Ly78BVQpFMQT4/fBFD/zvxkLiIgWiWcR4zLx8zPL8ng7qbBCOdlTizmoWZXGvVl9Ik4/4m
WeWsuI8O2L4LmaEdcUQN40nhuayXULt0OdmWO6Qc984512WZd5EheZfjEh2ReowyB6RdCBxliJ2Q
KWImcDdqHOdCcY4ckX/MlIQ7r/Vo8bEl+8vNnMEp30HuEk7d3VNMoUj22fQPwED9JlGk2mXHwvv2
n716C8yJG3RSBTaAG/VwUSJiCLnOrkf1Aw5tumSpvf63YLf56UrHmfZ+CoopSXd8SSNr0WWUKVi/
3gwHQ1raTIN5STzsnvDF9RpeCKxvm40B2+bhaY7ACsNi1EU/dJA3d0zRmZQvD2LHoEFMB8Bkq7O7
T7nGDt3suqBeo8Ix5Np/v9Stu5ALklzsvwp31JwnfXOvAspt43owlN9X4pfaXy/D8PBOrRf7sK35
nyU6XOF0wh92Haf+Cnj8T9jc0O9g8aehTnzJENk+KtMi0EBISD4Wt0F8pHZFVdr5HUtmuF7DjTtC
KzClI+FCXB+OqwsoXPmXbT8xdv0cIYKOFG3odwt3Y3iR27Yca7zpbrKzghgYiEGy8gt2f7gjvbLc
7fcz6rvKe37amXcx2ffbHPm7dvvYH/R/iAzUTPZKni8QYitlWLATArv++RzCrpwsr62IC6uA4oH1
+JHeqQfrfWfMhReqtgPctxebuV7hRSFPNhqLKLBCtU2WM91cC9OrpvyfKGrFr+FmS+ZMbxV7mJyO
Hej+mWw+FAaKKMqRHYASmdevYtxXKj6P9c9O0E6sFcjKLYuW9JW+fT83ySrub44B9bKnWpqesDuA
Y1P01CaYmjADcMfveZIvPWWQS7kij01nb9sVwYlgm96GkIpIEuVYzB3CGpzkZ/pa6ePNIos+D2bm
Ig9xed64bgIcBLtHd+83nnLSuG3sEcoyT4K67oqckT4kJPoWRHRsf0ueobTL4uHiiJYjchtVbSVQ
WBwLqSZLVyCRE+oOn055OHpEOgSW/l6RDRTZLcWe6f0SLYTdriRHS11ucVmvCMrxxVoFssa/Nrhv
8rLdkaF86YApYkA1Ltde0/GXEcgHcFqscSsmhjbjt12rKqWPHzNN2gz52ma+TFV8t7DWzp22mAlZ
uOd/lpJpkb6URjzSRNm1RmPFREgvO5gIjTjoi+ACwLH7Atsj1QJEDLX++cN9amr1HHGYXWkJGPgC
neC2aEltnu7zVfBNnHBcAbn1Uz6a/qxTKRXLMF6xYJbsXqVx5mLp8e3/EmKc00Dql35moW5oiI4o
KB+rIEWUmbeWKY2uq4kfjJ+/18Qlc/Ch1lpC66fvfyUkQmdz+OsYpbs7a6GY9jhzh4ygsDHXI5zV
6HfccOWcDmG+h2SJ8nfMmqYcUTZCXlx8L5dPZL5bMAmnCIpeFgnL2V0+U5rsXu3beFVurZOW2hkh
Rg6V6BmMH5Q5U1IUNoryNOaCk3Ew4D78n6AsbcC+nGzweSfWqv8S1LhJIYuzUN3Rhp8851nHCDup
9D+95tTU8vuzLY2bQwCdWrBRSbS7nAOmGTyH61arlO7YVQD365Vl3RO7a9HP1GRs4mU4S7vDyTJ+
KZIfIxECSEzXbOsVKOOq5T+KhU0vFm13qgHBaLwktAO8bdD/RhhSjrcI+KpnzhiOeC6vr7ULHPtC
nbUPpr4LVVtco2ElprIepzgQLoL95fRv0QqMJH5A+59JRw6Bcd+1Ndmmq+W8eqvAn64iBNzRILCk
nuvXzyTXaKW8l+5Taja0RqhoCHQfYlR230KCTAw1s0TXhdtncbq9tAiNGxpj7vAVznIpXaOqQaY6
Ndf9wH/PvWK4Q1BYfVpww3hFMKudX90uPQeeUSw5qtRTfKIx40wQ1sEJ3ZGivMLzJ+ue/z42/Wsp
euI9vI5rL5Z3d3TiwUMC/PzkMyyzhmNGypCffSn/XoBJzQRolXGlwmAUvf8J7dQe1HFyllNDBZzL
nrnomaF1HpL6L2/2unCBnesyrdWVUsdeKNtRTP9Pp3UUj6M8qG95gc3/N7olHv1ecJiV1alQXzpq
l0zJ/AVmklx6AEMPT2URVf++BcRb28eyuO8TQxZrAdbLjD/30EJHPDKCwsbvR8FGTO/Vef3AAxak
WSD6LK2PyM2I9OmOZpD6dEXEl7Y966yg6MaxoVHKmVYa8Zjqu0iJ1RzI/8d/JcBjuyDHRoP/uDch
gyF700wlile2jtb2KHvVRlMeFS591EWtXpdPDQMrWMFpKOHwFFZ1ZO8bs0EHh3n6vctFLw5mcAxb
x5zxurQPApwHXFnBi4DzL5BSRWspd1gvgNUJW/JlZFKp5fIc2aLzcxoQVR4+cGKmTLwjSk4IJRRZ
EpQWH1BOuCVExI6rxCghaBO7w8MuHNYBm7L3Mdi8idWcRT9/O2TvSTkdGTdnLYGK9amOcwLfxFF8
ZQUziYuvu2v4wT2lmb6R8ueiaW8rzWUbiduKbSg+wgpW38/7pI5Ie2ae9kFXnL9ZfYkEtGX47mEL
j8o5xL4MrvqrUrXmISq/Ob/YhgGM9LoZ3fgqEGbWF1SuRM/K5kSHuoQTTaOeyrLPguP1FMgkC8e6
k/IfveDZ7ApyaxqBi0sBfB8HRtF3DbPFdXJoZpi57h8rZIRzUXpttGh9r8pZJBifIJHymUD+OTBf
7U03Uti/03tBkpgTw9dBnvQiODpyvs3r705gsv7VjnFzIn0A2zscEAOQRPYCAcq+PCoTn4afKeow
uYuvZBeyY8l3kuXoWA0OmOVuvfQpSHMMbaGy09J5+2tmAmGFPggM4AxmDQHUTPCxPtW2i0P5QMwk
YW/uk6U/KaHJXq0+ntQKCiQhqO7wAQW1XfrAr9n+1zBQRoNH/u+qImxqah7NheKXp/PYghClL0dh
xxs0n1PIbOpRULIduWFarnanzs/Ihc1BR3au+yCLQ/feuKI8ZORtjyOIuHQWv/dJBnkTxmSe52Id
RcA9ADMOPRhAZHJAAa/uRp++FGNkZI8MYAVdDVkc2sX5R54iyfUAFsIjhhp/gE/w2ZkT/zw+/QKx
rx+PR30IoDDMDPlFaz6roZ7S2EaSDgvaDXmtGEm93fY+7ykd662BxDdMYzpfUtdi3R/9p63l/XCL
l5Ag4jAQQUjRfqYArh6J9d+a7raFteoq/9TkHkd8RHdMW+pCc9h2uMAoiBcSjH4Yage0NSlFSkdL
D2CttWqLv+ncFoB2+xnKSQ9kMJg9mbOr8lpts1tnCUTxiKeJ3F1i7TNVLV9cAC/T/v1grFHVOVUU
Y6LwPkJbDVkHNhtyPn9B6WP9g0jxsujkoHd6Cmv8asr09R62bzFKgg2slD3kpgd7QCAlBgspw9s6
PtOxO+04Te5CMRv1AP78nLMp1i85cmgTapvsaim+njrQzAUVtzAiBhmqeRROzu1BQpc9iwM4q1Q1
J9heDliZK/oDSsX3hIG42OgdOUFn0zudroJSqEMqucWyYP1ZbJOhA43ACk5IH48N/Oiedh3AEmt/
iH1Ugf6xxfdj4VJbRt9oxTq1n7UAS3C4KGUJh2zvcARqLmq7bNpqVMDJYLU1bgIVS09FWpq59YDy
FRWQZMhnZFwJjh1cZbxHcYpF0gPrrfIHaj7g9TYaPVA/0cItU0qnxrQYKEGBsh4LL5o7igjd5Ahz
po4ierOMpkU3JWCdfDk231enH9KXsmVA6x+lkKSt5LlQBp310rl52E51mOOllnMhyCGgV9eu1HdD
T1qtmCcHzcg6qfmuUFZtOFJlPusAqUdhBua6Y3wv6RA1l89DAmQ1USMOHu1tcb/k/QCtxR6pyNLg
kwx3i5fyv8eAjkhJ5aBbFZvpImZVj14chQCxGw7Pnw0IOlsYQsG4ldoy2jXYzWNwGwLmOvu3XZao
Ia77hvbBTH+YmQBPiNLhUMbnvbG4IW3xEFL9+KlS7s+LklF8tc5OiyIPRIUJ1f2k/0sI5N6mi8mt
NJGMt1x3Fm07v4QmI0H4jEvwOLYFUMnPh3goua26qoaCQ0HhrVWb3cFtRyZGB7qWg8f41UtRkZIn
bPa1/ivm+qNgPWsRL25xQMPbD8n4UEtedOSu/mQ8y6ZUceVmHwjU7V/5oz3jC082MZReC532lvVj
gqB3LtiakllRe7DHIPwmdvP++EDwvHBObBrdJ71Cyg+7LUQEQP98jG1HM/bU0tECmH08/7k7bXGf
gwffPt700FBH+OhS1Y3NPs9ajSgkiOlfpy+4V3VoXi4AT805H9kPeOACSYb1Os+kdxv2Zh0K2paO
RWEGtnFV+Eweawa1CWAAvD0+0ZbgoM1/qOfNJCnxctXNqDUutxGaSwPn2vkzGzPyf+8/CCw+M+BW
QKTgGMS8Md4A/WuzdFA/NOYiR0Vx+XNiDTDOemneed2I0YNFJ3YT7C2C5jHzxDVj8Da53+sUoVkV
ZncRkT+8JHLsZ8RTEg2x2H/rSxjJp+ffAn4xebkryU84DuDBR6APgryXgDaL6LBg0phMWlTEbodP
HFxs8f2IOwQL41jhDNHyMFmzxt/dNdhRCsG8EVvEvCEW+cSjKP4UvxQHsMr4pG6j2ypuoDA2r1iv
geiQuGA7/8lGAOv3QOCOfhXM5DXvsLWjrwkV1RNdx+3mReI0cujK0Kt4LbdDwYfGqWKhvQI08LXa
32Jg0kHS85f0PIuqEzojmu5s21OHlCDPdg1P8FHj4mtVyueiF65nPG+in0U7G/7cnAoo69tgTEG1
9sDGo6Zk9rTPyiLTyhMxQ7XGop8kbTvGkNP5QJKIlK3YPWM86RlLGxx0EDz4rURbew6EoR+v5Ahz
qNFImcBk0GhwGklGGUd+qwmsHQtH7Z9bRz6aea0VpohzST/5sabs4qt78Px7N4wYT++amsrGR99Q
ysS3Cy1SBrLv4j1uUuEsE2snenY88+SPL0HSgYKHN69PlQmJzupm5eDiMDxhLObtGEeslPETQ292
xltbVSdHKlny7OLuRYeTJf2DkLUdkJX88+EtoSMLzwOCQGbaDwHqzyVFzw2VOaBS5VI4vRYVUfZK
03w6f3dzxigskJWSOYMjuJnJIphusTMKt8LveeK/TzcR2bWKK8aoFbdyBlPAoM/Pds4/bpaWHAzR
40dxTwS19tPmRbOjeR83qpvg9ouL5KEoAcDMmOApiV4eFfAhySyEwUW7RYT5hovRY1YIcUZaq3no
CwyB//bWULUcwOB3lvcF4i7LnlkkcfYFnUz9WMS1lAcNooKFF4H5FGda1G7DHWKX+Q3mMgCvP5vd
WLmA4opuTaMW4iVA1hdLCMswTUnGZXrjswt8bN94qkkwAETnqlHXe3RSaS7XQPKqvCqLN7WhlPie
DouktUIoigkqm9a2U+QmzZP2Cz1/oY6EyhZVtQh5j7ZKi6rEB4zNt8U4GrogVQgo+55qCmxUNmuT
qd4TAqBCTx7zTqTM5XmBnAKu8fy8lI141zY2jH/IX6+iUX94iBBnuYKfosEPxXfwzmG2BSv4ArtY
7Pu3nkh68LiepzCSbdYQMZamuNOHLxSGT6YPEHdDCNkFh8PuASYpJF0MWdonom4m2MN92mYg0JH+
FDg0QOxjQN0/g+A0pdeIp+mLQZvsbpzDOgXFGG72Q0LFHVkyjHlyMs/r4xSDN70MsyxbszN7aeMD
FKkcmr0BEbFDXMYvfFh6xD9BoiwCMoGc60o/OFJt1LmwBbYIq7oRVnQgE2foi8GXgE2jLCBmPNDz
8Gp2SJ4dxBfgDz6Vv3WcC/ZsOTWKUQWPNgzdOL8mzcV1dCyWhqIYmY7cTYp8YfQxT20R19prw2yU
tvwfgZhdntpPK4/xxaozOLfp7DPNyoWUdUH+Qxpcsxu755azaufwA2rCr1oQENyVZ9oO26afr2CC
r8soGu9oyhsO3tHqRvReL5GEcmmQ9DlxYb8zZTLO29OGQo/39RxrxAfQoBRhnf51T4nd/Y0dFIxn
NJTQJTcNP71ZsXi3aeiwoQglJjK37bawHPKjSWMVJjXWI6VV4H9lb9823IIZwu8ZJnLRraJKYGG0
+JDNp2tpmhjdzl35h97E7+mFwKu/Fm8YQiS1ZB+nwVBGNqPlIBpwQNlOcUPauyq4Fug1YcOPuht/
9iQWYeL2w7YQ6tO7Mc3DFitngCSNLVXDDQN2+AZgn+db2l434vti/1DB2l8KKG9d9iiJalZPxhsi
t79fzVBwnzsfcr5ScDuVvVI3lLxTfPHXfU6fI+QomoJhOoHTAgAB2RORXjboiMNfZaKBgd8uAmy1
00OR6+6OXlRMsQLdFl4rdACHuXc5SeE2Cetc6K+Cr86kzrnanloc+Z1BxNqEHIPDcUIzjzGpMu6v
pGcdolnTlQ1dENNy+L66pLDW/jTT1huHwZFMQUkH5JoasEzmCkgWH6ass5RrUqmINkRycVlJttN2
VZUjKOLU4I7Zg7ryDenfPbHUyXerq5MFE3X/mRAWTYAnzN/g3c1loK2Lo4rlrBZaLLMBvxqw4WfH
HOfls5hNSF/36JTNssjKYKK6bn+jJra6Cs0RV2F8HQGws5MAJGetNg4We9DtAdamVL5Ji42X2aBK
BnOFkgtcgOZ6QBqBRj34gH6CiGE3ea2+ORn6AGxj7zzNY0keyUa6+hmsjhUoYZy6i3s5+ruap9Cj
uJOiiEYkn+cIsICkZOEWht6ei5Y2a6D8UcscoZBglkZST68wbJEA9bm4UodWesUTZR0pW+FQDGdW
L1i8vVocr2IBaxKAw0f5/y/lYztwjjB8UfHOw8EGNLZWLBJ4lrcQu4YPtCKIaaTPiwTmcYJvq/5F
fQYiAsP7MuU5zQjFnDIwJUaHkbsGg7fFaZyJ3JdZ/2rGVdZfp3N26kcILHgqt/VfRedgRK8pcZnf
bCHAf4Qi4uOUNBtZ2F+AeB4k9bfEGqPvrA5sM4ETSIYjCsPOhkGW2lJD94eCz9L4fJM/X62n/yFd
9CJsCMJl/EF5UTk1eLP5fOwRUdfDc/LI/RhlWAFtDTo5y4IvONibPT46OJeoO3FBjVPVdocaHSiT
8wAXzhII1yg5JLGhtpqN3K5OPnIRCZAyGhQJCWMpqMuURfNRyAVoPgcyeBag8H7EZy4+TZwVCLDM
xy4+Axzr77KsXu/K+dq7ywC6vW6WBMBMgM/uSmNk7cBxRr9hzR1HTcov5BPpIHyl4GFo28gnfVjJ
Iz8ZLryn0MTAK8Z849TYAwcp6bS8iNoIrF2Dd6qnNdZVlXEFzarZucOu84mjcO1Xp93CDaa7T4FL
1lWKgg6oJc71Q4jlMuNQzWvGuwCYQ1NwP2GB5PgXzm/w9xd86oqk3l8WdXAPEqTpz5gMyVVtRhZE
irCePBLtsq3We+Dj48UVYGFaIJLlOchiAHvDnEt4bbDMHf7797xvUp1PJHOPEy5J/9XTaaSGuWuJ
8EotCZPlZ07DX6X/sAETmdXGfabEZYL6okeySioKB6tL7BC9tXwSSPFYADIo76tF1CFxAGB5wR+h
5/gMmeM7sT2Aed1/0KPvmjW67w63UUGuiY5xZKmdrusHP9nOL6Gm/2b3p4Pkhkbq8gYyOic7J3SD
WCpRh/9dcOIEmhbhqWiOZeO+/sa+X4wOCuZGgNVNe0tGb7A81ZDzZbCQDG6gmRXX5jysACZL2wIx
ehR7T5jLnx0SNTrfTQw1OJex/hEp6CFy//H6LazasxKxCCAL+uPTzi80nPiICOMMtu2Mp83VUn4w
XD00uMbD4QhNh6mAAoRronv5d1D9ywTYwIClxw85RM4pDsuUE09qZdJATaNk+Kf4AkEr+gPmqxdp
0+p2/Nt/o4Ktf4XcwY5Y+zgFEqrWMko71Gu/YMsxlmmQq+pupjMebQ187AEqYmD8Yzim2atffNFm
i5RPiD0UTDcnhujNDvoXK4QtrZqksB6efY+RZWb9GbWYhfkVKvkI9hBnVtFvmfWNf3baU8voBQuo
pvTqe2ZqlboCBYECP3N/QJUlxzZAx3VPAXStstMDKYU3/9cV0EiiDLq0WUqoVQ9JwlR+iHDrnZr5
nwpRxitvHGmUPmPXs70E69Tt5nL5mJ/4Yd/4FmAg6clXBr1Ypb+k4bWF/+ifpD2vmZCieTP2Dzg4
Z9ogRpKTSLiZUkdlMkiCzmBqt7VZnfxNcYcsTIjOShSCCnrOwS4TVjEQ7RIHe68xfdTlMZwHG+Qv
rEd/M1hXXSACMndaruf2S1YFfClgCiXIm58W9pM5Ji/PUtpfNai3//vXVmIG8M1Z0IyazEvPurtx
y1uYdHgdHF94qI6J+5b29Te1VdczlHbaUeIz8gHt5NHgSHBR65yUQ8ZsS5ktrv9Bh+CG7Ozi4KsG
T4r/n4jfxwaaGVTW2o7vyn+0xXO06TjOsxK2lcKVVceF8RUcefDLl397fmeiwb0qn+Ob/YJzKYjl
dMggmcYqSFiLB6IF52pn6Hrh1rWmtno9xuMljc3y6GO/Hnt6ut4Lib5FfeaJ3lNbtuS7d6c4dZfy
FuTcLO/9N9bPO+wvobz5o/ta5PZfZ2jFwC7dVYED7Z8AAi8ZeOecMJO6Cr9fUHFhfFHHPk53PlmF
5mMLA/KvjVarvC4B4d9nEC1E+oeUOcnD5B+3NQN15fyhWy1lDfob+npgh50DmOK4aECftd6vjKjk
XI0UHSZ1Z9AQdVh7wjfIxSd0etg1Z/hpLqX/BsosrBnad90e5rlNi7po+i0xo3QMxyYSkAgiFOM3
L/yNJUQ0gnERzddgk7rwmWdW+OsS3QVX7n/kFiBygaK12PFJRU5PB64L2Gne2q6STCCWnHriyoR9
BGhXZiTWAc3QNloWfTB9L/D7ySjc3X+MZmgreV/AqO94KgXemZodccWglg4JzXUFQjuUpkX2b8yH
yr1KX6cEfsZtYGRMZd9r1iIEhiI1GNweW3rE3roCO/gv/PInVetpPyeW4QK2wWjHHkjRwpwAtnxK
ivzZJe0TT8bL0TxcvX7OMag2CbyTF2/VU9cMznSXM3G6fxlLfsZ/rivnqXih5NPyrm1+lFwPcH6+
1NH13KfAtn9PxJnMUWx1fLIznHZOOWpObu8xL1UpjBUQDlNaVgTqRRopRb7XnSZK1IUpkFR5Qfqz
xvYI45bWosiZRqeB/ItnTVDjfNZhWXD5HBvioJAeSt6X1mgn5xdHZYlakuciVWn+QVEeYknz89wc
YqkFi2SvsnvZK/IR2duSUh3E+fuV4iK6uB5T7HL02RRP6LXWlJjbvYg9pdkIIHm9x8TX09r5Tm/k
tGyvCPzaeeYgYNnZAVcy1Ti24ZsVb6s15BTDMyyFu0Rh9mRH6+xAHzqrv7veSv39svSd2HZZ297B
2QSbWhNuy8v3cQDsm0qaLgDFQY1WDgPhhda2Si/L3p1o5Y4r368kP6AZ0Dun4D8Y53qq30WacI4f
1MOFTFuhOf+2ngz/r36XUTCojam722mmBo7/K9Bu0nD9stDETPggvxdVnQ5b107vaMEm1/wE9cQ8
4JVvhFV6W0k/WKdupo7rpI+bGKE9+0xp7kH31A7j2fq/4uQbxn7DP4eitXR9Lnsup0NxrO7103gj
Umyki3F3aHGgdxroNcWtoWLw6yThfdzgqS+yClGCQ1tC92I0CGvzvb1JZTXyhC9hLOz1xhUOyZsp
OTx5dsZCBq3IhjTKIZB31spO6M2kvS57kTinSAf3g0/hERjQdfTKxr01V51cZSYV3trW4WV/5kDh
ZCAyNYK+kVuWTf8PjP7GoFeR/jd+Ai6iks7gq6+aiEfXpVYYKisJ7Mt1Lfo6exc6XL5AMkSuQInP
geulvghdM3Vk57S5NmQqj61Jw1590DlduKFUTmfVjQ5pwmHmkLEJFeOlQk0CXfA275D1XmZJ3l8p
qCebTM/kUGhKcDB6pcV1vQZEnxHkqASe81Q8RTKRRavui5UDsKbPb32Oqik3yaLFPKvUkS2mDOlN
QqzSH47pr0a5ve/yp8z/kwdsE5hOz/gWStDxOdNuxPs4Qi4zzlzfcSMrDJBAM+dOAOIZ8Hs6GVMo
2WeRzTSJDHy1Mg1dOQ1U8PDAISXypKAS0svh1qGTEPORNPqD7k4kyhw2t/jNrZ1nkbUWcdRoMH0C
wcE5ZkBaVbyFxmy2hhAfL8X3k783cT9+U9RWf9Qbsw8UehEkEfsEXvvxrfLbbSfxjybBWvF1ZKHg
qCBZ7J3+Rfvd7MGt4/xxbucJt/sSiGCyi6IM3mZqdJY6Zbg3iAYojnex0kV1fI8evzUJwFempL/t
lLLuGyh+x/9m1potenFbqeLm0s4hn1p5n+jiEHDVO2Ovvez6fflb2Y2o3xsxni8ESTPaYkZfa89e
YHD76ojuM+iszG6+1bQiXH638wiYBt667m0DuOja5v9G4WMp4yQpeAYqLDbQ0By+HteaEZ2T9rWq
WnGGvqJwz/ZgeRZmwb858XkUC4Cvom1TSiVfGh/C/9lEby9dj/NrlozmQRoTrmkzKXdxXky6bkc2
D3ej1RBhYjAwuhnnMMTMWDZuEx1Hg+/8r+7FWXPi+9IM4NF32417ZS3TQ/yoVvd5Af4KHlWc2nFS
kT2DKW2dUtFW0PAKh1b6JjBcazawMKZOFOeiVZ3v5ncF672gBIUM2UR+L0wcjGoeR5tS0nA5g06c
WV1Q/UtjSUFtefLJZDpli3dFRj9p2TNygtPltJ/8BgfWQXDfyAydkBuoRbJZvRTdyM853AeQ5QeB
qsa+Uj87Kgq68V11l0Zn9rkFz1wWHHk9zra6RlEWRK2CA2LXalpfkg039yH0DekdKfHyiQWG9kJx
ZDzUOSDcSKjd5l05Lo4EqshTkToUNp478ImtyG1PEIklochid1y4HTmiPBMsrIa7FYeYvi/qV+4j
M30p7+7lnJhoPF1KTX8+0JUGHS5+IE2yOzirajeU4pvmNS1a7HPX8F2y0829LA6c1bF0x3BQCXzq
eCyA605Rc8uUWfdp/GSQLMQPTwR8H361xAdxw5hfDRY6KCrepvdZY8Bu1gg5IkRgd9izMEpgKhZ1
ZO1D/3tYwTTxF7v6UXoho+b9hRJC/RKa8cYlAMJ+3Lasl95DVe6i9o774VJ6CQW+2gQBfGXMP0eP
xfpARs5nqmKu65qhfEfiKTc/GkmvxZvEdi5lXH49Prgy9BSeUxrAodCDhubjLTJkWKak/3Wdywdv
BT8S68izTBVItTA0pXksOLgsv7UI4Q22xRwTNWa5uwC1wWDPiuka/FpghnAFvok2czxfUuSe7wsC
0UvBKBBWk9PLF64zx5wKeAHMM34HBa8iV+WLe/G0xA6/Rx+fIdUZMz8ZfZEGPFl1H2XPmtn/SpgS
cXpmV6MrzhaGxVB7vBpJT/weDX1eaJUZFy0AzBMOLSmtAUsAkgWm+oL8IOf73qnTE6TZ+v6MHQzk
Dlzww5i34KyRdcFsRcJvQmfdIdfSnu0keF6cxZl2SMuXfiA/Isvih4qCKh/s1KiqSYIHmRBJxvjn
CDxs5Fj4chEwUJZOVy3O9aZfaKGlvgBQ0XEt6U1fLi0JCYlznKSWs8/mlgmCpFLFIIxLfFpPzLcW
svaKPdOb5MQXfU+lvrPUV597GBYIpblqM7SbDgJM8ZQE+jUPACMPnHAFujt3d7FR45GaknxmDU+K
WO3CMALqoyMPBwcKtiR/kcdG8Mjb5lt0L4sMeDnJRUZe95b6pXHYU2QOmUSQITAihF9GCDS78T5w
unl57AjpihzBH8K1GZW15K/HQsXMi2/vPeq7cgIvO803j3gBtaseMZN2mcGWdCuPLkmxvWhKQ7vO
xbaaheW3dWUQ1Uc57m6v6fD8VSC6B+nm052xNEMVJkIoeY8CdN1fBVrWyBSfC5U8EcLJRHBL//gH
Y1VL92IX/2+P4KSgZgjBocYaaD7WQ/Yv+eeKmFLOkqjlZjCFocDAf2skEAdeQPCL3q8XwEXnxe1y
kpXzBBcQkkWdwKYdsX7qvxjxXvvB19BfEfRmVcmtdY0tc6M+UqskFjUfUoAeksUInJknAvth70n3
e3GznrkszxEDvWcTnQIb84/nVN8JosDP2fCnpuWswlw5GXqwTcm5uUIGnmVi1s/u9laNmFzM68Bo
rvhD4t35NO8sMyZPu616GGqnayIt/bB81kQJRhd8WPSmvNB0Iy+KtMCRhSQHn/BAYP+4dQsurH/T
EBbKURQZhg894P5BoX3jqZn7iSVv8yT7sfZhyZVSXZxwN68zCYuAklQQM3P9gHY3c4SsvmWG2PsR
XkAR6kRNP00r6DJ8ZHm5cO1vV0tHiniArhXn+PZVtByGd2KDNKCmdQYMj3zoi8L7XUjN/bBbfuPB
SBSKLwvsmwhQbI0HUhqEGOcY5y/VqAIrVnrMi2hlv5tgKMh0fuqB0mZk19yM2f96c3NQfcs16s6r
rQPRc6sdkU8BYUHnWQ+FTOMuxCb8s4NLb46X5M0+Mxk9fzRoC02B2BcUaJwW6gOOyqNjxUCVSr5N
vMjr6+LuMgb6DI4ge131f9BBTvMxoTa9y1p7gD5fBCjYLYoX2OywnMs85y+SqzrpIPg+CkI8x0xd
/Nyme9MXZZ/eba8cclcMF36vNg1C3AkpZNTmfaM2fiFjlwl8QVioc9a7nN2/WwUx1x2yBsYO/ucg
0SfUWecZMs7MXBQN7K2DAtWQIjxZky4DfFLTTB0+DQSHvPloPDyz6env+p4y+gJvXCZJeUmhua6S
Ue56Gut2pdbQWWYh78beHpIUVow9IPLLLpKgAV4solr9GgFWQqGusx5SkkbmU82KOUWKDfZqoekr
M0K+l41rYF1WoetuO02p3Fj81YRNtE2S2d7hto8mCn9ymzsRpBUcoEG32ZFR0d59+pA4XnLrQqYm
ltTduAibeOpPip+tk5A44W+olGsEhuUYhS/fxD6eE1R1pGfSqaVefVUjxr6adgalTNXRmcU+v70Q
WKWNF+aWQjz7BRIs52XkUjLlMucJgKV9GXcsqCX25QMa4CnCKrqGIfiwX/MpFjZaAU2qrxDO95Dl
0zNCDKINTSepUtNqQUB3u9+buLR7V+fjBJPBeHOhI//pBO7JTIcGpZ2hBRuIi02qoIv+vtsb+VcX
zH/Jg54KUC1a1fj6ChSa4owEFMD72koTCRzSr8ba26qGnOIJ1YPpQz404EbtMBsfbzx8UcJ7mfsL
oei+xu26mCCXEIx2UEwzlQvdStrCcWBcnkkf1l3u1FeKCk14lvhRjTK4aHORJOg5Phgrxxm4ump8
Hsfm7/qtqRY/IrSeFh0wCpQj3+MvMvdB2R+FBC+i+rCjtNsdg79tQCQzetxP1OpG8ok8hmLlepM4
QBzYXULVmcoI1ae8D0KhjcG3n4TFkfTGGD3NOMtOFRUsKpQRw/8xi1n/W3Q4YSJ5UPQdz3PgPyNy
4rteDbCAJ4GyCj1bPJ4DkJc7mdS0aU+4/hQ5yv3/CebiBOFBWkXzfdaunhpretCoYItvHjSjXwLb
AMEmdLyv7zIS1dUvdnT/pMsJW75nxPxDo385Sl6WpmCeG2YgeoKx57Zr8i76NrmmO4gRWdAYXSw6
OzrVvkvOdc/ijPU8miaftAv+SFyyHsW91De6h9f0tAvvi6JoDHtk2fQt2e5syCQR0oMuNoD8OHUu
cFO/Rt1e1SpYJvMW0T9ZBuRvnFQujaXmh1m+bzQ3F8dmGFk875UsGe7DKNbBdrfNLN+51AyNihU/
cFsRVtv/aqwgtnnmp2olYLX4fr97qYJTpDGEI5BB0OgKVUn8fuH6ChFh+7Z4HtwvvjyViN1Fs010
9q0fpb0D8EtzttOYmV46K7Bxm7nW2R8Z+9uw5ERPxzaIEjheYwBT7RXEe+wniRw7Ftp1Kl7f7kwL
cYDTzUYCxb/Zt3xQ3IbycDBk8niFSB9PlwefqX54Vp8c5UH54ehWsJ4gYsYQ+z5El7doUY8WI0Zu
xFR2yQr+sW1rKpcla1MyHi7hXpGwzjlVDOZxb/pjKyfSy85GT6uXgUnz7iRon8mR/rOI+9tgHJfs
WO82ixVUzGxw7oXXPh1NtXHu1R7mVBvR8rZLc9LXR8RSnXAxB+UnbUz9hhl5+dRlHfKfjYvvVIQ+
OwfFilBMi3690xEoPEYt1NW5hasWLzu1UIQR2rfmok+ck1L2XsNtp6kMgwQEfSuHn+Z5Mx55lmU9
8CULr79YYJ4B4yh9HdHbzBy0qw/QHs3WGJbSMCBHKy50CkgN4lZEZ9BpgpVsLED2gcSM4H3oB2gA
5riEZtJGO2yy1BlfpUjayNM98M39HBdt0+i2U0xgEDR6yrphzx1eJVi8c6KDqs9uGAg6u+K4akfR
SvX9j7yu2F9d9h79W1RTRUr3LkOSc2lYMuJB3B0UlWyqnnk35pwmsACb8r4E0gzU0KjX6f4yLG2z
vjXuOW1gN4G/Cf23UZahgNi3Hxaz4KACKSkWVMjP4bpfeP/oTWxpzkrYWJcgo9H7BA9zFSQjpV6z
IoyBLQ8z8r4yKtTy4QChQ4v1VXFLM7gCxkz5GR9JMF7SDV2f5GWxXAE2Pj33nXR/TPz1smmqFEZf
YpRISWfR4WEtLhBT5/LTZl7dPx2WszcvBpLHCB4ft1ywsuvPB94iBFhwAKRFP5YrBaZRDY8Y1nlD
FcYpjWCjxfnLuuxN4UpkS7EGH/7mBru83HOoWurtBRavqK5CKXxUSOOSrpl4RcMDrPYIjFkAdiIE
8GI53UIAgOKmgSs8U1v126TV4njKbYbQdS/IEm6KSf3YHQ7Jzyd9FCfPlKW2NNXK9RIHG4dWL6iR
Cq0ijKEhHx6JsyDwX/iM+42yp7qLKzZN6btVJYPv3gEofkqVtTY8xwZIZR7YB+AYe4jUddIg989U
5EOIIG0+0J2jw576RwPAmdrVKW0LcGTKwBlnxXYMFIMK6xei+8yUfEzlWbD9BqrxDWXF5wQ0S9+D
AZ+QB5ZAL9KubllQ/AMmALAD3oVjCxMiUIuybmhPqECQdiWS5Nn4Wg1qh60PeScRRcC2kvH6AXBk
1kzqtC0yUqJX4Q4lJ1jz649Rab+9izQwFETwKw7+wUJ7aOCqcFgRZ3qT47Eb1cqA2ag/CKRigGR4
cjZqoB5sP7+urY1PhDdqSDv1la0er46aX90Vsh9PpLTYFZMYzzcjC0epAV/ZHHxarOZm7p6pf18k
io8FSeSO8nMU4suVYSTP59FhMElRyF/g7TuO1e+UQ0MKO+PA5TRRTFIRS0BSYtQgk5O6Kunfg9PS
ulxcZfHTRJKQsEMD58kk/EYTB7wepsosV3kaqdmvNsI7TlEeF+fL+6zHkKx4WFML8uOAB1RveI5u
zhmlDtLgiHm5CSbr6b02Plhsb1u3fsyQnHlLxO47ZRnv8qKFUQzhKC8M2XGakbd8XiCVeFpDue90
QJFTNRRlTUPRapRf396MI+9+nAYDcu7BZNUK9zZd/1E22yESGFRXJamay0ckegu9PgdPOdDT/E7M
T9x9IU/OT+cXsYZribLrQbt/olmoyT9raPKEO0xdZJZyzvN3qyIdBzN2/WpuqDZ5Z7tKt7Knz15q
kRMvAMN+4GPHsIRHXwSdBS8XGerlEVTX28V78Au4h2yUVEs0pEl+VRhwMsYVlEGqwJUEIyUDpCXn
2V19yhMfwrbjIXYzwGySJ6JbK3Id9dBcSoFzAJy6OBLe5UNWwNM8jaF+ooTD/sEnf6X9BwXYKXEZ
8J70HJhTewPaAl5PQFypRyJEOIcbYPMOLdjxMhKGVFc7UfgxoUhvFIXv42I8fxTHifJK+vINV3AA
DrqY1QuIO1Gmt92263spIwYu4AVDJX3WXN+4HbiU29RJujUDATHvnsTNlMfVbxh2UUsOHTKf9ocD
t+vtNn7nlKdaAzc2vhgChHs6iNpmtj+UaGRmw2lLtDJI892MBnJkV/6ZacQNsc3lMUcevGU6CeuX
BnX2kbRTS5KqrlK6KYraKfCjm2cZBZtGyCJoIWGS4RRlI2AWyMZp77qR4jKuF1HSkAbFrs5w7mFp
AAMI8roly/x9q7h54ZNP42MeQblF1goMk4WVFvprkI1S/fnHiEyqAREPYDJq7gKKoV8Bc9OUimDm
GkRrF7XV0+ydN+Xu24i+DG+dB5Bqc1eHKYm62PVciFHVolKTYpa8NQZ7rXjRrM/J+XJESsFRFafA
/oi/k9aB1ucjn/oYKzgvGv0ct1w5LjCajFFh6oeAVmGdrzgC5S52VWYo8Iqvm/OFWXfOpun3XFvj
QvpZkZDKE7+/GhmiWbjhmC06sci8tvPNYJR7tLC8O37YQhi/KkyNHkgplniskYT0XRaz0vaXB9+s
0JINW31SKWvVzwnZEQJ0SdECuDZEG6/FEY5mXJU5WdhtueFBy5myPkrZNSCyAL7Cois3QbmrYwtN
WXRXw/euHkccELMdYuwN8dfFZLE4JBrqtlGLrBXcp5ngF8ud7MKSGDljG1rgkTCWss+Ak6PyySAQ
sJPPi1mNazktbcdIqf5xnEyjuPZ+ftke6GJX5eyaxOj7vKqhwxrlxKU4AWw5dbwAcJWi0X0BU/Bv
MiUgy0IH5GGrWQwX18be+KdBvcgTJEtKYbcL2mXer4fidqjVTheFuk2LM4p3yey3U28LwEol4EbA
KifsssICHOkuzqmGpP69kwv7bI2YWxMS89gn1hPip5tfsDjcweeOAnt7jG2/d6CsV3TXYfvyddA2
3ZNRkfXQ4xe6w0IWPx1T6cGO0mJu/PSqoDAKAmy7pQF8OBgQFfmuyjC7PjkEjMRs7LlU6kYPwncR
yVaww7JgrwsbjmeQ1aATV3Y9S1fSJQUe1HMzhgP69xLchfq8ijGcOwSZPvQAHGUAa7cK1h2siUkG
L4Dp0lb3ksCjIFO3+h4mS/6D1VQCiySFE8bTbRG8YVPHT1TFJGjZv/jh+TOmnCOGEU3CSx+QqFnY
iUsBuUdZTtkLCG1eZkm0KZEILdWjiKX8LubECuV52KdWOTBP5IkHVrqLOVJONKWT6sTfPseaaJ7b
0WPDRktx13eIbiRjBQSmt83qALfBos85ix7qsi9LYSB24XcnYyObWRxXP6IvlUfk3p/5B+ASEKjM
7kdNMi07rYo2s05p1ApKt2fFLWDUgDF8rbCnrGJYKyty4tHqnwZaHeG54D2J2pD0aAVLdeomGUT5
ZVkFIhrmD9umVdfBei66Vkkai/46nD9/nvl+3kBHxWw2t1QXJjlm3xUI++1R9BTT3YoihM5JwLOa
i4I0kO6pGcg4br12Nze8IDAtHmOCbaf9ot39W7QCGsOTaODxJBGtAqlWxho7Hp6NzKf0xQ35bCMK
THZOBxUpMJhhSlfv+pzzLoxC/QQYtZFUX5qybuQ11y7UIZAaWCGHF7fhktikbOenkeguvkW1KE6U
m4/BP7/xqyNsQFsJ+6ddH8vNNM8pl9Mv3GoUFzXRp5b5Zo2Ytr7FNkoBljxkqKRG4QI3MJX32RSk
YH1laslqOu4T4fAzYtmU9h4ZtmBuJz/AZEcT2nmMoSHZ69PC4Li5kivtMV1+s+HhUDR5tzQnip1o
YzIfpN5pr1mw7eFsxT1H22gr6LPGmXUxhrISUShnDUZFdpLNII72xWKhmD7lFC36GyblKh3nF+0A
Y82fYToOizljWuqAmIKPgZdKZjdSf96pDhwdet386NbZydX5gRskLuos/ofm4GCNMw7cZ/5W0wnC
RwO3viNnVDc0h5crCID/v1AcS85RdaoR037ch9KFIoKJ4aSY+TzWqRWIztGaiRA+NaNupcDU+BB7
pwyL4VhDROChZAK1g02ZGGgpBnycLqbSQDnOHDTHKmkcDi0HZ0yaz/GvrmNUg7Bk6qs+4Qze9rbn
1F6NnybjgrP4+scRys0ekxEzmm01n36MG7WtB81YboExi63g6HAe0Nke9Id6V6/B6/S2o3/aC2bd
sKSiwPftPLknNST/4FLsqURDWQ2dczhl6FL0+198Zox6M9jLDvKuL8JLT1GazLKjVp5ypbV5ctHd
klye40AR438Sxca57HrPnlbbaaO00QLFCq8DkYO1jaCPSksCxf1xHDAZiHSL9D3PSWS207Kyn2cF
cNYMSkrvryDvcfNxxipjL2EP/zEB7yNRHgDBZJhMSTj3WMh04QPzhRj7XZ/5heZj/x0zai8iQY6A
HGU+zRoM7yDKa5Q16Qimg3Re1QGHLrxdANc86HIo+4TtxKW6inwl5oC/atpE/t6qTD5Idh+pWaA0
O423wOwp1WA6aqs+pKQ3l8/1rLt5qV6dWmsHntj2fVuKW3G9ELbUQWn8k1RSz0bInmgHrnQmjrnM
m+4DcR14rJtPHR+ydzBItDBjXvE8QMHeGBsRcvqp9YqUq2gQAFymnn02vlQezkhJgwZAMmQDSKkQ
nRlh3uxzOmhoLMgKQk7Iw6E/W2eIn739oNAMWSbQxeDsRJpECN4DtqvT+bnyD03WwQmG0BvSJffa
VmhmFW7lKoQPlLzR7O8W7iAPOxHNMR4CRdgH0H0X5B30+D0qv0qxT5hpHEY4muAsfnsIgBoLUixz
MBXz+AAFqlGspSEaTxwzdADEu9ut1wyGY7zkW2ckj7GrHpCwe+n8RR0iIadXyta9Cw6ddefoK6f6
DAUCoBXPFZf3hCCnD2xkXPgmJRoXOLOV8CqhTzb6naC8slFDRop6znzsjlLnDdxbvRgU573MTDgb
BxBrKjYGJHeb7FtfY+sa4UJa+dtB8mY2DK5bEfrVSxTvgHAvh1VjKzL7Xi5JBx79NZro7X9dL1fP
pVwSQLgk9AzHzd6mE4E2glnulbtd23Oes0wuwxBiu59NvGeMOdOZd9Qa9Wz/LyvKexO+9bhRajQC
uyzPGcNik4pQow7I+tI0vN5YbBUjJV9/dOK0xfCeYGcTqBfkO77Y/Lj6Mnr7oAm/o+fYY0zwAFhh
OQ5oLGfRmcTeynHUuYftfZd6oLT/cD1RbdnAllh6KAIbiMdvIbDLUkZocE8R6t9yKL4hDn4bUZQt
vtiD3KnNGcvhDEz6GOve8PaKFu7RLQ7uPzN/i+Q1Dr7AsjRkjHdrUgcUxfeICdCjouydP0Nro9+S
413zkk/YZJBF2eNSpJ6F4aPRck3M1Rud29KuwF5d2pBXlxPtgGgKkydJcaIIFH0JAT9sYCXx3rFB
8GCvYeB/PFDeBSppHs/tCGJgvg5b8taXT9WHw9kMd7OaUdSPw8yvvyykC8XAvNlozpLWs4bc7P9r
totOoMDG6AvRjJr1/VjbrfwQ70t6Vg7HMaIdQ3+b5VJvS+jb3EEqPT3GI9dIvjq7G+DEyzgVN4ZZ
oYuhyOTuTvMvhtP/zoIMhvL7RTB/e7GjUtQVZxnFFRMsMiogd1WV85nqOaygtYMcNCL+FGXo/OEd
EmkZrGIeVLdGnHGLJi3YS0dsmF+vC3K+quwJRcwn9BEkQLuFXkDkXuirG2hlTX0G6E2/Kbiy95YH
4+yzqbjrjKvusWHOfTx980nnRjTAp+/wDV2840YzoDLTI2DPFIuoAdq3Evjn6BLkTP3mNXJw2/q8
lxU4/h2LNHyMPqNOZYoHGZ0rNhjBMSHB0po/L5X8Ilpyi7WPmtZwzbmK6s6V5X2cLEPX5QRrztaf
YYNNtSrPccCJKHdGRp/eYq9dc/Qn5UoUyGSpBXe/u2JLPrkjBv8X8f9JCb8jVyeJPGW07X3GBKJu
bOkYaY6TxqgcGyewZLcyJbuOVRl6wsdEpbw/KUIs8nF9xRaSR9EUqwAC1dV9SaRbbyaRSiGpGXZH
S5m8uBpfiqdAzNVq8TD1Ddk1JBLRXn/SwdaB36+c6vp3ICTRtF2JVlerPdbWrauVwvZwUeiw//jF
tihkoJ0Ph66kHdatpRZvb/jrOu4IKTwCeClmgcEC7ufrIIaJB0v0ekmpwrHF0InC6vKlnelrxIGl
rMx6rO7Lc7mH7GjnXF3ywhNVKUJoirFApcwneI/3wIJvB0b5uqGzOcAvG1XKcoWkVQ9UHqQfqxXK
HGj2grcLSIIZRMrE7bH8yjmwYoKJnL2XLQBklQyxB1/VRoMg1MTkyCVohcv1Ut7xmWtZk0NlfZ7f
pzvRZj+3OcpX0+kJOzQKoi08IP6ufzKHjjJKmfI1mlzGEN5bj3wsAdueFJj8nBVKd8hxUtHfklGr
Z4Sl6vxZmuRmxqTVucVhf7DE8sHiq5EEA4rYGXE5Dx8nHxrut7jERW0r3equVvxgaC//JJO8mj00
aESBEhL/OZS+bx9Bg+3ww3zGcmX8NnFitob2LJYv4YVhWSZxRufnE2ucko4MpgRGqPeKe8CQiI4L
z2//XcpapO7DLU3N/td9zeMkN84l6ybV6S8KDTfSYDSO9VqI7ZiLZMYbjLe5LY8tQ0VC3k4QMHp2
NBEN61Ifpm1sHjQlk6RUhR8f3uIbVwDbjPqPFGyfvoYmhO5SxFIzBboQSSAUnRUV/+YgAa+Q696N
DDCJJnOhX0InXZRVL4G9D9If2vUMbpHVGj+ofyW1/QznI+C6/aRdkqLJxMl4zZa6FaMaE2lkFaFS
wuY0VpWYeh50xg8QZ407qVonPCUy/guQiGGVif/Ac2s+nMYn8vOE2jUk7HL1zRzgFq4emsvhkaPm
vmpYO81noTew6FQEZrpfUv8EGA4G2iWA575FCWeOdqer8G1rWa/iFY3JmMDwhSs7zJL0Z6bZamDz
xCCiStcGBpGy6tCT+EKfst5zpkbCFcASySGPASrkfsTX7N+OaYdPnJp+l8PZHzlA5xyMLG29OSkW
An/fRFBerkfRsmxXeKlZXXByvOjVXeHZRpnlBu/weeZ71G3q8nVI+2eBPbtRymrMg81xTSUiiRzg
pV0WlwNBTQpHpEQIRoovJr0DOH1ngwOedKbijH20LreF79owyxJoG/Zha3nOWLEFh5u3BbZuIrT0
m3rdDI0IEz8q2frhCCTV8HTP/AphMsZUBdyCf7IAMlHjn+w2D9Omxe/FHCYtbiAU28aob6RJQqD5
1WnI4OLncGWjt2jhbKViCo9lcO34XW5aZS69smcVfQfT1tgagYhRmif5i4NxcRrvDZBly3qz4Qww
+IYvLkj4tzO0Oqq1XaLgHvSYYcIkHqHbGS72XzxzVx7UQgrhGBQdok9DikX9ViJQ/uCkMgHKnIXj
7ymUcvqDgREr6yWZa5+O9N2kULzgFRe77WXEigpoyJnvniXDhpXtGwpK3OwaX+gSy6cO+PQWag3w
97mF9f4U12ZVLaf+Yifb/GJuCduFfZ5wJdf0dQy/bqazt+ecdkdkAN1hU906Dyk4RY1Sl6MydPIr
lA/lGVM5J1vGDmZnvjGr/NoBg/DpNU2ofrQCxFNmUmTmcH82CaTMA7TFiNz9GKrWgG5I3co4d99S
XJcXD86fvaCAL1deGhMQKVou/KaJiFQi8am/abEYt0rOFMxr6cDE/7qWjBcbvDUtwC6y1J3jP/bM
2Jcn2QcDJV8oFZN1ox4o/PHlfozWLgHE9Lfm20lYwyK8KN0lzO2b9l+R5igT3CcXrVwbrj60haRP
tRryCWvQpfVs4o1ZI+W8CbT0nMEi09Ffh+a35c3UiX/HyEsk8wALDS72TNwM7kLbDy4cuoshMVk7
TL0yUfdTDU2OwnulxUuB79/4GjvVPsgDrFllyDNTu/G3QLO7wYtei379dlamVJPNh/ZhOgGeX6v5
xu9vLho9cNfACR+pDPwFO5q1dJHJ4f2Ba5b0nvvmGA5B6zN03tgulgdzcnt9IZi4DuYwS3VCnBYa
YX7fG49oOpOx8fYdxn4f71lBIaxgiOVp7GOGDlrkZqxNeBXDg5oALbfT4ZfPmsDkkCG1h1ywuBjy
o+TnSsyYSSnEZjWkRhwiTc/kUvuhMeGBi1BMs2RneTa61KX9tIUSUXy030A2vxSz/sRx5PcHA8Lv
4G/H1sgadsjnYyLeT697ZvLpLLvGoe6Tc342B4W7cbx9yOqhzAKXLLuT6lOUCfSr99IB4nZ9pXPd
FoY6cuhnEtCgh962GwtQ1a7/ecLycME+EPANV6Zj+qdXHt5iFzgxHI5WpodCrRbIhSGsJiLR6vSJ
EDSYDQjbVq3d7TKQUV45vKe3DZYcs8db0aXTM1DwS43zDnuseJJTS1wjoKh62WCSLwDpUcQD7gxe
N3jH1Xn4gomRVzhmXsWf6OCs26WcKJzx2DTyySwjIBXKUyY5G018zbm5DfE6DHUt55nf5kS8D1AP
XpHmusRlmAHWXqjQOBQMGg3w+1Ea3kIZR9n8zIToxC3LTIUyFk/E1bYbefR8iKnxadakUMloNCO2
9/MOujfu30G6kLfbKe/5AIeEb9pfHc6KjEIvdgutcMb6y5sK+j4z1elY3z3nxBRSz2lTMvle/awC
PcR9yJihKZVUmwCP0DtQwLVsUzj+bGqGpnaNHiJLZYjKoB1oqr0H0Me4eIUxZ9boME/RkRO3ZuQ1
faoLZKH9/3hJlGZgWutDQHxWo/D+7KUzepwWG7R8mjFGIUhOZWl4PbGLTZERXTzSkoOC5qzPuUwk
pv3ACqRPWrqRj/eHJwh/NIX7ro4UW4Cf/NcTMbOpbshJZTSpt8s77oFLBsfwcKt7zwmCLL3UbRSU
MZSAUrGSGkLnOxYbyjDfiCCqdESZN7gnhNSndVJNVYLGbwMolaBcZr6/7HQ6zoRJxJz8cUmEpjP5
ex+Tv+q4tF3FGWy8XP1B+bmhcAYkbz+Z4eV4Bj5ZfLr0+sKzIrxMJ/KhS/WzvM5aTWwt/rNfr7AV
MC8tQnf8WFYer1B5DyybMsujGjoZWi62zlrTVmLQdix0kwt5zuJdCWn2dmoXjei/W11zLQTwMFpt
asxlbISSl2kYwfy3yFtT+jznTajrLaOsUGIPDncYzBeNDnCoHHkIsFm4+IDzgGvAWVyWzSUyjlNC
Aq9gkKGQxsomAtWuIEOoIZ5Kookpnz9mA+BDRRvZOiEeqIbZnxkFfP6vfTRYCd2XyNW5FHkFxirL
An7QWPJoRcMP7fSk5R2T+yyVS3W3dB78IVczxlUV49OTAbFMRJrwQvToCPnC6/O/1vVUFtmmwlsl
zBYKRp/VDGdtYDXEsfjn++pwSfi+hgDJAIIphpPyUkD0vZpb+VoOG2rZB24bYUeAD1OlxuDMVjCk
JHWTzxHMnyzdT1j5oJLoe1u3MOQjhoSQcokXFGPPzFX583e9M0rsAKhi2EJau1rVmFLL6XUGbBld
pXwNQ1iwKP89BtNV5s6C7zYQ444IN++03t8HxpbOOL6ZfxR9oaFNNTCM7lMH3Cs+JVHkubERVI7n
hkG/Ps+R8q6yrvlAYODA2zJXOBbtSyyWEaIr2PnzOqpuFKR2+ZIWdfwk7VJGnfYmRitWaxETX0hd
Kvt8+xmAYfgdp1Et7VjLDM34CsGK9tt7NEHue7iWJpCVdvx7IuFrjYS8eY2spojjaEWHuG7lSm5l
iBmUsD8YH/Z2UwRzduBgrDB9DqxQyxEyPE2IQ1+CkqNd/L46VTA/CCD4Z6e8p19Kat6xjUJGyHoC
ePPnILEmuy7BehdyITG8bBYvskUigNbbjDYk3B5FmVDi0KmVMZ7m7QIy/LUWxH+bHfhFm3HflL12
ZVSCAXJeOpg8JXVKG3+5xQx3Uggmz4sQ0vzdeOP+Zrs8aDRTVkZZ69kkP6HpsaZBLs1T67j+Iq/9
VEA0XqL10lSJAXka/55q8Vmn4TMAlAFTJfvP6mxo9VTSwBaVfhKsWperGX9Q01qH+oMbcmao4FN4
3qu9yebXErbh9xb/qhe2u9DBx3XCRZhYyOrtDI24Q04xmk91a7jdbntKXC8n30AWakKHC6O9XYkp
t29tXuzFHmfgxtihNNrlidAZAoP/4nzCSUMjQM3u1VWACD5/HlV2Wrux0Q8uibGXkIhNShGC6XRe
HIHEzi08vgB9CBGuhBDjzes4cfi0eOpEseRuRVJ9csDdDUF7+p111V/j5jAsyOyqiNlFZeez9JRn
8uI/0ga0rsmwLyYqSyRTDUsEDuGtXZO6KBhmto4sXF+sJE/e3FmpShvNgCGFc8pCDa1PjfLdiDk4
anv8eUSsb1eOgQXSGeXv/aXfbZpnfw2dPccK4NvEoKjQT7ZWQlI5gutDKZ+AT4WPVr43KwaYqgsa
kGAb2px5P8cG9ty+9MHd1QsH2TLj5txUKtENk4ffwpar2DTHsQVJ3K6ovcrvac0fu94ALQ1Clw4l
lJ1mWs9CT+rXuU9dPCCKug+D0uILUhnL7XDybNZ/uYSFLy/DEg9yeUGpsZGOcAeyhuHaJAML0mSh
W9dBragAhMsmm26ZWzjXmYNaJmf9H0/SSJ7Sqdpwia9xBgybuIyqIjrI3A3A9RjH1/2qXKEZ8B7h
qBrfFer1t1sa2lxm8f4SxeQpaHEs7+i2XLJ9UAwpywzol2dnIqTKSy23RA4T3SyQYJ6MHhuUHiOh
8h0tz+E2OnykmTkb7CjMt3GPexZVENLowPMrDV3sYZ4GNDuOXsJToTjp0Z+5Z9RhibQThAURTFy5
bwa+nKjRTqDpIqylO6l88AHNkdPYu1q4hSr/b3M2kT5OJkb25SKbm8C45NUej2GE4+Btc6d0rCfW
DabCUyDUkoIgfA9Puh4yTQAe/qfIE+VuXQYa1MK+JH1w0JdcV7eFTQlbLVL2VO9aO4fKQR8b8S/Y
ET7rNc3z8E6Ky70D0/Ul1JlTl5s8f3zOxeA6m3ZwAw7GydwnlBmNWl4hVUYFFd68RndJ0oQYDeXU
sRAVhVFjRNnnnBP/BqdHzuqbpRXVQD5B+DU7O6RbXbVxmFJWRvTGzhbYjERssAyqvBgRi4pEU8GH
ML4zxhspxzMOBfhD640xdvcuVHroDLQW+lRYlp37X9EMJdcsPdjZ2zHFU1KPYcreDKqgdx3k4rvG
LZz24JSTY+yMexyYlB2r08ywbUUDAiEMDoi5fr+0qEt3BE8g2Cql4h7GiFHmvfb0ZMStPjAsVvtU
3yJhu+j6R2mKpNNaNXQJHKXK/tuLZHB5xCJme8EaejcvaVXslnRZnMMv5AfR9rmBO060PmChDLVR
dViOHIA/A82uufTIJdA/5EVYNHjCFcYFH8PxePPGsE3LVHsAtcEuYmmCFXW+A7LIV1iPid4PUA9w
W11Gr1dXaDxdoHW4ECX+5IZeGkhRkk68E00p5oOqUaaHJc/OZa1smGQQZTg2J8V4i2H5zDxq222J
NdcBRydQml0aJIj0DdutvKnzejXUL5uf44gK/+rBrO8weeAQ+obp0et0UmZBaso4Zn636dVv1Txu
brXUAx+cyovjpR1QHh06ZkeL2Sy6byFX+vW+DvXX/CFTArLPw7ebhAqn8ppPGaBbI4morkeqiVMX
vI2ic7aelAjLeDrH+FUzKsEFL5wAVKajxkkg9ALdvWM2C2+8rxYw9JjCuHi72bEdAmbOyX/OWfaR
83nGemJAgQMs9wK4+0b4dlaZ/DToFnGYUQnEfhVxAWktq4ibwAsF2qkYj/+oL0XRZcb7UbJUYfxL
WdTQ6MIcpbzfO+R7yAhmpe/z8CM41H0dGA4GVCB69wPH9/3fp/R9N/CXCScGdp/0yclfOhoYr6Bj
q4OI9nP9RQx2vQN1KRhf03yot+mzwMZGZ4iRLurP0A7ZsyuVaIWiQFUXBKXeuyk5WxWyUSjGv98T
HhyMDna1vSDAoyoe4k/EW/0wt6ttb9wY4iNUJGXmkeyEEG6ZSIIhJO7klXPMdYqCxEWhBe+EcWlH
PAH6wF8WkY1saBPYWUz0u/+D/xmay0CvCP3xHYgyYRv5mQXDYN3pShTx9ydhU08ugrWWV+9OckRa
QGNNw11EBE0jbn6f3HqEN0TKgjMxkaz7qG33MfBLgP37DeIhaJm8ESyEbtWBzIlclG7APIGs0iqv
TupccK99FLmE5ukd2z1bnY13C+cGrgYYw06TXzmQWq4tLQ0qEGEJxRbx0gplEeFV0zY6AKjRN4Ye
EcJ1DhEYzgg94MdQAVrO/HGOZoxML6KSwo4f48eCGcxUrspqcElO3oqUS9T79ypT4y/Najw/hKaW
wFTtbaovpwyMZ0Es3TIHScNZh3OAoHMm4CfPmSu8egZZay1DUeIsawZhGxRENPtxm/PRtwVTimew
jYxSH5qxN7l8OD9X5rq0UnrDt6O0TStXhYlS1n54osXqS+l+SQ2fYG7syGU4IWdmj6Lm4JgDV0Qt
5z72yAdylykIopA8sc9hrLVUI4L5ZscNGIECenfpJcTTuL+9gd9GaKvbZM1Hv2Dpb3vDeZVtzrer
FliVpKlHi27HLlvPVoSpJsZtr5GtiNwhzGDn7ZwQqBHA4OTDZuaEtmvh9E0JyYzDBUrAZaA4vt/R
BQabMLjkb/EEjPzvzw5G39acdeQoY/ea+YSXM7CkLBemKplzZ5rKXnI+EA61qrlLgfBVdrizHDS3
SmyHk85z3Dz7GoAtUbmW4BLiBWK8zl//LqPF38G3dTm12E+lrFxS+/Hd/WAc9WNigJJuSM4JIO8E
FWTHWOhVEeAivDqiaSoYAAbt5dF8qTePQ3elcd/jCsFHPLdS6/hVGIEsFCsX7mNfZe44m/CgpX4l
SobEeEEiUkUbsBcy2Ee6gUwUaAoRn+0CrBcyOB4+rIzcd/H0zFUAmxKKLR7ZlzEcefLtltv3mXMO
+4EAu60XPmsPc8A6qEgpI9mlWSdSgi7v6elmEEuILOQgEglXGETzygy7XaMUpGEwJYs8QAgzcIKN
4yGaQLcYRiyHDdAbGcRI/kdzeyMPXNznyEkHA8gVWTYDO2CKD5LBzUYw4g+x933ctFYj2prvDWs+
JdBhXlsbjzD3/2P2ocpRblYvh9u+MGyAkNaxJQXjRU6aHiJL+GYDLreYGJ3t9KtfDvtrswiNIymP
+doeJ/GGaQQu6a8jFkxt8wylFnadEuCwimHP3tntzxhEwfYQj76y/13cAvB7q6Esv+jdM8fiQL8H
738J60vPkzZS01lysEnsJ0chYrfAg679kp1UcjJLa11pPITda6OP8tGEZ22up2mMYTfJkYCC/glS
MuqSMentVufuZyBq+HYC6hNsV7NZysDEm1E0UjrtO84ms4GpkNPw2BZESt5Rvv/A80pJs6r6EKJY
UtI7jwrwsZLBXWfC8prRe1Ixabz6zPPSVZ6qtrwfp3Gg/rt2qMYl6oJeG+GfM4Wf0whia3laXZHv
3zBgs7tKh8oKCYLWmMY3jSG5zano0m+0MlKFpOceqXnd2nzZuPO8e5Mm4t8Akm7esn5U6atCy7C3
Z+x93NThjT9jn3FXoR/pQOLwUsptaY5/7BAvDASvGCupeW0mIXcsjKQL6FWbyA1KHoToH65hJvzA
kQZ7x0Oce9k4sYIm7RG8V7v3SkYTNYaMlkIIpTLfFkNPC56pqewiiONcwOSP8LufD1MUWrrH9Yc7
zVgP2+JraulP80XUMQv8QZry26IJePtvWvweJXbcEplNo8lTJ9MipTut0nfds3H+0Zz8D8t5Ob54
1HUx1MNoFEX3rjk8H7dzaowCjK831vL5QlK0GKgQMbWEuPV7irnJCOnaGo/2MaQ+R2DLnLcmYB5B
48IAlec8dZoMBrvr0NBvchchokq4YdasyBFVuvyZ6blq6T+IISPwfqI+QVkVq4MVzYAgzF3+F3N0
e8g/spGZNGZpRN3qRInCxl83efLXivSizjY/XDDltnt92uyrzjR9pKrUXupwuyZ7qhefR/orgdQo
AHZL8/CJM2oyt1zW7WMqH4BoAsp02a3XPUdNRbur0Eg/Xogn7GLjdE5RwAirRWjMCkzPeprSanfb
V4zHv05j/6C+Sx6hoHtQEUp6eGOFK6c0NXYH8s1RxJ2VmCUlEq83g65v1yzSg//Q/LiKv1I4EzWo
hEZyV1iomzdSr7u8H/Fg2vQ8ggpDiVS/qHxjZmI/MqV58fWT0O14aOK2+gdPRUxGqtSasJ9ug4BW
mUpayVU/CvKJugBrQDYDrdkb/TPTDSzh7ExhMXf6ITSpBDKxhKp2Cqyx9cKcKta8K36T1KrmVBE2
s6JN0D/aF9JCob7k926hC+lt9icX1jxLXQr2Vd3UldxaQf6lzZf3mr+MJJoWL2PjyBN5SjpZAF50
7oi/jVE3vvETKnzLNOBsp/OdnHEqRr8X0aOSaeRELXpNgHPZqrcdBmOATq3HzmEmAgOZQdJcrTO7
L+bws6AGdYR2jfbJ3qZzBrUpUl0G4B5TCYzSkqhfvQzHBKeyz7/peMTcGtdyFSjqzuCX5Iv7ZUhI
hw01lWSrxZSVDmuIPsFqp2IHFKRfHcNJK1UJIFFz3byoFn4EXn6OY7e5OLcQNmGnaXcBhKlMdZ7A
JYvHbCjCLupuRhA67O+mfFrYWiscrXGHC7aO3jYJF689wFZD+j/yiAwJMfFu07jTxFdedxwf1b2B
tOr2IwikbRWUg1eF3AmOVEVAQ6i7hlSUBzU8WIVcvxaZ92gWQ8YEhh7vrOnJ8bWX+1JAGm3G2X6b
/uQhvMGGt12fCZARK2thnBYoIIa43vNuHr1nszp1qt+kUJMHGD8WzYcYB3z1MCNjnwI0COljBswF
OWa0T6vy1Llt7RTr/sEvK2diqsCPJD83KgMG+bfiQtc5YBaDtIOTLYSSuSZpzfQ02P9mtwcQVKeD
JtkOvNt7qIlztc2p1fY5gkwFOQDlieOCrmBravhoZvebnPxM4jMSdTe/+bjAdKI7VOM/7r707xNB
CFNuuW5u7OD2mB2ZmYwg0s3mqeUw62dRkQ4g/RsV2g4m7t37WDF4afmiBg9DtOPofYYKKqbFsDQE
ToEu2FMgAnCSgbnQMyKNbKggVhhb/I/JgD3qd+vBvsgQcIjtX1RlExiOLunUrR6kJ5Wkdb8TH6/b
BKiXOd7bAW9ebdNwkSF1bHfJtKK0QaMYeY8mP4BTnNiRcab/LiTu4pgcmB26Y9wR9UeAyJad//o8
QRuFM+RyDj2ng+6UsLS6LAb7bIDqTC2+hIFiiW+qWl0rBZlKUnwcFm19ZiGF7bLABynQuLwrj/0d
PXLw5sFSH9IIjm3c70ocum5AaO4HWeIaGFO4tl9dKSzfkmvIXlLrqnKPTt5qauNtr+UvS56mmNt7
fsk0My4Z+ZHlPKElpshftBu40Vvjl+F8OqBA0mAdox2eOdTIXvBLa55PWZXvEww+UA3jsSOqblA8
vFQ/sBcRflGQ1d+uPdS9lvstfS35ENqBQdeKJPaBWoy7qVxef6dXuJ1fyfI4kbxDEwfDi/czxxh8
t2HkM+kj9bm/AVLEMjUPM30BdeMI9qVSKbiagZitmlA0xXQqLYgOSJd0poa8oWTTsjesVQJxRV9U
7zt70+9ZdGx01mjwVefAL0nxTmyK3LRF/Jj1vud2sf2RaaqLXQOhhRxmRrEsqrGM88zG3otPEgj7
R85gL+JLFgot/LTt9pN8J7YncdlNpOLrV23Yo9+dkP7Np6InT83T/rpLaeiZ1mgKpyNOyBUmXVtG
rhph6CDo3yVnSfqd6RkNVvx5j3xdnxL/I35YTwdOCcqHhTgy3cSJXODf0jCCXEBQVKIUbu0oAd6w
xaBc95E0cFb3qHydO4gsYdOpr+qI2HY7ecZhfp38QTZG5VfwiPfbbv6WOZZ8qHW8jtPAeJFKueDS
6FluWkZOG3upYdKTkeQPfPpjM9ShtgKbXdCXpJVCQ5Yn8b+KkvWp5fEqGGzdz/YGktiV30gD0HD0
JdGm5pQ/dYCDMceaB09ut14iPuqzJ2QyorWyzMGAflOCq3CVZnwhitMISOgk1/2bPsw9FpysZTZD
1B2baUSnvdE5drbXXxao2u7JiObEejrxfQSgdosQG/kJSE4zcKLNzOLzpfO1DBg8TKmUG15m3FKM
V7WhItDjoEY3/K6AGRy/+YbrAHudowCXC/Yl5/xY419Ygg9EaKACn4K1gT5/Z39XEJVwvgXzSf6Y
eiY9AVtA/oZmalExcSwPUfETTzbyKvmLU7yFQPL0sUaw9+hbeY1ETOB9pkoeQnawL/ul6dHU4Jo8
Ajx5sPtIpQmdw+H1ffA7P2G1XYsOpG+Oz5HSyaF1B9AMhNN/ykVqwFYJC/derRuefOBXHH2f6PEl
Y8mdjXvM/DTd7I2hG70xWqSSejIkg4b3bVOO87/TfpA+VAiJeLLhOU2zSD2X+/cJ3parWX8GGcNV
hjG4phpQakiU7rgMnxAvb6Z48jELI5eVfPDjs3YtheFnFb4+csiCM7q9OKpFJqX7taNuvpFBSGin
o5kjrQoEEZbjS7jExDv1hvztk/QZpAFNHmP9y4fArEVmnCVHU8qqitg6wHtglYkJFen7V7nARGz8
UXPn8X5t8kO35fe0UaNwRd2R8nGjpyFWMPm83ivet4Yce4/cY28lIdrmvBDKd4AFI2Db0SXBvVEk
KOTyRZuwt22e77HSQsS1xiexfsuNL5BxAbiYiQbgTD/DoY4hlGvFXmVc0t7MxIJ8n0l1mKZV7lRU
qGd3efWRQr/fnNmLBKNgdR2LHEQbyyGvtrbF4oc1N3Fp0rTO6fdFL0XxIy7kzJWSoQkQh/Xa2KWt
gvrU8BH158SahhV05dnan1cP1kcQZieZch1dhvZwarfVn91BHg4UBLucqCwc3AaX93ffy79USYrd
cYBGPUkhfEJouVrWJJcrmmBUUQheYfngXnXo2XFFHSyeFI9xN9fXiPet4rZW4HxoFspK1+0FGHNt
D3dLTyYtcHa+XJmRJjEn/sDKQO67FW1arH1zkxumylEhOPusFkWv17nxQkhnqmEXhOULCXaNhlUE
3G7/i9WkeB/0H9Ue7cmk75JSu6sGCBYUsCEhyIRoq4yPkZwOCAetWtdKZ5w7K85Ah+B9qBnVmpAe
wQ2UpKt6ii4yRM1MO6cWavELGYyzIag1Gub1w6ba6oJn8KwFO8yhCLo+L4tb0OFpVph8bqVZ3iN/
zGFdkREkldpNnCMwNOp7d60ZhwofM4oBCb1QMc093+OWYpaCII6sf9WoKe5E1QhZ3h7t5GDEUEt+
pjEoHej6ivToWtzNs2aHUc57CMnTltMgmgTPvKlkQ1US/v0Q2OuzpJVgV0lMuVtXCDDGe98xVJNe
cBX/4HF1wKC8KjnQw4wQZAxj7nCy8CPQgfloSm6+xKuxvSbtmjf/vKPMdOcpZuIkrXW0lSWPDd7i
eeu5fGCr7jM8r5CXsBBRuK9bM2qTFxhyzaYehFN6tgqXQxOTtTJn4vDyYXoO9tKPTHC6gCAkF3+c
eBO30QsxxRVHnn0h3ngv3wDXBlQP2l9ny3p4gTJ+vekPFoY+3OcH5bbqK2mdIXTl/eTcsxGaQDVQ
wv86rLsr5TtXDpwDKs44IeJXg9VJyuoBS1ECuf9zr21og6xn3kdokCVkCx1pFe6nPX2LMp24Kj/J
E2mX62uosrwgp06wle2BaJT9Vd4RvE/T40Tc4PhggKp53YPrxqTOl/dGoWjh0Lk3c24qCh9Y9d6U
3L24LiEAm8F4tTJITkOAIYbHTd+kqw4meRx7BHaXuPx3A5Yl7hgRNvN17eDFI0d8SYa/qpDsl27l
SGhebbonJ6UMlK9X9YwuTxGlkv931g+3LSrn2wOd3Ky1ZCTjNKHRAZzAL1S8n/iWKHS+kLeJFG7L
jfQ/lBsBgpU8VkCKMl+lVpOC+dK5sr1rzfxjfrrTYOQGDUNRY/wyz1rkPMSm0/N+1RsC7N6rvTrA
464IjMXbCNmIwMKoKdJIKK6sTrokXFv2i/VBskuGv2UewLBB/A+Cnuar8tvatPRqAtu2V2D2h19S
QYo6cPgx/3t9CNMnnWMw6DV3NCM47rbS0YB2UGtFwt9Sun7O3Ow65GrRyyFruGIoLsk6UuGHLCPP
LlmyvOrGB7S9O3a1VedE3dYTs1YnXvd0y1xwHv1+rESaO4jfLTCMZ0pMlQ75m7qUodzLEcCPXUGe
JL6wuQEhtJ+eHIsMPEcXGIe7de5k5SMf8OBUsmpRNZTtcZGs/0e7TcJZGEXycCA5VX2kOzrIB53M
zn5Ym5JH72WGdqcx9QiMiGamhZ0PLDn8XPLaa6iuxAAMFFp3NC4iuf9ObwBVR3uik2dQ2da2PYTx
pSrSBZXZYmhVo/Wpkey/UUHR2zlTFjRPMOHYOe/A9lmYhgEJqbl/fBqG7pXI4IXKsBmHLRy9PLbs
RIrYUB0KLKsBs1tSm/ayaT/RJQvWSeHwrBtk+/sFVlbincdVBNv+9sKSOG42ICB+eWDC3YCR7UWO
wIK8ITv481UHpkTAE7gA/6El9NZ7uLHFFjalb8HVhDmLZ9EStp2/MAs4acuObdmbJX9OJIuNEa67
A1MWCw/HzHbZsxByfXLHFL6q+RZI75PbmuSeqqLchw+PxU0fVKw/H++yaNfsLMmNMTdjoEj3xx7M
jhzVwaVEWSGdWXIgwaqRcOLyoAlUiEA+uJpt4uZnvFbyDA/rTzQjCtuieou3pUT/NTGCC5NZVpfj
oiiabzITmLNFuaWajrkcb/CQWYVU5ep5+7ly1G8cYSTBptrUvwEYGtl9sCc3Rlvno4RRwB+5VMoY
gaqYGiq1030YdvcNfeVS0jAPcX+Y+dvANoL2Ki4NduoZtb/UXjHY9ca1l6lNndoxq6NLpKgELa6e
Xvc5XEXig2o6d9m5x4TOR9F696wEgRBw1wpBtstXs8FPFCJ3yHB8V6rw7UPS2CmVcFMDxdFoZ3Kj
LLnPOcffYVMWW9hHsed/X9LOq8XB9wOJRbA9XxYU4Vv01MyfWOWKcQqnqRH3nKivdlmEasFt18sl
OPtWtM5SuHHHl+2XLXdbuJXPW8TvHa2XHHe5nCq+L4Xu/Y9Tgbq3jNM7RzS+kpcuxejt5+PV4qV4
o4cl/Pab6oG+fgNaCxeTdxqJ5/5xR/zvC/u/TQIJdSgZawpzPb+vQ2Jtsq/Gb8Da7Fm/XB8Z9oBW
4j/3YvMi771YeQaLNvVQdN9+Dxckw8znSxlM92/Ub7MAiN0x9h2/p1lqr/O1wJnoG7Lx31gQod6B
ChEIaRtU6kHXbIuF3H4YXSiEsJAp5ncVBmXu/afH18Vzb1zVP2xT/b3yQ2y59J9z+N7QJ7v1/010
NPFMNb63S5W6Nyqe3gRjMpU6RB5YnZWpamo6jQlrDGzoibTrcm0yOS/xHSJwRLt0dZXFs90iLTdi
keBq4KYjTRS2SfyhoE2nKlpIF5a+vKCEnj2izkkkGabYCp33BkLfwfF1lNAEpee9mB+i1e+fczZ7
frzfJzLCJUcoKYzabwpBEe15L1HyGoBIg0U4rfYdz7vxqFc5u7D5T5oZVBUaHmLJXuzH0k9AYphq
hgS9kQXHw63NImaZlbEgX0g8Jy58W7f6fj0VcL1J42nLbd5hqptzvyAat54hR8TMIFA+N39iATG3
wW7BuNAcEcn4WgJJM5AwS+vhw3Y5wim+YCDxnkh5evAgkPs/qbHOrgA9+X1JtJ1MqHnH7MAbnIde
Dn0xL7no2BEv3wX2Y0AMWEOQhJ4JY3b5MEYZH8+/cCz+zsY4UdbBwKhz0IDPNeKPy9iY2yN3EH6g
0CcYq3n5sYneDUxvPQv+N9CJOMIuN1B1EC9OuLYhQe7Ni0LnAo3rzIb1yn8+aQr9eamAta7/kS5m
FWS9MGr1fxh2ErfkaT9+2Kq5xq+jeWbpF2wI6ZHu7DvtzMNyZ8WpO+7BffMM9uOet8vryIc5PJCp
FPs101+BQicCbCmEmrpOTw3c6DmINvDcOiw6dJX1Lg/NJUrf3dwQCu5X/syHylAXoY5KlTSNiKkX
o6TDBp04yrRsR/Iia5ACmCLR5uMVKaAAB2IRfA7xNr92RI/9QJNd4pumi8HeIiPH2ltmrkrx2iZX
bfnA0XpePDXdkSInit/7FAHbK+f9rCyiuY0/g+pdMPdUSn9aG15zLDpia8IPY7wTc7DN2d6lkqfN
wu+sZTE7bn+boUvxoIlbAsBnZckToxePbQntTHVf1oMuqOhcRupluehUHGymVKK28V6iKWoFdfkq
O+1gMjm0dggcClpxhB/V4YftIUzSpk1gwFNKNHU9FVqRm1C//c1APyYv73SxDFpZkUCxHBFszbis
3DccqQY/M+lOl4019khrhVkpJwMoWsyJOOKCQFZwoE7siz3Z8/TqILT0+8IGVgwskwsaafUcJsL4
0FdCv7YwyqW42gZIRhmaTadL+AaCQ7VJZM0hNORXFk35OJQ9OqmIj/cRzZ1HTpQf4M5+FBVclokM
cFNR8KBqU9hH1WDPSUC/Mr0kY1XKCPsCul3ZmMymfYXOBZE2jUcw54hHaY+cXoQ9BLcykfWjBkTJ
++L9z+xyQ7tj3MPFm9X+aEImfHx7kCyf0aShhXDdqadrwwlrZe+vVLB2IMGgpY9BZ+w3He3xH9St
S6gOkUejW6ZKwOEPufYHbIQqRyIEEzD4HRYhK7YgS2pXg+5ho79xDsxhQplc/9mCI7Tiu+u4cv8n
YeAlcho+JOBagPIg38/K+rhES2PJ63h+QNJQHQCkrtlAhvaRBrSNWU88GPXAaAEVDHkE90D8dvG+
LDi9ujn9xMubGGqfPJ6mmBbUoU3+jiXClKTGUbFIs3i8oiOF+kq05fL7VcKtgqEKMqYSDZcZI8IF
Ti1baH92esbw+44i5IQrpMO6gRiBp+OZO/68loWBrOOg+l4mFf7sS/POUs5G1Ss5NW1e9Bd7tCac
OaNCq3sJt3jUCVTMkQMYMAOokLmibngEOly76IWHEsE/GrbQH3y8zbc+8v6wK8eGy0V+lZlsC5tN
In8q49GDKdKPFBG22nGfYy86Po4/ASGWPsIwQEYS94NIgv5tnuUZyezmR6QuyJQLNOmDxY4N3mju
QCAtu7K8b+L1qZC5eB92MbA1MpSuPMz3G7FGvHeOi61Hj5L93mvSWPoY0dIY5DmpQ+XV4aWsHHQf
/oeS0aB2GKDtzU6XZlWfM0qKdPKbpeI4AfWrqA/2lccFPpDeTrm7vOv1Q8/mFj+DQZx3GwV2mPK5
il8iXkprmyzSe38agmz39SvW7mFKbHoyNcE3RRURHH+nvtIhD+wn9Z+ApPoLVYFtX99KmS/lKC4y
3NdLhWVclVWmtw7XCp+PnIoVp8yjzNUgf5d6RU9hLmWp/0RgI/W9Zow4/T7Qq/Dj7YDjGtQ5k+E9
UPQfxotwzCBxtFxga0YUgw86Cz6QFTVF2XotSbIAhLtGVJM88Lg+HZzVcyxDLK3t6IOOtoQvIHtg
uWjABW4K65SFzkcd4j4LsMPW2sNG5yStxiT0/xSF3xkZtJbPygvkWGVs2P5tTLGmW3ZJiDb0uhGz
cZm8iKqBoP0yq5m9EVTEug+5WpXjRoqD/2/IG34ad3RflW+qfcIJRS82z3ZmsqG8FTef5HHfFwEh
1JtAOSMQ3gfzcVyoG21r5d3BwGLWb0Bgh2Cp+5G6SZDMPysR+c7wXZl7GMsJpkHJMriAWfCLr35N
MXQ0k9C0RsocDKL1G162h8KBWAYYnjWc6Kub23wb8i6JAcfnmxtmsSVsqKqHnMfM0iW5XMJ72f5U
9hGnk8qnWxSTFFXP2d0vtkSbJo5FJl0LIg5FeJA66KJMamyKH0n/QjB8tPXaK87fgDOt/ekdd0HH
DkOstkchEuZi1sRk6r4rSdQu7wINrmjmo/Iok7UpczN//s/BN5S2YjTYnW3hE1nyMy9DxYziQvcR
Yo4XNbQzLz0KZ5+8f0l/HfX1SU9A6fBGT32i+I0CJ52+mRYMTTwGiRm9KEAyYWii5nd56ikQ60l5
/a7hxO62wo2Tl62vK5jzUIzLgAY9Ju7FeFno179YFCYn32illpjck7TNxTBojwa8r6D+afmTs4kW
Alift8QNLhpres67NH5gmRxm6t81K2hNMz8K5kIKkxy1lE2TZ9xS6r44x3WtBTW55N6HNYuXgJsU
huGYfKJvfn9o97LnbC6bqgVI/VsPw5JJO/1kEisqG7d6h4SieELImJVPaFulDDJHmhNfKQ1sqSs6
5u6MVE5+nOgM4FN4HXDz+ADUL6yQg7meeFtt1P0VtDQzPrOvCt0jCZLi8BLZEphAIjBEPNxoyZNn
L2mokko+jAjvg//+6DX91+kRMmX4Z6fGuXMUeZLMJMuh0tiYdaRm/+W3LcQ649+38FcUdmM6XSVl
cN+Ow29/YlvO4MwcqheB1rKC5GspLzlsQJqwu3YARqUuNmKjGQ+dbfBa8Xth5jrAoJVTV9qTDrUn
smTW5lhileVOH19CU0EGRensztHeKemeyBGXhkyYxsr7QKd8G0olUI+NJ+kArfUiEaZ+f0GB3IIe
srAe1Bst0clMXnB1uDaUmj37vz1uGwbBio+bR2ukOY5pbHoRVnUXd5MfEZ4zjlhRBjzwdHZGxdo+
Ky0BwJ5+ymo943gS9oJuNSkmtMaN7y3r/iL6mZ8BC4IbtPUkjBgoxN7uDtWdMcAiWmXwLyXoPGUy
fbSGS3xukn/YHbbagXv/My1jyc3tyIwhZKy80XqPiWoFuzmytlDpadyZgFKI7dJUA1Io/wZzIJfQ
8zi/LXrxJeKzPbZsOX7mDQfvIVZPF8dk5sQapUongq/RrAPbNnYtg8bwN70r/HiUNVCtfIDiCq3V
4DfCwwDrYoZ2yGy/vXPcYlnhc9O6jGz9O76l2P+1k8QJxd4tKmykkYpFcSTU1UJoRHb/Yrc3E5zZ
Gu2Dfn4N14ZWhC6ZsIwh1s/sDAz+Um+zUjTTz5OwSzvetp1qU0J3rgD+B5+JQTfXrcMd3kIQeBMk
kTlGTN/ZKZYmLWPWJh0ch/emjTo5zFMvQR/2DZbAc672QcpCY9TI5whlWgEiq1aJYhEDoaH6NgOW
71cgAq71qJCjllWl24v98S6p0TG2Nnfm39cDofhueoONfEs9m7gTDV/0mrmffwx+xa1k2TLlt4+f
nWtyvhW3Kvru/G+nUhrWpLN8IpWowCZCTmxbQYzqpTyfXHV4aAsgdEw/MNhcLJPmzp/0rU1NtWG4
70XW5u9Uage5Tbtt8WdX7hfoFN50EXqy4zsfyxwwIoepv/mKK5tIWCA8wDXSbO43qklEa5ax+uYV
LolXzSyW51ljPZZlhRmAQ7aYBIBq5RU+CN2SOCmnEhrC27z+UDgT5gT890AElBSOW7HcsnGi7BfG
479aqIBuMaU51hGmByxx3524if+Fj613aAjpXO9KD+g0tllzvolxhugun8j1JMN89nvTzHHHTt5C
1bZDnZkq+Zi2RNDYG1msaMj/ZXLNv0mAsOGJfI31FBwLialQTJCU9tyeVXL6OVrp3YQlx89hG7we
/el0KzcZr+/RMQ66bcVVQGw/KkLHjjeb5QNP9LJuWjNQ+Gp8PivW0y64R3KYqKlWi0Q7ey+UR2RS
TC3N3upXSL5am9neCzOc5wuaGA/S3+2FVGfLJxJCXxzaeN7wnedqDH1ko2WhN8NersZb3qbw5LPA
ufAtcZWP9tj9cBf5H1MaAsO3OqSyyMqEVJl2KLLLis6KpwLwBxB3y7Vls2cEWWSiElFXrmllSqvR
vyn36URYd0SrRBZ/u1FGnA4+6S8D39nwuXRzS11Ta5FKyXTg/hCtAWlnCSRwkcZ3hSsvkZVEAMQo
qFGLFvwSN71iU/asz0hLFEOX8IVVOGLyWgKkIuz+87I+2OrdHeLzwneacF2axQwRdgjbA4kxN9IH
UlabyjRTXp7rWe+gnL+kjJzcjahY2k+V3Lbp5ZXu+vAluFsvPm5CLYgUd9se8y2obpUCy09Bt4aD
p5nd9BS3Qr3ImZw7pl9H7miB9WgcPLSZic6fTn1oSTWGVcI09UurfgOCJnnlrkF6MhBVFs/9RSlp
9r484y00pKlBc2Iwsuz5aInZst0ny61wbLmBcP498YnOkxQ651GnumypBZEpPA4qxJHogDJz73VS
BJUlCNv0FRHVHifRk4CKTk32t6HiUu8iqXu6nd1a8H9XTvIYtiMy9WXcQ/cQ9J3DTyhciPnkDR8y
oOTerTBhhPDyxxkUj5G7H8BBTDYJku3n/HcNWdeToYxkSY7GTBanXBHtcCLTDtMZ6IFXkEm5N/wl
IQNI1XvyjAB/gKJeW/P55iMO9kwk9al0IwxR44bRrteuML/591UYDe0T1bMspyRffRpmeimwSp3o
CwuGFAykqXphQsD23K4xzIb73mzLxwJoJxfhCa0NCxXEX7TfepVRC9QGskJ+WQkSSQmcITlla/xl
L0THTjJTKa6YHV1iZQ25lSWZNhmtY62wpvwAwcnIfIsz53rCBQFdo5zTzPXiez0KmL8qgYuItL8v
WkUF058hfSSSBZH7SxnQ0czoJaUvYUfI5nJERWU+DFsdv74G3cWWDclf9pcGkXawRhuEA6spO9ff
Zf704iNEFSN+jdhFyPJKY0W276b9zmlG3GpuCpkatLDlUBdyDvQcSKzJFlNo4B5CELMLwwhg1ghP
RFB3EV20noDK0Q+kmP0JcHGos2fji1LYuRKkMCJfH26tXOHGO1f1qDiWfoW03dgwgS6uwb30RgFl
fqRx6MmPKN+0zVmSON4oZx2Dutvuodr7a0j23EzhoOUOsiQJYDPknmk/o84D1+oSAcxYWLu1cs0K
6jT4X3vzKIb//dYYzzzibVNYXq1R+ktmKAfWaPNICxRyqF8SeYFneUCThbCLIElKGN7N7dsS0XX6
Q4qgALklt4/bHjhuilGz+YzNum2Y2X/8B0x97xHcBMG1WX6fqGXu8bOixEywwXMr0Knu/xkVXDH6
nQOb7apCSz2HIElzvvjk/mozp/VuhSBagObywcaB6a+nud3ON/Awjhn/J82Ax4yZT5pW65WWbZHg
E8RsbbnWJ+es0kP2nNZhrbbhS8COM/X3wnerPaRk/ARnXXYzXMOc6gaIDqOA9MINxaSJysUEwXMO
GI9gvOdrZiJgU1Gc3Vg5ofL3ccvXBJ7JjNtrXtOu2rL7jiiUQFXoNLNr3CTOr76bAJsaSn/gk16l
I+051gBWqPvUudlAE8y2EHv+r6+81D1IghkTsYi+RZRf1NkpDzQY2VC39vosWhtQU+A9LKhq4aC2
rT/+gj3xc8G2lb7vTpiXr8pM5DzlxbRkatV2kxJXfW/cVMgR9/Ce8GRfK6aGHBlwm04TpxQxxNIF
QuP88wQKQeP31q6FxF4Jf/ReaVdhAHbUseIRyn4nMrvj+PFCNSOj02J2u9FOlcb4/7fG78pWsT5u
zLWSH4lExwboLt/0soXkzJkqicw+P3yL4HAq3AT8BU59FN+xsteyJ7Kb9WLgKLx0RanNoeEiMxw4
hqdaPG0RkurZe7lh0kXIYwc4YP4HJbMvnLSee+L3zaB03wbfleIP50QC5zgo3JKpuai3at6Jp/MX
y2DDxJPP4/UtzDefiFsldzhxucdb1brxjdGpABPphYPRSp5IDRJsTjcB6EsBSvdKYX9t064MEVHK
SF5Co0gTkStLSWnggP/Qm3mP72zI+2SzhB+Br7m73UCMfeZcMjgJ/EPqkO/s9dYpBJSD2CGZHNGb
sBdee2psTi62eNwD9ULpYsnAEZz92Em6u1rWmoSL+75nXqMTzxnbZ+376aOsbGNjVBzNpW0yxECO
frSJhWbf6vR3l1l+MgoVpobOjX3CzT17J+Q6e0NNc0cfyIP+TxoieiX5BvJnY9925Jk8QU3XehbC
1HqflGh0o7UkKUFayY0dJ+FLTHiMfrN57h85Qx6K/+MT2f766VTLYZHWh3KGE+iHzlhNdArgNHHc
qIWVKiteLS+et7zm6U87SZI8T6VhLHJ24UsB/TaZAhOs3BGb6CIOchyhSz9EHFw9VMXB8pTXoUJq
YbUltpLEydy/A3uBog54MUS9mMxN95RtnHVnX4tJdvPFLUEDizwhi5bhhvDP6Dnihsvwa0LO23o/
74X0L+lt4Rk63uRXq2UpLReXEVkOzl6xXUsgsO8xgsoY25Jh8xCj8a6hBjw35rMaSKYyqZXyy93S
wbOXPLreP+ZZvPOqcgKJCVJIbVr5YnjuX2eFJLxKKujqXToP4Sp35f3VS82dchG4tviOhd7H0cKV
RjQobP2zv7Y+J7i93p/FJxYbrJ4DDtStL7i5VZ2y1TFAuEz25T6JnXhmxAwBxNEU861UVjV14hDw
JbP1X5seavHoG+J+/m95L0j3kSxHt0Ba8hKZ7dztiJ0N2r/OBuPrSoNiEmHl1f/DgLgF3PMz+IVP
MVTD39OU8wyhlkClNAEdGaVoYBIBO81AsjXR4QtwMg991gy3LNJVzro0+hUR0pgl2qj2LLTqNSNX
A8vg8IqpMPj5fa4qCGS97DAm5EN38F1IZd/R5YiGIFj/tB8o1xP00AIY+m+vRGeVqNUj3kARAL/d
sItIZeWCLRfqpwlsflez9VSrEyGqHg2oCrrLm+AwQPVe1Xrqf0nE9v5553ccODvk+//mmwXHAGUn
D9OglR4igbsSeDZbNqDuMjlrJb8ZMtGFnS+K5DmHmEnsaKlCK+c8HIuNTs64cuRn/nl9ev1fBfmc
I4gH7POsEN92Y+fdVoyBHNxW++Pk42C3REo3DnYoimFO1BTZVA5YlZ0yR2jCEhrBeJEb218FruIS
QuG3wDlW6xvfm7GPrnwV8nGHuQgy9cZbVo7vzacX9djTkyhNTqJqvN+3kgsLE2d86Da03BTXewds
2Lp6+mb40TsEH6sYOv6m1r+r+YnU3Jdsi3UPokdtKmKl1ueyKPjMEfL35INPPvf6Sa0bu5w+ivEi
cwwODVhlYtxaSOVHNLMF6YzcsCwvgZayFUJUfvLw9mOevDNcvR4xAwd1koXcNb28Yx+H6QRsXBPp
QF9R42IndfgTKUsWCGwX0b1rEDKYV6lOnVlEsCMHeKhYWKcootGLBlh02SFZ/2mTQy50jhUFNuAb
uVRmeIvO1XWTJez6LrQGsJiT1MZY5rTTt5OxHJ/sk4Ss+vs7hbMhev4vdo9zHf3JyIdHN8J2lhzL
bLHXJiPfKro7EHYjMDwaPZA3DiIRsRGgOfFhuC0nfOkIj49fdHbpajuuPHG05dGHSOIYVGtGyfm+
5DERpGpv1Tmn8f7TpwGIqDh+oA7xelNBkjxTSx8xG03Nt3FmJvZfBo5ppENpjvR5hTf84tFIHLJd
hIMKOnJEzQTIIXyxMzd58vEnIVG7r6bxWjGkVvC9D6RDoQ9Mj9CAGWs3/x7eVVWqs8u8H42n5V3q
pXyTLMXRhbqPEJsipW9hxgMWZT+gcowx19y2oVokBvHAdJ7PrMtnyq0AZ2jhzogP/nUOjtebrIsu
6/vFEpe4m3uxvgQFKzrYJHJvT0CAOx2QiWzfTlZwDrFjBD0qpwbJQtect6AwhmhJo0gGTvRWdgXV
kwHI02KC9I/PCmaZ5EqjR4UZ0cQUcYJZjgInBP0o39BQZRuMz5rOI1QKCB6X3/VQR4l64n4lrGpX
dCdfzjl6u1vRFts/dYNe1lKd4R8dRbNMVqRmaUEEVVqgUGGb2b1zqYj8YKTf3TnTaxxnFhiwGpTO
CcktedfiFF4ooZOg45pHyU+u7EB1UAEZ40AJaoCGxHM1iKldGD6gUrCjhWCj9QUPZ/S7XKWayRwM
aZiq8MxZdzePxtLqnEY9IR8H8FK6OGb/j61fS3WMZzHhf2qBLqUZJnCtDaj85yH7iClwNkwng0OJ
bHXRgHg9p3OCP392KeWfX56xYXXmCR9sJazmWz5V4mtvhoNrJdaq8xKtyWmLLiHRMJ7gkejQlAtY
Cuyth8+LdASqiRoGU5zU4Tz07wPNEvoR4nwSobA0qRspP+1bnGBKRzDIDRiIIcy8m33M1BkxQVf8
sdvVZ40RW4TE//nkQ4DIXpIEQDKT8aaifs5NFVW377F8Ty1mBWO+257U4v7wffa/vXXDNOF8s575
qwllaTGZOFXTHyn4o5xa9DKcB23mV6/luMdQQ3iDqCzvaKWk8nIucnbR29m1WtRbglm53MIaUYbn
lCzpZJFquznpBpBqi75twFWPEhT/pLcze7ssRk4FgxsX1ZN5uy/HLTwMGWPj3qZHk0rWsW+mL6ZN
3dKkYiaRcsDS2iM+JqJQVsqmyge7QnCipwLcTwN1UDUrZmL3MmPlkwUSEkamQB+afQLGHMRgAoHO
ak6inWBosF3XQe+pBbb9ATKISjDGEFyD4Yl2r9LMoUg7slEVVBIKL6S9Zqltt9IeDzGvBPbYMS/7
y+t/9nNrHKEJFjtdBb2sbMDKv0oHAVmsitXYscUZjfVUGVKlM9O+ou+8B0RmJ+z/HIpjX0yTHPZ8
B8AG6FuJGfnMaQb1Q0cjE/B0mu293XNxDhsMUD7DmrabssiZ5+AV15VsM5WDAGvajTNO+baWHGmw
fZVKPS9FMfH13rtpWs1gSgTc1/93bQdr5dWEHbhuPuHWwvJRwfJ1qghHDtpOsshHsHY0XncaZtPl
IXseB0YBQhIPJQqJqcOq7xGNin0Qa0vH3jBd/Xc+8+EQDGqARR9z80gl/q5pfjhB9HTqDDWhZsrF
fX0NQzlyxDdAF0icotgKqNRXToOAihBA+IhFDPcL/fyEKZ3aG5G0QLSnc0Pdb53UAU/Wf3tXQ7+o
weiuMVegd0X15d/9gjseFS96D2kbmSH2jrf4McEs+ZHE8nY7fvEsHWbsILprAcLVv2BX9y+2qNW8
uomGTYe5vzF/YZZ0xm9y2skaGlIJunG0w3HCLquV+K/h1srJ2vrReLlLsh/zYkJWIO+1owC9a7ZX
Ymev3b4DNbyBc5jqE63gn2t+4qHe1HaqNZnU+dd5ZXmF7cw5skMAegZ9YVB3ZIJo08CbvSjEGng5
Z922B0HdOEbG6DauYyEbfdpQjbPjEyLpe9u7+6ypcZciGzkUe+BZcfwpDGCFxIopIy1PAN2iK8k2
RKTGEmPRs2ry8AuK1aCrU8goyVGTVGgzgTn0fhHa7xIYsuQw9SpCiXQMP4E1qK5N6yy+EdAFOJKv
Uw4BA4txMku8BarpoSJQvZ034Yw76w7VJ7lxVOZnsfWBW1X/qgOKAmYe1yPdbVhV1hmU0qKnSLRw
Qf/kMqN9OXmvOaFiW4TkO0D2nCTy9XzyLtPGXDM9aZ9UkF6sm4pCyK8VA1/PJ+xUf8IJ5BNwQ8Md
ii6XkG0GOHuO7gv/YRkgvvcDDQ4K9tv1Wl28Arfv6/BPbZCJ9+B0PqYQYl5tcN2sLlcsUzdKS055
Vbidu/MzrsgEEEgmGE52f6NoHUa8MaSNj596AAQ6ton1aIO5TfuVaMcA1wSm0mDkM6TEWIxz4/3g
TxTskhIno4DmNJ9d99+LAXWs+yD1CHpraHkf1zUPgFPmQxYRdopl+rY6CFMNUqxnEhMgQktKC9H5
DzKn/HLpEvjdCnFVsg85mUA6GAawg9vDA+gK550jEbsKBOBbclpwqtI6FEtvuT7uzO/KpSaO7VLT
5QAUYl6y4UGxykIwwTFX57aI00yX0Cbbrgwks8+vbJockMO0yYsk5t/1Z2Npr6S3snP/kF+mygkr
hzAmVkLgh+JgyX1uEkvUkBU4+pP9G2PHq1TrgIvQypqhJTbm33K/cZp/rd6btrmLSx5n+oYUafR2
zmliRc2d2twr5sq2HZ0vNIYkEqKokaPRmM5J2m9d+gTSfKrMdxQm878foCF/Ue3VVGW8gW7c06fu
1SArB58p1er1UmdQNwq0QHK6w2TAqcDUhnQJYe6XtaqC0BHVRvgTRghkG1T243h4y5dmoFOP7Yjp
NF08P2eSGLBBS34dmi3o+FcuJME4dWQmGneIuOcPduwCwFL9wIVgJc7w0xt/dPuYqcKo5hJk8ljk
61YpvjIF1Jvoq7/6o2ERZBr1qXIlY2tOhEMMRjVCG88UZKXGzUXceDYLyO515uOqmRkTKT8Bca6k
mNgq1ITYzodHqYDMPDzx/H2Vwa1jOAun2z5zjb30cZ6MxY+hazyg8icfYYV1Wnbua2BEEzD1+3DN
NsHHLzh2wBk5+gxqy4KpJdwlou1dbVsXB9aSVh88KhP0HvbtDD3uoGHy3D0uwh8TKJdBJa/0Rv6j
UEG63h3JtvIxbSiCo9GJ9AE/2qhddL7gJyXHReANQ4jdAW417WFDqbavUqo1I3BBXkSDUy+59lxq
2L4QdG0rdiUS8A1iHYkXX17MYRXzsdl3lXozQmvgFft2XF52HV0y8Y25boq7j5P3nXhT/PsWs83g
qr/sdZBCVOd/DBqGQPGWqCAwe+z94ABMK3Zi3ZEzsQ45wx8R8G3OX6PZu4KjHJMG9nLUD1udm817
AcPfjqnmQP75BqRF1H7hc6o/HhI3ja7wqA8ArLT6MiQ5VPCIlN5vM+SOWK2vN9h2LmCcb3H0Cru6
90zSYh1babfKu+/guEo+jORuvpcP+ERDZhAqM/Kjwd6V26tlRwa3qMMxH72x7srJIQLHOnw1DcVD
Z4B2PyfoJzm2Zyr0Xy8JM4IMz95zh19ql+MpyEGcp01rywje3kE6S/Pl0YaDblWWhX6/oxjgzAH0
C4CsdsY5NKOsRd7FsR5ofz0NUKsSYUrFMZeQPIbPoLsXcwWAOmRRCdmNB4rFtuk6wfMS/mZnA9Ko
QEJtcB2BQpe5uEa58mQNXZqasAGDAuvlDvSdf6bALKYDAAUuf0+p57aO3HsyeJb7iP0LCSqYrgJX
sFa9RNTzU5s549+85dnXKXv9MyeaMbcKkd4D57Uwtd7jElPUFpjRkwVSV1surBtJDEgtbcMIJDLq
ul3E+AadJU8bmzkepBL/ls3+8R/L5zn1J3BwBfcGG0HaJKLIuN1S7kZktM9cfPgCdIFfGfd1JDBm
AjupBzQpjDV53Pcsu+qvC2h0cvxymA7Zp9he4WHOHXOb99ydV/QXbEIfS+fcaNl0IQCQmfCHWMes
3a5vrK+3iV+YNqTnQOCGyETppBKDEkuU+rQEIXVzwPHibT6D7H/HiK2yM/n/fziIlxEZTfY+57eU
i4y0B1WzgCLxC9M0dh5XCFgX1ZGpLozcsoZcyWpcQhYquRFW9K71ZRKDxrVExHM/sSICBlYMWEhP
0eBFoDlFAhb/VRvZifuGTgCi2rf35e6KdEK+genIuR84ItFisaN+U1y5T5pLpOohCzirGp6DtlOa
QQ+5kx1DLlhFefQt198ePEiCSF6SySaxjsiQr3zRimBUI+Ipwz9V2xCcOZRAjYQ8IKTURBNrf+3H
OUgjtqSVgBHNHx37/ze6WnEMSgmuYB53uesM9WPh2ambi9jjpB6DjnDh8ycfLMCBSYuw/BSo119b
NDTadlyQT6jNAzwyXBkQ+mYn0ElQxDBHdwVHvZxViaWOGFFuhFolz1GhWvCjhSwYyK9+GWPiUyhc
orprz2Edh8G8zvicB/0w23V5/HCgFsr+XcYY59J18tbUgSMvZ5O+Ui6+AG3oznhPuVodXJwSQRQu
7QytmyIexYBLvCzKCilsSmQKaRCqr26/NP3Rb2zgt/dUrKbtiUc+yjpOAfLMYNAR9Uig0PZXNnvC
mwTe4qKL2DydorCBwu3keQzG591LRf8266LUBo+wgv1DmLKkLj/b21NNJDhWrSz1wNrlEWAOadey
Upc4y6ZiEdignv1mUmor8F2vED01HOP4GfPpVSO50CXkYpOKqAXd+un9Qbc0zTJGd0uibRM+LOIb
b/FakpEe07iGTFCRfrCyvgfnqRwvMZPui94anajBOaDt2OTQ6aqIJs+RTqY/nJzOTZ3zTr13mrFk
c0sFnIiOiDkZpvt+h+4oYVTMpOurSax+PhGj7A4qPA4X0LyCve+jmZ7lBrFPH01eFe5J1usqwoUL
sHVXklKQBliUPAYCo+6pxk+yQCtfSKL+W2vPPS8DDF6l5hcBiRlhfSqSxoUDmfmVU+JoFQyDbvVt
/VB8NfpBgBRW8vOaDi0cZJDY32QACLTZPdr/IwipSuW6uW/c/gg/+vq5Ui5J47DUzyq9lwdTnDvo
3RFJTinah8v3tG3uWIen5Gpf7mi86/Gf8vFsUUO+dVRSsKd7UmXxqG7yZqMRPeDeCjcIJSGywfFc
wN7ig+22XGukft6Of0Zeu5fH8cr8e28cQtVIG2jMB1F7f04hTRTyX6XLQt4grU+H7/MNvL+aFTxF
jax53xJCWFbvuf1fugIRMvAc1scErSDFXB4A59nYNgAk1GnK2gv0+xTP5R+J94fojzfaEQQON7YW
PmKrezIrK+VziOnun+rh2tR/ydJ0MVaFQPccGfrjFwTJkmvxMf6TE2J6XIz1jgvYNNRc5jg6ZiFl
BpvIdg8/WOg6lVB0KQn+zkuRUDKuxnnCbisP8oVJNQAKOPifOjNt5AWKnROhF11wri+MU/R7IAVH
wuwROaupmC4OSchy4B+Iyej60HVJquABWihHHEb3FiZI1N43Ku5U6t74lSVqoEhpD/xkQfzt/LAZ
G6hTkMTwRUz11dFCQDc59JUI4kpL+OeOKBONySLEn+pAA2VqjAL2ixfY3VxamMpM5dCYjhbdNEFD
7fVVGyy6lA0zp75PDAfaajdQoaPQb2x5EJ7S/SGbQp4iOGIwl+kZ22+uhvuYYoiAFxfR/n66hLWx
51t7OmEWsSzQ/Eu8tmFzvY2dF+8t7Uy4n/+ZRmdqT4BBBzSsGEvpTQuQUVPfBGMoRLcd77i2TUSg
+4Hf9FzYP/WOaUZ8N3K6xwPcHOI7TBlZGam9ZM3fLMfoz4WybIgncWyLsb+YsUYDsoRRMVmEvO/8
qOp7u0NUFOBjUV2SgdjFOVdFF403A+lqHvThAzz5w0SPPQLayYY5aENp0OYqaZgByrbMx1DuJUzQ
Lxo8LQ6XRhNVCvfH1VRcwmOINFpeHASGS/1G2xTFRh746uJxims/FshDsoo+kzO84Ytu6oG3i1fM
bbKU9zMEToYMq0RsZ+YTT79qGZFIWNHPjlh5AFzQQnzOVQnj1AgItHKdrO5zkfywTBZjdK/VgpJO
EeE5pnSmM0WLzi/hSOHLSIFOsXkyvSYvbW++MGuEnzin+neFE+cKs9uLzsgGstnoM5t/qJ+jdzqi
jO2kaiEQhg694W9v6b0eGotVPdj39PEujkttduXGbnjHsCbYvz3/HTRDlCANWHvSAxYxjOp2Ji9x
AMMJ0TVdbs2qJ0m4LgbUn+MKjcwTnBpVmIi6u+k2byGLTOdbVelc8gj+s0Ul47cDP06WcssL8+c3
viMOslqvXr1wPneyiJ7/uWbv03txoE+IXN9rpxGw/9hmax2bu9wKV/8uhum3N5C7jiE3Img9pjnt
SCYNIBkzHC2DeVnJ2KhFsToa62Wh6n2C8SUPByYl1j5V4Rj7krV4VmmJaVGFrzyLUUW4lyulk4aT
KFVsKGFUvmKXWzahT+hu3po2zc7bBTv/27eAzTLD3hpafrmgdaeN00o0lBEGIH4lnxJ/3CKAoGm3
A9vP3hO5Jh6KUwrwp0EyYCK6pQ77KVC3lylo60hDtSD7SZ7V009lXG3pKsMVqjf+3CvIlWDKwE9A
PnRLcTh8frhps7+sbUv6Q/MJwVqgrgIkExiKKryrZeRlDVlJx/bhzYyA6HmJGir6MSz6rkl8PptJ
3T4/+h6t07N/AngiJnHqCTtIPjYDTonILOf8KBtTpgUWDZPIhFAPu+658InPV3+qUwDFFOmy7U2A
+c0OZuaHSlwc7gq9BsaZIDNoSJMjpdVLKj0269nSfaAgm4/LlOnW7JqX2tvRZ4SMPXROhiukrD7j
mbdYGgQN9Ny7N0+7ltj1VXAEDC9mhoK2SM7kruqHl60kpf+Uf0aftJYlYQAmXEdtdOonF0MIRHEX
ryhXZpVbb89yKSNPupq366iHWcnID03wc48aL1iMPYk4v0xa15gJ0oCo7g4b8Z6sERw8wcFjeFtZ
eAr3aWWaEfGSldnT/fY8Ft97aAhJoM2n59pw6xbColmLIF0lLIk1Sqx0ggM0ot/5v8ptasWkUEqg
r2Mk1AJp3mIbZXXn+28cwB4fCUcACQNAF0IxRd+6u0gzd4mPl9ZgX+18LdTrMPb2uIPuOCY2OAeB
VEJQxq7n0MTJx+t9t3qBO9VcCvw9N3o/L2O/+TnIhDhLLbUSZikyNsEHy5rx8Rx6kwpvPKy8c6yS
bwLpFWCBT7pT23LgBB/dFDaZffL+acKLtgEZQ65ZhSF/FMDaIciXcCiIH2rfsvsWOd8OvIprRX50
PfkoxD9PfVyqi8ASVsUfAejOKN4vQ7cDQN/ziP1WBiZhYfsvFD1L+7Pr7nvnFBRy5vkgnOwkqtax
P84iEKuAcILx464n/dUbqF8/lzpvzuJITtvLPTEtyeiiUwi2TnznYQyBxGkf7W1LRLY3NMhgoCer
LXBreAiVu4ox23UD4E9EJXiyspLUJFunYlBDuD63bsmVgoDY3DgVM5h061DCT+7pfSKQt7X12oy0
IjZAALIcw5dGFop4i9/71gRPM9ziveA/i0d+PBJT+E7SSoHqLMp8RwSwzChdam29/s7ulMKsStnz
ZIJ8HcXgVAibE6TcdvEq8MDegmLgxmZ+BHh8NdnoLm9wtI0Ka4GNOk7rnWS7kKYcaCBCuYGvD0b6
NuYz16T5FlyhBTZL8H37jqqw3fThvIvn9Knd9KufNtDCSPUxkyUKZz6CmfbmQVnO8EPrSI7nI2aD
0dzERf767lmSa2lGfmiHZrP4BW61O40ScCRvfWgIo2OXjh6AhFvrF9mEGbK3qnvqfBpHb7BrRzwT
PKoiFHOIvXvszRdkfFRvBcvR9bPHGc3yjncbyXnvY1dCiQI9FMOpqcCDiURckVySbHDdT9UMuU4M
VWO1dsticvSVtaRFiIeB+Dc1NLO1+KnPG0mJF32gUk+8gIbIIv36AOharQZ74HS4VGHlA6GKYllo
J25J3EekBAjXrhWx+76GuUfokgFr/86p3syL9HAN9fAhpMk/BqVHiUYtVLEJMhuWzvAe03siwB+i
otrZ0BQR0yf/gJM8kwRJWzRhHOwY62E9bwtKJl6MBeMawrOrwRZKOQvU/MQMz6uLjpqMwIGa18gf
8ma/HYehUQcXkbvNMSFuuGhtHC/bOCLrYLNYnZvzqompZxxm9ryOlaM0AKOL2jci0MGNIVp/tTLF
7PSGqpEYHJZKOsZ2OuUPkGFfo9aP0jgS+QoSipbEvebECCQSdZMzk7r60WFrore5hG0XR2LnxL2F
fSkqM4bTpIJcWDBT39iXzqVPVaBRBWpkFgsKEJkPYB1CfYyU8cFDqBdTjkciFXj0BEDgnc8SgfHe
4xo/p1/scTOySAYqCURO1ay2s7RtejvKOszcZfIpLNIt978qLE9iBOAnW6Nf7ciI1AJk+fjD2VTf
mGxkx+fzlyoCuvO+3JxRkehjcD6come/SR2h5qkUpUtvNuusX9WVEaYOJeJG0RJdW1R5g5oc8vQm
FaSz4nzuOgNPsFKwr/Fzw0zWdD+z5Tu7zOHBG/d6r4yKGuNksnyQOG9Jzii2WRNh6mVYOyf68w8H
Yl/Sch50QS7IHkMhnyvDerH0OAMKWe1a3F2UJEFN2+KkQtoN1QIjdbFKnJzHfy8c8UJwX5zZHw6V
E3AbtNYUqvkYHT6by+7fR16OAjvOPHu1vrPtnoI7JZiAbshSvKkjhi7T2NVN+gUTGIAtLGGDAUbo
WHN4q4++X7FDMNCSvfGd6oJafsAx7LRgVKhlgFVnZHGNZUejsA3iBbaGQL8afPU8xl/0hGLBVRHi
P8XthfQfcV8VmdB24me0RTkY2Bf4EDAprvjdJQT+xh0IBvElKp8dLWmpiIAdmUxL3gVLWgLlj1oB
sFjFYALyRPf2pZmDdi7hkGAzKVEvwzSDcYalvJeX2w/X5+MZWfB28Q3EjuE+ZcJMjxZ6XBPfpiwz
5omcNDxv5+DlIEdTGUfCskbulQ35DL3+54R2AadacNunA2zniENY2P8rNhPzBVulLK1iEBPNpZ9D
Oy0SSCoF4vpKjaMqkuyKQqd0Lz5udx8BJuTSASW1wy68m1a3WMjtimQ440gT0jVsjov4LYmLSZWs
C/6sZeYyLxrvLSOlUErd5MsJMpGlbCWbOhEzxjoCbe8MbSY4NdVs3v31nWu/JVlGr6Xd+UfCU6c7
iMw80yncntt2Z1oUxGufhxCy0gmVFXFJ81giRyRGN8J+DNl9LaHViIt+tj7fcD7hZqVcPahXBexh
eOmjQyNf5krooy3VnOudwKQR6/zPx8xdvJIHKDnSY5EGgRBjuDwgOqVZ7AD1VtVq4zMI/CGUEZ0+
6nJgOMvAcmBXrt8A+9XHgs1NhjGRciJJMo47/eSs1SsEpQYY7oAXHTEYisB2ZTE0Q4GQAW0ig12G
OFthttuNwKt5mCtFYG4WbX7EaC3VLLCZJJd4tunuq21XfR03aYTMCFOZQ0u9exuu4bj1m/ED0CWt
vLHB3A1FhEGPyD2kjBZG78HG8PXY1jRmgo+iPAGGqk4pPu9bePoqEcWHa9Nfpri6mn+J3xtNkCgq
oltusBcRmsLtUSDESXJgdBIXMJ6WpZU0rzS8LIvnuGLXXo4P3Lh29x77I3Ob7Y35npQuvgICtPhW
P2m4vkFjLBjsCTkhTunG++502TnmDk5h00esr29otTMrGfcPK740/4nxoTC9fmSqx2ZfCsYbpgeb
BhHS9931/JLZ2uyEPKYqXydG8WpIPzi12z8OwAH45FOG9y3BPp/aaqA2OP8rKZ+Rd0hEuCmLpMHO
PV4sj+t9/vC71H1Kdt2cP8ulZdzycPA/ZfDXcXBBl7ie/DDvtDnL+m8iUpmTw3mGgsBbXlJ2t9UT
dEqqK9CvNgzI7txE07WRbntyzJXGimPplLcWuMvWkDV6sgZzAXtmdx7MzO9vHw0DyBofORhRA3ry
qJ6xGaMszkDEQBbAbAaLa9npSVQsbRMrXhuuXQUyJuzmWHmYo4DEtLG1cfe1mFauGtppbRmGWjpJ
/hpkeOnoM89LnIINvxhbpnf9hNINqhUE6fg25GMoomd8tIcKF8s5i48pxJ+fQoJKEStMO0tzIqUV
DV2zllKhkOLbJ/eOuPLZaCvdsqKyiZDu6FfGcmtMquzQKazqW+jlA+mX4HJoCkR53pcpVilT4lG3
U2f7qfepDAQe5gn6Wr4AiQLVCyj7zMfarfQ9Uc0nSkmc7bHU06NWPiwcz6pce9t195hvRmlaE8Fp
MUgjQkl3ft+lzcIyeSnUSgB+HRJVMn9i1R3jV/12wpkoQasvk+q/XljNvsJpaRbj0bhLeHZuUq+n
7p5iJ4U6KvTuaYmTaOw4YUZx+fyH+gTuA88nRGCPc1ZOISLtAzt5xsT10GofW1Jv8qSzhg1NsdxA
ub6DRSkU281p4s4VGY4KY10Fzp9JSGbZe25yUa61ABkn8ygnUizqCE5ydLWwAdHDrS2AEw/2TvlC
7LngixmqV6tyLTIvF6IQwSpMMuYYqWkkqgztQKIcMnxgSHYFb39m0geN6pT/JkyjNAbcxHjlQJN8
k9fRxINAi7mCH6+8NEzJglSaQGG9X2a65gT3y9opvTXZwLpylqDMKnm+mK4Z9vq7r/ddfwcPRn27
IRtv4LdEmPkgkHfOya1sUV8RCp0Knjydjbt8ZJdoxjvGzWtCWnuSfmCh46bOFHDgqzmOQ4kG3jHL
HQKit5/r2AGjxb1763HEUSYmS6QU6SafcOW/ATzAqTFyNF5tL4FBvbADCbfU20+eX+nvVWIZypq6
2jplfjddVWS8vkX2dZ2EeHz0h2EDId48bHN52ChHtYX/vy33c/6fvHGCKovDa1i4khJP4WUyuovX
qjvH9h7ENoAkvPPjHooZp67Ks9GzAFwJNAwLj9N2eGftPymg6VMzJzVIY0EatvH+LMUwNmrIdgNI
7oTYs2O/wyaljZAZgECsr9jESACapOqb3flHzXVOszbdwNKMSp/phbAf83RdjxXj2N4ozge+J5Vb
bEkurdbzvnDsT1JuzSXtkeXmr2mFnWLKcDxnO9mkxmVIG0X5bzrP3lyQAAwPHXssu3Bd2TCYrW4X
pqgQ1ZpzWt0aVpfvXSiv8RkGohCvDavfcNptD0g0FysIcd3BVlpIolyYy4OOS6MLRoeJDNjB/CMt
WdE5DMxRiDoSIORISMXuKCsZ9s8zWfNWkTNM3j7sZXLNngdVYNSYkxFbXeIpc2OH9rRjSMBE2mGo
tt3SuvqcVQBI2gl2WF6wQx+nwIcKYSNH4WitdOkm7Fena88KNq8K489S4mitIgtzVNMzVbYFikrF
p3Zmnb7Bw04zAJa9ktDloSy2WP1j9SeocUDp1ttpn4eYSqcoc0sBKHncw3C5NT/j0M1tsOmcSgCq
BMTsuHR/Twv64A9TeVm1tROAy38fMhTzWLWMUSsIXQXk6ukwAgrVFgoCTv5New2/bDbjipEkDQCu
tWYZ8I75qL4MSWN9G8QegNcjeGk29gRCWa5++c3fPIInZE6FZnYrAt383Azlk/x8uYxdbUg/cG+I
lZ3du1E4VJrarACdTyuEkZNzOHg2Lm1E8wOE9T9WmAsbs/sfIIRX5xLYUMk//9DDf/fjXwVvqJFL
qajfVInTRar3F3JY3TJ1X90bkdGRYOOiuQrtoy3DdixVkFovEdbTpPyZ/6tTQN9l6QqVWP7FuoRL
Oc1bSBmEAjjdPNO/2GoCN772gtOHYRREZOBLQU+D9kJGO9DddN94e3CcxhQbZ6jQOL9WN1m+7EIC
Chkw3x+INRY6TJvz4LBrTY8jh0NbqWnq+oPmFp9/2OS7EwhcPAXf/md0c8qvypsvw4/+11Z6g5Ol
5d5j7fQHWmbVb5OW2DTNrrTTDAQrzok5NoaKw/FShr+AoMIo3z1WltNtkKJZUi0w2J1Mn9xv6a/w
8+JZYabV+WyOyVs7QLM5u2EHYRDsKYR+E/1RZZyAPlupkqkyWiw12SZoFF8A5H+IwTdC7zEveiww
2Ta38KkF4trQGi1gmKnaTzsp7j/y+tv/lodu5DdhGHb0F+3jJpdKgVsHMUBynnfY/62xYrb4fyfe
1yuAefvG6IlFxzJeD7Zv5lnkV6sQtB9cRmJaXrkTmSb9MfwkTJ1dkydbURfmrqfO0HHyLnuAD3bo
sGAI114D0ezp/7O/rL82Nd2MxI+8T9g+70ybx6dRP8FFT45zQ2T2kX1PszRYm6yMrHynQxRGXsWG
4Z84pjDNBnwcfAE3lkLHvKtkmQJBe5VFB6EfTvsVEasXcMBvg2kLV77u2hx8WHujSomfKY71WoIg
xHEXB0LBlVe8rud3q57xQ+wV0f6vbLo8mhvTsF+vSLx/KA5FdiGkkP/2wDlPvs0AWjePVxvWW9Kc
F6oPtdFdoAw9nwjuELiiL20vv3bUUzGexwGp/m3wtppEDeaAujUmd+mb8TzGVBoTDdhIDrf6sqqQ
GgxsIQpcYd8+lW2tMguo6ZtS/HT/nrj2wmtHBCbzjEXc0IIpgkXmszPs0TsBPxIMXKYGrC0zNDZg
l8PfmqCP5SotKwtXb3ZvAbKd4TZLyyIy3W9gaRujooIU8xwxfqWlNx82OINVHu15zMpGtkVenCnZ
1zx+tA8Gp6M+s8t8YaBg7OMpGauIPl7WrUuIEbkYSupCU9ntDq0nivYTsi7HN2CaRHwvxNtsvuO/
K2Avo34OK8zBdIqL3SisIsfZqAJtMat3Wy5xjcEe8SfLqP/+8qaU1EiCm0tvFMfYifucWz7EYJnV
oO8K/N+RdueOd7s2R36lONr2pLVgp9yhU6Yz0Lp/5a8eT4mdyqDgozxjwZ14KxShqIS/mlmtZ2OI
WcBg3kefxFrbTDIbk1xeYoHln6l+sXLdL/ZvUiMAoSPEBUTTE52GMkbViMqrlR8jwnahpsE/suY+
LBld/XzVKn/o5rDi9Rwvi+DRvWwK2SnIqPl0OIm0IFdWBubAumC/n2wbz6Ofq1Tjw+HDiwXDLhRC
UfE4zf27OXDfMmzOe7Z213rXKwIw1HaQfuoE3vcbE4HjVLqav+Xpb0+xwDDZzsQa4Z1BO22d398E
aQ/TGJWmMcDkuijZBbgfNaziuIGQb8mrh4Crxi99uHBgfyQ7adcJd7C8ZJx/hLHx/NoGTxfcLNOn
Rh5bCXKYm3cih7wE60swR29Va3JOkSjLWLxXbnyJ0UPtstkPHWq66K1ta/inv+mYrmkAgq1YSFIx
ebV3LUNkYCWBIIObS23m9Omrppm6bHCKuP76KIJancNsaCsWGGmjxMVglTZl2QJ5oEf3CjSU1pi/
TQyT/vo11GqgZP1DOO5Z2Aqn+FBZnDHT/MIA6kWJ3+Fe+1iEP6rDvIZKirH5sDiABOBx53kB5H5J
nV9Aqdm5nwZbXEnQDTv8DrHvD38nGxPXQUcgF3sdjLF1latdldHJSQm+wxEmLurLBEJ6BiirLCs4
gzkFdDQLumOZ+KmW+g3BIE9Zf6PFduDD5Wu80ha1MZqgd5BEekafSp+ok4mVvpbLCbzrhJwLfNmc
+eU1M5gjnxBYe6oqzcKllMCOucrgBfJRFunJ9k1xDy5uYsN+FXFV0KgkHyW32SDmNY81X9KRek/f
rd4lu7D0fWrXky76XNt1DhBFZ+0C/lCQ8KexyAi2EzPEKZwWwJJA0AW6PCf2QCnuv7g1UgRl6fSH
hg/0jiqnF9tKWQ73Q+HrkcQOFOtvj8U7HlCOQhoB3c4MIBQ9Vg1kinfe914iHPU0SaPG8701LHry
L59rKb9MGXwWXRYMjOIffeavpYI7If0og9il/PPVfbpJlD0qdWzyC1dsYnddkwhhbhpVqRDA7yUM
jT5rMMuaGHnLLdqCziw2ob9/T937OGQNlard+jprO7ujDh8LWOx/z9FyBZAF5qnthfH7FW7t54p0
+rjsQenWvtfSpGrTa0B+hCGMgPDWdfBCNhbVKWoNnqxVMkbx6N5JywUQeHcPUEVUXkP6R2Q/6alA
yG/5uGfQfImBK+mm6zmUh71WBUqwpQARbIOXej4jpvGpj/S2pu++9r5sXRxxt4bmQ+y8RqWCikaZ
U0suco2Qd10JkFrl457dJsbIqrOK0m2ZCns/JXCEdzk+3DRNnHRuit45u1gjVUgYo2xfOjvhHEZs
fHHdylOFpZxkMBaKlV0kTSly7/MhGf1crj5Zqkk1EXVTUhOX/vvnwnuYlhRn2813NQnmp6tyDHLn
/sccPi4nhTFm4nx14ep8ItsJauyztVYkzCTqjmCJVBbuwWYTkKM2XZUllD++ftJMfcDVtCFdlnS3
it7cZ6A4QhN3AYFKTAB1nS0W164Qo6hrUU+JLChuetulKYl2JiNhUaY7D06CWZtiVTFJYM/YJ80B
8wtpxnBoSoKQbL1IDkfGBDiPj8HuSGaQbx/V26Ey9sjXk6y5CqQrS1+U7dGSESNeRIIAykU4OEZC
LbSa5niKk5mvb5jVi6QlCUB+JlAGZQn7NffuqPxP/8OLhKMK3sCkl60CDWQmR0vfG07S3xFW6+iM
1nmQqcj+4pKIAIZtpRKH3L+dqYjIsYYg7Y1VedAMJFT4bvDoZDA2lQZc4Aus8cvNqORqg3Nm4Y+M
Z3F2EniRF0F+66bKgllpxnc3selwdAiiLFcOzbMJhrlY5oGm6bY6SaLLBoT8aEZhWr81KOao9WLB
nT9cltaVSJhti+C/X8fLm8UPOKVXFc3F/1aQNXLRdLd42bC5DFUgDjjrtJ1QVdVsIDhpjV+YYT29
+L/8gf4IcDPLx/bfWrP+j3+W0gjVcWjqejWXc1KNJJjpPX7L+bEE/lhU1ddWYNY7agtvRpC0rF4D
QDXpruK7x448dN3K9zY2F31FvnZ6kH00g5CoAE1ADCx8tRW5ohzSqt3NHVXoUSNdPfbN5k52jBN4
5aN6CiymK2gc10unKO0zTBcjxjGLiEsVjOs3UfTYq0CZEvyHhf2btuGLF0a5NxKdtnJD8UvELcaf
iQ3GQ/u0NZpI3xq57/9ht23Hz2lEd9LKEvk/FrawDE6gmQoceWHTo4Td2jFImNrDSKYAfWZR7F68
7Lh+PS9dYP/iakg+KMqU41wmI4goKs0BH9Gju58mdt+h+mIjA0S60EOOjLTV9eryySH/dw+/oyMn
9fEvP8NRUKqJ1Y13InRdv50EY6v8rHP/48b9QOufjHR5ByUQeBa5OlN5UCFN0hhZDSmIe5w3SJVn
buuJUuis4KCs3HCJzNoKbsx0Tl2JfFuP0XacHadpT7IK7hewCpCPZdj1Sl9Zv0VvzOf8zjQ4ZHXx
A1zUnxruuFrezfrdYBV59KzPj3deByB/6OGulPYwqCEjYtEdNI2UNJDcaw0MYLMbuAQKTiDn8gh3
f0N9TtZFMBynd6EMNn7Jgasw1CfgcmbRhHHz9cLKDEOKUpFpMvcyqPaGc+L09GpYKp+AI/AqZXa9
loEnPmRYoMiNzqM+P5yBei50jSDQCkWPUx35Gh0IlLnDfKqsmQf954WK19F9cukhCEVX3jia3JqN
+mZPjWp+ziZ3BxpAWz8HQ+OSeG8XS4C9+01jJnqh0/UawTOAfmXmit6Dc+8zQJGkQp11TkpJm9yR
4MxD5SCO5otYK6bmapFHX1ndZe7G9BSob0/CasDqL808fGPkObNTmJ2Pk8Tm/x/JJQXgQO6zX6+B
aIJiLBbgn8GwGIvEuUdTEjwOXNrEWedsp46+RHxfnQrLyFXgMci3LZXbNRZcwQL7a/qXQtj/OmVV
kfm3Ojse3ZxgX+3PW+ac62HEOb0wMRH3lKYhatzBi4znpbFDAB0DRK+Y/61znq2qSLNBgB2414zf
K2h9Xu6SJcHhwjODNjBAx5iQ4z7m+Fg83AezMuzX9TtRZOhiLd2rP+LAgSH9LGZod0nfYl72iTkh
jOxzmM5TXOstmamJN4GrVCV80eg9Jy9lG7oVu0DK2ILhooOX6QZ7eeI+RXhZjpepElk6eyM/AH3i
O+qplzHji0TyqZLX+nlixO5oHVBym3K9pBgMFNxFGfDWHY5LbbYiQ9uEwNvR5gcnWOVW+c+BPKky
dGUDTy0EzZCZjR8OTISkNxiRyr6quVkMx4T0E35ZmyIO+WgHyul5lUliTIhpAXP5SXW4A4rYh/EL
TSlxkFGDZjWrnckPEzuTV3tR07yPLx/AUSxVWO4hGnu65KM7dIctMScf4G4T/V9fMoRTjnOzEgBz
6Yu8ndmr3DQphMscJB9XfUtMx4wXEJm0CoQyltadCXXcixgecV2+5JK7LrTMV461bXvzSgca20CD
MaY6L5OU3d1WZ+xRn5oumC3nkZvKlq9WDFigKIVaa7+zrIS4KkRayZcBa24hvzrNTGFZYLKCkvhR
rNBqZCVanuaFMOsIszzhLrCxM6j3GC7gKxj6FdaDdLjhIwvPLslz7lXCPHVTgkwiHj2O1ki64RPD
RAwGK3Bi+4nC6AjlzMtBis2q/XgcD777p4YGJbxSGonO9pydvBxfJD6PTs+6sRTAUGvNoyP9F9al
zsuy4W7uyT5Mtc6r2fuSNU1PgZvCTN6pwlDO5ExV2jElpJS/vgJAKS8wUOCr8UWCG8kNRoJsTMUE
+lvSCCQ9YNlAb53RBkpnljrxUfTpyTW/cOfMGzDB647eDoy00haerdwG5KkWQQ+glMHySCUe4r0i
WxYefBXxB+XgqZauVPyxiK7O4XFA0Qr+AhrChY88FLxDFmHHMPQ7tuZINJZRqLSib77xlDs0ULGw
XHIjO9xKrNhDWA9CVE+xcAgEKZGSL77SjU+NguRsEC8h6Hq2dUTmwaUzjHupYflJq/pKH7LoZYJj
3JkYoYQ04R2UkVNvk06e61rVwx/6gmefUVDqtK/dvv48v7/yfSmezdjrGt7ccakPaPUN4+4N7hgW
nop7F/xZz/6E3QWqwRAISoWatCsH4BdC0gCgkLSJKt42NeMoLhWIvPYcJmcFLLvlwQu0AVFs8Si6
DB+AvBfaWv7N5iQTId/8Z+UvH73K7qyS6xxubCZkgxDumByv/eCI7eb1O3uNIM8CGRwLgn7I7E6B
b4e7RXb/mkwyW8HDhnbgKEt30VufIGjX15+TPFKooDoeinkCDU3ApJkcnqX+y2jcuKkL6l3gCi7W
WQvAG6WXgnwAkmHE/r2opIrIH5GGUnGeoCy5rwBjKn/zPo90RjNvTrkzjpuGQ8RqmO9NISdbYjmU
d89XGEuU4EH2Y5q1DkSlKIET8dnRTEVdjEVkCL87b4q86y4WpzcczNEMvf8XNRb8SEiKyb5zW6Uf
P1vaEYwLnRFfh5VFo1r9FOCst7ffZKdWx0XhMjwN+9xLzxtmpL8ZmChsxKs89V3g5+ZzZeLNeX3O
C/aUZqB7GqSXDBtitVMLIoVKBSqtJQ6oSm0UZ9C05QJHr94Mh8HXgSWLMJD1pFilCw9t3FlO9YiR
7GI8bU2Ev7wD3DnHk2NVhl7TojG6AYQ6ZCrA+YqdDMNwNyZofr/NV261n/nu9umSkRYSTsiCajBr
U75i16/zS1l2i2ZL7e4enjtbmMK+u0+G5jAzuqYSK9Nl6GReKQ7+a52y3/s8v6BiUp1ViR89xhxB
YwgWGAPO0Ha5zqc8eYQMp42hLeeYMya9LAN09VckLqBC0/CNj2Dp/ggSQyKRAp0/KctwUwEdfW/d
Hq4W4b+/OQ/Z2zzEbsgh4Lgo4xR0/2hF34K3CSDIStb705/StmACyK2qX4zgMvin/wgmc4yVJDzj
TIICvaWJWJOGdSpTs0PYytACN9buIdzll+2uk/92V/d20ZzHfVBiBig8lc06EFImaer6QiqMLpAs
lqgMTANXazbxR5P2CZ1uClSHa+D0Zk0PRhFlcFJfcOBrFo4TxoFXgkrAMUM/mE4I08Wu3HsFKIhs
D//Z8d2alp4DY5CZLm0Xv1AhjSquyIyQJegundc5cZE4Z/54vSkeTw0CK8cm+BOKd491lNhb9f5u
994RumzUsWQn3fv/4zeaaQXCBflTu57dgyYQ14KtMiq0DZkwMPNQIaM4KtHXPY7DN6gO2IevoTcM
2Al9/mFxWm/wUzZvO80dEIDZwYTZbhdG3PrvQhP5gGmsgaruQqqvwnJHUPyJS12NJP50AZyKpwUY
gT12ZZKB4dkg+W3c+G4UZ0oC3x5Os/CTw0sYLiz3JsacwAP+/wY6YZNKmBmulNVOVeKxzXwveKnI
4/kqfzihlF32ZMmccxgng+jxXCalFSz2VDDvv9QPJkfczPh2m8tLcX8JO0BN5poJdRNYFhgDI8Ov
l7c7KwGQEEanG3lloEwcDEF7K8tPEV3KTkd6ePyFKsTC7XTpA5Yu9dfqyFfJGWTXd0+cAXSIOQYJ
wvOm3foucCqf8To6iR9o3jL3MfSzGdWXMPOPkWWeaT6g5ldPYU56pTEw+mSZlZTSPt5p0reWpWFG
xjFTo+xPk0EjR0hviWlh6F0h5kIv6HH7uRSAqjVoVcXvaDA3D/QKkIFx5a9XCtw11AK9A6LzDeN4
vmmm7+CK/5chwIJ7diDYCxufJQM2VrgXZyEDM8cT5QMaBa5HxyJMvJgY6GIlXCb/hBE8tniE65l5
U+tW2m8A8QoW/uPjeABVam56jCnuEBFM5Jr49CWjGpzQm179g8Kees/MJu4ixbhJTmtGQwbp7yUH
7DGDCeD2Xfl6OdNHAtETLJXFVCYTgSg6LKxfXiV5GHJscsVmYgoIw1BkAmuy+4ENbY21Cqghh6Bc
kV3qc/DLbg6RZwsnKAardnixHnovFKauqN9u2slh1AZ/quwn5JbZUuB8qqabvwK44iVLdsClp5JS
cz9PcdQEDklsoQYKVA5QJ+lALiQ+kwCJJ9u/09pp0++KIedTrKKRcxVjqNin0wI9an9izZVBP2LS
tGp7xEQSAC8gZNU6UqB1WMYQE38EL0gjqCkWdTBl/Upe43DSS1LF7aHZIHHjXArDmA132HmxEnmG
QBkbFs09Hl0UQLjxdOxREYd2pFEouVtk9XXB7lXNA4n1+hvlnMNgGvkrLn23yBcI7yBjTVVq1w3b
1SaCMKDDuCihpN7A7tHCOmgQnDCK5oCnsCS4bjE4jQZrbS8NEqueyLIik4iH5Un+g43e2uWtIVMA
1i2tkNxqMdC478r9qcZTtdzJhyj0ZlpPT8uNdf3dPZ+/E3bIrK7C9K5qgTfmaJo3irYPQ45MjFEB
FghulUxqh0ksdyiTFUnp3wdp66z9wWxoQl0NFrJ3DeN9LIXlLJHje92nMCxdX8XAg57LxoroeUOI
zdl0IalbW+2hfTPCkfF6QQTWcPLoMAegQcRmRpIZx5DXJEX4Nm9n4pVHX+46taaoORxshhBSqape
1Bn8oeKI+jD0fOgasTDg6pXModCHR2paG6dqDgpHcgxEP0Ncb9MWFiMfnJaeufQ7QB0bzIPj5ZXr
fpl9HVvxktxDvcR9ukm5Ltr54fDGzP/T6jMKArqY0pWiy42XLIu5fRANwfqZwPKEwVujkcRkSPsH
7JuMHo5Y4dLExnhrjoe/E6xDZNdqC2B0EaV45A+5rSXFyere/GnMmgHwQg9ylX7Y86mKEdpQYrME
eEScA7Am/ikRfOZLiZ1VpI8s0WkYmmjxpsirrHHDCs8LQUSqqc/H9TL9ZiaIp8tgcqycqQhICwpD
ilZsrguaSExuKHIOLxxxZaxA4UODWZf2TE056UdVbX3hRfdzzrbrTaM0OB3s6cUY4yfJNHZI7yM4
p9BeP1VmjvotnTbCR6/gjjHnRkoLLjFbp0KkZGqBzAp23/bKOHJ7c8iDbcCucxZ83wX/G4S3b1Cz
UxAp4xjYZk89q+LElWQdmtk4lzQNcyy/ChXDuKn2bChSkYZkFbu3lIzU8rMaVX8hVwBkfYuIaj9x
X7DNBVrJcJ/Kp3znK55A0WxzSTjwE5mHN/ndZag1ULauoTJnxnnyfpG5/m1Mag+7nuibHFde1ozr
Q0UD3HTDFaSPbBRI8JpJU264SiJNPk9jWcwwaOX2EQhkc4V90JbkMAValLGEsoCOGN7tvNVH2/J/
pdie6xvqFftfQ/uRhRsh2upTa9GSTsymx/Uh9Fbll6JDXK4/pIq69ZqgXAM/jf9B2DlsWrpyp2uB
EWm1bsvZ2ojBbKej+GTmJGtFlqz8z8EuZOqkqlPyCGfg6nwzWBfFuQj+ZQz9a9UMKOLDBaoRNOZC
PwQ0YyFDhArTCQdEFxfD+LIVz/TYldtsVrwWf+D6EwrZBySfhFTSPUqcUyHkBg3pmw14hx3iGCzl
dczuKco8BkGvQeot191SZZ8d8TVzvLpTyy+7PiItDLS/dodauskUC1l8u+HCEbsd5M0Zmh6SKqne
iGTVq+gH11/Jd094yr23dlRhTbg/R7rh5k8W6zWkZVEehZQhOu9LFK61NUp4M/eKw1OfLCsVADi5
LIYAy7Nvj+x1PXIJGhmz2iX8Y43QrVn9hvTeJR59J1CgCuJKP8Fx2Ijoqz6VPfMyuIUuo6by1f/P
ZNyApVBoPNC107WqCClMVgDaMmYBaCGD81YduxbD3viF3dOCW3p4a8tUCdjWg4vdvKDkMQuSjB7J
BM9vvCy1FiZDWAdbkcFsaRk6414/8mUQ1Gqx67pCgabyL5l61A1V/LlctdIfCWPg9ZpbptfZWIuq
57/YBT27Rutb5FYzvHdDwOlnSpI3lCv/Ps6E2uiRcmrz4g5AvARQuiUE8zC71OXTORJM3R+cRov9
5TUzsREnSocVwVjsrLIGJSy8M/NEqmhd2PXwcLV2RNeCB2/nsT+TQF1qL+S4aCA3vKUOdzq/At/5
qIMjDKVjF4JEOoRbG39QpYVdbptkq67LUaIhunts36pWijh3dN0BzV2QWkcXasImymFp/50duM4q
nQuJ4ux5CfJwF1rI7pX1MO9md2Bl5blwI3wkvea/jAPkyDklwyGvJOS6JD1jA4f6s2s/bgt+4hp9
DLrCNmJ3cbJlvUzV2P/mSYo683dTrKZ5tUbgsuWNgIeVQGXJSW02BWxgXv75o1pj8+VaVYQDyJ2H
0cPE2JDcfTGgwTkCVxoA7p9w30GSEAoGH3z87e20QymdyprEf7VjZxpSzcJlF/6FNdCTBj5/M2eK
yi7obwpmcwgNj9sf0cb2HR3A8hg9ZzaaWVWtNf6UmgoPKsZRy7uG66m7WyWTXreCLspIVF14sSnw
RJm0W1bh4Ibr71XP/4Qj53bbPgFY2YxPwYmtwSyCVyVJ+Z44RRLKajwlg+lNJ35997jTwZkv3X2p
125bIyg9ljxMfuSVQ/gxVFNCVgKMwvo7PSGXMOhgIlyG6OdSojvpHIp511cTNhRWHh5djCSHBqpE
3yn8CjtcbjgNzsXbRGZZ6L/a2xxupQISXzjkbw81nF1SmfAhnbtKKdMtN6/8mBrQMmG115nGFlnA
AJp5UIJNiNep47V1HGY19JqvJZwcMk5KSXKAF4GZJ4kIj7c4wFL9uPU5XWshInowvI8l5Pf4IZTW
zSVIxR4DhRMdsoJeGI4+2+YGak7CRK2R7MXh45Qio4gUv4IAvbDpuaehiCOHqLFdUpHwnFiSwh2l
jVq47m/loNiLio3FckTuSZP4vlrPdG6zetthcj/N9uujsPnpF1EKZXGq1k5q1LOFl9tzjUrJY7sD
qEXYk2ccnbEMfmG2QtlZzJjkMxWw723mnxuicTp9PYDp8c/VTODrcWNAAQH3Yua81WVrrcn+vOe7
vULVF0tBAiB/aTI1fDj3fQcBmUYVyPf9jw6LJhGe+uoySsn76jA/ilgdvAzTfvmHx8xgAejXRrzC
MnA0yaqLWSUTANCmK8AsU21wJITx4M1CybWaCAAc/du8dRPR6xiPvCp2cx4txpz3URjkb4EEbqg4
mYYtky6ief7celpkMvEgQDHunlanOAj8xPuQDDV0IuHKIa/UeLG2xk4iRDPE4ejvb7tLE5Eirci+
k06fgt5CyZH/kMXxI0QqFLae40um0HFytFFayC/W/RFA6B9X0GvcfRHPufIfEqw8KynSCWGBMc87
0DBa8gxLEPDtXaxAdWXDi8zsSkBDc/cnGvRvzy6O/2VecioxxWnlULzPF6g4xtPkyXAXkxVwpn6N
AwdH095+dS4CVZHDzqgxZFLYBw93OJRYEe7N3CLoR3WHeth/cmvWo+0s0PDyZRjT8M8hU1LsdTo6
8xh4r+o3ScVMm1zry/a/8MxcAIXq4ROUcyGZtv0PAMymr69H15S9WpKHNAnNgphlQrj/QZiaJbOf
VKcHoks1SfNgCq9Z1pViStSai/mEXBzCsyqdkQPyRMZyYMmOwypvvWHtLQ5wy5gvDa17+wXCXXUB
96sBpxoVewmxhp0KSbj7opvzcycKWQw84eNc/l+mQxZctD/kDzgrnuLFVe75WOtqIepy9EHpm1FG
BPw3KxY+G31YNpzWUKwvmkBCrejgkUIInvSimqMqCVFFPhigjmnTflaOL6RhuhdFD8UG9Mr93E9D
qeym2JK1ZiLDzLRwx9SgW2m47VOkqAeA6xvLRo6PmFjczZ44tEnys5qltLZx7VPOYgoDIEQa7jL2
rO2io8RHD76ft6gIrReYq9SzcdLWAidCCWrfqBmk59kP2ewLtfl8oqPxlwRzZI3j7CHH+D2kgYYu
MphLlrJ6uk5fFZSFr0zqIuKgFcAKrgeC+DpoMqjb3TMFnUg5IjGjERViat/Ww7VU/ihNUTuMSWza
kwzk5MjeG/1sjMgqh8VkBVbzbvu4Zwv17sHDrZrb3DV1ERicmbatovBrQdTveGCct0UfHgU1XoGZ
TydnWy/y5VjBlEuh9dow9EBjo9S3AG+vLh8vD5euAfIlwKIx5/DV+kzN1WyzKbKeDwtTN4kwm1WI
S33bO4+Kc4RWVhWIxYSR+S7T7RCgvFDq6V6a6nbmiVdybfjjrs47swdcb9mLezPgBZBZ6YSSVk4u
gjzxSN7+nYhehDRJkLn9KsPzZKch39X+Zc42FHU6HnAvquHrWOr1/S2Gu9Z1fgsO787dG9cyH1a4
zEm718fkC0OfMw3nWXMKLZfX2MFVq3/yH6StXKrufd9YnpioPpz7rSrW5B5X4umhtS+5Tz9CgI/f
ELv7YkXfv1ELUkUCE1MCphwJoReYuewK+ItQAL7wrb97y4ZIvp00dGnoFABDfvQM0y4hMw9wRTpv
TwBUvZkHbBtzXL5EDvkADUOJFQgEcKF7cb10WYz5roBPvANW5UxxM8Bk0zAtItp5CtPJurLDQSKr
B4ZZD76gy4wbSPe2g/4n4wGw6Onl0uuNC8SXaV/IVKz9N6D8mgaHfHw2kTjGmZLzVoju9d4T0mCc
ABRq/063At7TpsIfd+zTcLGWpOT2bUTF2u2QCaBbhtW83FO3bPn0rnxb+hW5eYDfPo7DM2H4pqR8
9P7fWUUfzImrXkmF+FhU5lh1DIsLnHbAETiMa3YyIAPBTybEjS+EfbS5bq3Sv9ZTKMGFjXlMm1N3
iCMoixD8fkngnTZw23SY8kIEY9dRlhEoJra0ux2xm0rnIn/qebxMwOX1oA9BQbLKrto22Rb32UtM
MOL2eVndsYYqQmwh48I6efsRJjPXHzGQbNdgfJIn+dCSADgI+fKADOZa08bzWs3Chv/yt7S8Zuo9
xrmRsFoLPEZ8rktDa19yFDGxV79M2sSF381uvusBbUMc80on5lVZqmXUOBqQy6uRSgiAjImdi7D2
FsP8YPyVZIAqKzjO8e9YYUMX2bi38tQCaR6k5mrCW9TDJG03mIB9ODjqi8M6TGe4InVI5uT6NIm5
h8jc99LgKyvO9mBPjrvNAwmzjBXGSoosVySSvrLUBi1j+Ca3GDrMqtWcW/P04Wt8YQy7HJ9VwNl1
9kWGYGYZhhDqMPMjFHvaazmWZ526KlXOJR6gEhpe2WZPxUUV0B9WL7ttoKtvkORUfn/B0m6aVkvb
OK0N+B73y2VyXuKer6aKGPjhXqfvl7y5EXP/YJnBeOWJXHTIOgbk4q7m0BvAwSkmB/4/lCFDW76X
MCoJQSFA6XcEftHbPFlNgevO4qKeBJfG60w8YJPo6uSVTFTOoxQ5AzZ4E9UTfU6ARNhAt2LgK2li
JYofVbA0qh77QzWipVpMhcpf21ZzT+mzQfoPKNL/73KCNtsNeVNGSBz/PrbwXQ2f7vjI7xOHI0v8
2Zr6Ec/SLa6hozkspUB2a9Ao05YmehTzgEJ4YKxtrGJ8lpRTYE60erZwC33JbzLcBLxh+4JYjMrT
useLLOqS175x19Okv399mmZajPfgc8AVA/a/fUB+mbjFQA1I3ZT1pgywY0fPMTrwcyuz9YJSX8Yz
i4SUJO33md0jeWBp/z0mQSlIqC87RPD8MOAYLm2/xJM9NiZEMomj5Xbb86R04eI3qIYqPp90xSWS
tDLv9ncoVQQUGMCfOxNaZAGjT/hDoDlFWDnXXHPK4q+UBJpOWFN/G8eigYvRR88HZA+TaNzqC++5
X5umo35eI+TdCNSPASrptxsTl0olRiK5MDKU01Oed4YN8F7BIpG17f7nHdGurx1EyMZ7c2w44C5P
UOjhlPWnfKQhqrfg9RT/UUF94QTZBn5WNfw2mtZFk6vIlQnzZsbAR9TjeuBd69Xsix2bnnV+wahD
n+hKImB7sW5JtkZ0j52PC5HF7+uPejNmJs3HY0gjXtZhiy37XjXSbKt9ULIIfrResuJCMQJqlDoD
E3o+9X/vgPE45Jxr7dxcdYqo7DS1cJEDnJeISsGVICh8rlTVIE5Uf1tsDc2vBwLrd/7hLsGHoZzl
r7WB3b76OioraXAbvOPmz5QU/UvF3KiGoGV4f5w1J4DfVnYcKAI48v/2LBYpjRJsljmeDaZ9JcFA
duVymeTqlGsHUi8yHNV3j3VMA0KYBYH8PwIib0ip9w6Ho45iQuWfwC6Kk+FQRjulkYJfD7vrrq/7
+N22/O67xyGAwHTUCwYK6PBENVUnajxFhxj5tEpcp8aV6iMknzsntYZqB6b7w+8Z4fcYZr6xDMBD
MbEBcx697gPm3aJDJYhJBTxeXZb79Sx+US1opLtm/S66m6nlRclet3dQfKSoqumO9NHcQz503a5D
LAQ0JdDnLG4mFQR1PqwRjppHXRRT7FgNsM1WWLT9SrP7krW4LU0VbJYmJ46ubqjmpI29R1EZuj2E
InL0xUz71w8W7iY4Yx2QEZHlr1BAvG+AbNaD22dzmopdwZ1CftHiOcLc+KDJBXLl3SbiXqGfXP39
tn1WWT44qHG1J26MxGsK/JaGaR1FnlNcXGJaghADtaOqTq/7Ty0telR3P1tr8lK5fF9C+V78yk16
SB9er06CTRmf53pZ9mkmtHjUyn39GUQUzOAOudCfkaGevbRC7O46cHsuHagHAIx5w5P5frK1//Jj
qjFMWH8IYovx99F85qN+rqa1hWFZ6kHM9J3zqH+LCmHwxw6azMwMOoJnC2Qyiyj1CNftYREYuw+V
XdeW0ISJsJRanO/hv+O8gLYNNN15xvtXhEUkRz1i7vetpJSlV//8g4THCBNCq5SsUjIiosgpjgqM
8xIaxkSUOWB+zDOuPQWrGdSL5kOazUesrGI5us5YWYm3Lfgm3RBglfbRf2OxPbMQyA+pN+6WiWKY
NTd9acgo2Z+LIIfdEgoESgGD0z6Jawsx6NFFmgYZ3zYpyqBfGm0ggbnKKmgo/+qrpOu+NzT4835A
N2f3uE0DKsmDPrpTDtrys37J43KJlGpC6vml5Kx3OaoLdzqK87oxbzcztYoZ35XRK0MarpO/XA6K
7+BAjz5mbihZPxEUn8fvQ63jDPMQBxmMw2EPhf1i0YMhsZU+OkaP/fyZ7zKNsn5rl0y6/HWQbVZe
wR0sETKedngsMu1pedHpsLAqQZ9e17bz9vlB5jLWcC3jLvuJXbVj/UtWrYYAxoS90GABWz43dq3a
oKEif2TC1y4Mt4s4iI+38pQYS7y91T3q6eFHnaSn8P2lFltcxYcldyKGWQpPAEhs4huEWK0qD1j/
L5kONT/WJJjY37qvEIy5L+xcyuCGeqdx8ck8hPCPxmyenuuVb+UNYxSy6rAGDu/s3n4WNWxEmNAg
/HNu+5boaHbMAcb6MoHOf7s/H91VyAB3nQa67k0Eona1JLvBAFWxCxQVvVXHaEQ5/kdhQppm7ys4
cijSoJLysOsCKBQkn8WLCr3695NGJXj35tMjF2xnmbLbW15oOL/CNhLG6eoJchXo98+kEjF5RlWd
fffzWjeocTl7g9LDMREoGV15g0E8r8Twgx6p06RMaCcvMDMNKOLoP69c1CeqBhHDm7mTS360b5D5
NhCF8VAIgSKwV2Qn4wBZNarVvufEiEvZfmRFjY+aeSXIN9RPlVJT/VYmQlenuzxw3aomFrMxRblF
5wzGwmZiYxrnLybJOClFlJUw1QUMDd+3iwSA2fCGYiT/gYqkXQ7YpQgVC+SPO8Q8iL8M+CHRFZaN
65GNHQD2RzVf+8qZ1598NweeO+2w20rjudI6JLVyIiD+GsBaR6RuKir9/09wEZkJDvkdQtukb0/j
/yyumygHiFkoVC60CQpEqFY3E5xC/w2uWgEO6cUM1I1pVrzXdu7g3Nc3O2LLlIkuMwgIuLXy7Qt7
/sFzXRtSC7eCCv0KOWLuz1SVfpQUnVncC6cy0bQIOARe9unv3R8Qmw/N1PEp8a42ipORaqAiVPhJ
jT2A2gsxf2X27oAsarA6x7QTfF+D04weKoyquNvmIhfQrV+3eI2nmmPyKobEUgBhFyzkG7iLpv+J
DP4kfnHwBY1e61uqI7aHFP2or950cl2P9329FigwWXKkO4wjI1rDbFDP+xpzneRs8IpTVAzPZ0xP
OuSS6is4vjcIZ58ewdUo7wI0lyekgMpOUlSQpsEhXFwR15qE14pm3Cq7rcjl3NufIC7WJ3bHSwZM
SBxac2jipbCDbTiffbw67/N10lPxC+IXXQczk/aCI33scMH8r8PGgylct7vAd62fhcKnQKIXNgmK
2AuLkTfGYqzjq9B3GRSp88zkb5BXwUxdtbyWfRsXbEM5/Qo1wo6hxOA2UhjXDUwwLQeIH330vX+H
rcU3KIPtbH6hEdaJTUs89rjTbkUZYJjCNK4O3BCsqqY9pJRwe7ZOniJsTeVGndaxAvhVe2a7GbCR
iy1dW3U6V4LUNQNsbDTR1YL7eofMkvT/gLfngV6uW36UNRIFFtRXaSqkZgA5CRFL14Iw0Jlm4qpQ
Vmjl/Ci8caluGPSpBLAGYDbFeHrwcllhfFmZvMj1kq+zUpjGBD4HJ7KWnWzIQpQ5chjLXCZpAYpy
btM6R7Q7ettI+zM5q7GFbWuMOTHxTa0SMGdkp9GxlivkvHpQkOFMlslwjb+kiZlF1bRsmPpfZ7v4
r66wzzvEMhyFJyi2lSIeJfNYRNPOodJAZTBVSOULNl/0hQMYfemYTKGw7cBqJarXdI/SYDlM+puW
y2HZ3xlNxvj7as7N1Hyxx/N1o1aHh5QEWK8ePxjwZEMHh1OQBJAcyVqkbX/x7b3Q7v1+3UYFuBmR
e19KIizRL3OOa1Z1a4oGaQsq+lkqY5HoOxiSsZ2CpJiuMyBepOA+xFX5SVUuWzXvGwBPGVQHaNJP
fe1Qcdn4HzL937OPd3fSMFSE2njYZ11KLo9dgXh5aVj4+GbAgJAD9EBOzkm8ffaDXHYZc21xUqRb
MkpGTJWj6KzqNTIZ9m5cceKWfP/4vZgr/jNQxZjyXPtWHDZXBPybPM1hxQ/q82vd/mbdcg902vSw
efMQzxZ28RvOCv423qI9p6XNbgoTZ8skaFHaM6pa7KeGqRpf8tOm4TrOqCSDYDIFYF5xoXGNKlQx
+T7vE5gZ5Tb8O8xoHCjR/au47A4NxW1ZiLyZqdvxzjnJM4fk7LkPgFsvjmy1LS+LvwZwyPefu1jN
HaI9ofJQsDZ6ipxyRjade7mFcJn+NnM/43HcASiDCFM+220iczqOFXNxs5iHMH143qlTpUHqcKyq
2ZQVtCY36ym51h2j/M1UwuVR/5jyiKmIExwAc48i2dlTRzRODkvU33ytehoJbHs6PnCPOuT8jXFc
hJoJPSsC6qypScGFSMZveYuiQ+DTh5Qzv3A5WL6UxgbD4w0HS/91JZoeTK1KWAm/ixw3402gn3tL
8RU879N9NSf2B4Os8JDp1e8QSTIOHU6JeeAfbOgLX7dULskYg++I2ygsy6eqZuiM81odBn6z3uBM
tbyllZgvs3rkho/rrIbdcbPWHpKt3aEyYrXONDx5PVu/Qs14kwfsMTthtnGVknAEVtpr3CTdmD/u
LMe/p8km5PtMi9Ig0WqYxB82uWl1diGhQcqAqVJvv4nT2XO01M8FrjPc81XC4CMnIU2Q2vKbxKln
m5lYqf3CVFo286SIPaPcBzSZ3VQVtWO2QoSWiZ130rP7fuZeA3jOROYiOc3aV0N+nvQAAf1i5o98
eVW7+VWcfp1lHlLqNZsMu/8DDcDowdp8HccMgwbo1ypo+peSIPICFf7TrafEL5EV02GAt1D8oZbP
lYwMlcJZsR5WeXaMJFGDLOXAsw/JKYJ6FY8DGCiE8KvKbMmbFL+R10hl6C01kaHcSh1Aj18nSzcX
jU/XrOQmXWxHoguHqmqesJEvTYCiGivX9P3ToDDp2VjogWArwlzlpiSlTmV7JgMMrPBC87sGdxDB
nKbTi1TqBTlHPdtHK6CEgpjQNFrtToDcuZIZdp83umOvV0Q1F6hQLI0Z27dETm9m4XcvpQ3ACjJG
OsTrmj/2tx3FOFZQFtArMZ325/dY+V6PH4ov4ds7xjhgvpu8U4FDoQRdx5hYmMtZjZ90NOOY5kpP
i4lf/LUd3MbN4OJfPfDep34ZjKU39DKJ1yLvzA9BgFOfxiEdFGvh2HpFyv3hPFRLEqRornsP1LJy
jgSslzCPbSECClu6olxjFhUr9XHbPZ1cCCpiuHrulX5MQ+fjGslLqtUCwvtR7AyW7POeXjQt5DWP
OyChMilpid9/RkJog0F73G0St4dc0RUr2ZkZUcA+sFIHAcliMTDBQ437FdKA6LKD4SsZE473CyP6
RJd6rShGw8lzqZ/cqXPOlBr8TAfzEgvFRubYRlkciVkUvQ1sckzEXXDnghO1OBLDP3V0Q6g8Valw
mMB5Qkkv63Rs0BKpa/k+GhAP1YjJu7JO0MtVCigkZwy6M/n/vXaZyUv+Gs9/vN+9/1I6PL0ao1ud
0/k9AdJB6zgtVm8TkDp2CmeGNLVnWybtpPnp3Ln/tdfxiFESeoaX54IoZFpVKGKstS9+RPWrbaPN
o+L3ZhULqPsXQXLuoWP3SqaZE4IGzSByieSIl3h6lXuz6d9KEf7dfMJHI7mpRKwggNivLUNB+jps
VcU/W+3p+LAQSFnVhdFpZ62VhK4P9Mz8FGlp0EKTTyuLuGLMEc/Qdl5z5sm1KMVovXPkiorjm+wl
YLWwGg1tRYbWQh7AoPyTY0Bsl/fR0hcnPCcdXVbJ55j4Gsa+yZbLYYUIvdm63Z6yBo5Uimh9OiT2
uWwnNbNW5eiwteA79BQIKriF+/2gosS12aNNGGu9ponYNmzM1QJQyS5Y0cLTcqfYJWZBBlKRL4Ww
2FO8nLT957fzedGJq0EfU0SFv1dc7HYHBLQ+Poy2KRde/57k513fLEB/2gvEt+sIhUXEEMoCojoW
Q43pm+M3ekaExBr+OIgL4SVN+MK2uBb0xlaAS70iZhMyVG0xT856Pt7EFRkZl8yAEbABJSGh2tt/
NcusFuWhq/zzZe5MqRFjmntUuadJTQAgfpePIJPqbDSCzfZyrhTkpOHqvad4v3UnF+4nLj2t7Bo/
uAb51kqXrKeB+PJFsg+3xxnxwOj6Ahk4XDYYJuCc1kn00XYQD6HsFymAEstUYLAOLKoxItoFkfS/
Jch4+9HSczuYJlRG/pDg8uHXm3GOggsIhzkh+Y9QRkCAvnQsXRS+irOWvBvoz2zp562vHdlqrHX2
nkdAqFUjv9/Kc/x8E4e4RagNzviLPJdQxvA+Mg/e2COpJoh6jAevPLHjSKmBsHhgZmgYx8csrHCe
lSGdY6TO6AJnKuWWhQ+BWiycJBcSXPKYoa+7dieV1tiohKGuJLRpxF1EmR5dlNjLbmx1LH/qJTS/
OAABpDBE5sfSbCsbmP3V/GHLuSmUmVRvJ/vMehi4v6irj3AM54kbWq/9/lZf2oQbVkh051HkL3Lz
yuwDsB2hQhmwSj15v4YUWpNK/F2SemVOdI/drNVp/eT5ynYUTXB0si1p6XgOZYa/+NP5EBNESGAp
hHyNCt/n+vYwtAwdO8kQzMyUe5x5Csc9q4asnjZV9ac166sjwps/WdIBqHtopuXSnO83Q6iCRmQE
KAASo5rbjbSHzT3JPo8gbrgYk508J37+p0DWRRStOYpaZBc5hkzRmKlw0M817UcJ0OzukQZG3FmW
QXIkZTNf8bjNng4FyXljUnw6/QZkRto0Pp6DY6qTmVAPfA/mwtqgAyfMbLtEAUoD4rwSfY72IHPs
SP8NEpLJTa9N/Sqa4q1EcdWbWDBSwHvYtjibtxWCIGP/7n5ltiextd6qmYdRhvAEgglzsA6d1Vtd
EA1ua8jUERluKhSDLzmeIVEhMHK/H3u9aSCVWgdjG28eVlvWCIrWm/0dHgEZP7mP14qYSbp1rNJp
USUD5KpsSI7Vyj5d5ah+hd9v7l51b89nu3ziaK/zmSu2nwu2Dv790KU4pQw5tAFoGsMIFYYGJmqv
6jqcfO004oOTTOp38S07ZVeBufCoLWNwx8K6IyIA8qp1d544hnXHrc67//2k4iAHxYMkB4YeGKDn
2mrX6/bQcRl88R7uNQljOAIDgXfWSY5LFPPeVN1VKUwOmre5TXgRJi1G+wkXoW5Z1BnQigYqQ1q2
n/CgTMYhpKoe/sh6R+GLruvUiQWN/sp3Uo/bBM9wSTkpJVExLeCbElyVXj3Jcu8tOhRYYqLg1GNI
wrZ4nEFhtYOQFW7nOjOtmv1fz+O9vmH8IbXA9vPoimW7dY2zyoQXpzF8A2QNtgWRTq3HRAtK5RXK
U4OMKW8WSsiLfMAjHjtZIEY1iiix14JQdVDjUg/2HNvw53OFLKVJXkYBU7bjWDTF2ZxXXNI1dVpy
zr6yBJwSlc88HyYCwpOUBo9bnM8Gbor3iMuSBShq9Cfcsz7wt3wExvB9dcns4swdQTatH39384yL
K375mTvpLauWZakAQ/1hpvnEci1dILqpjzhvaFnA2cTfbb32OM54Kx3U22ChxnRa8uouMsu67e8T
HWB57rWsVyS4Vv7c0wp2KEOPr2ME035f2giQbMTldCcp2LPFUsWs/XSAgi3zvL+xwXuuBK34mIoP
ZNjlARFn3u8XPzMkBxGa2TJ1SDs5oVge6JqfwdAYGAKBgiZQLYJoBxbGAs0OBvM76/VnfBJOsshd
Y+A224qx1ZnCVT8GqWgF+2TZZqpqj7aeY+7vYdR10frWAqnyi8qPX4bqlbedH2ZBXbAZBPzv8Kpr
f2Ki/CTFPYQx3IrURNbniHxu8J6F4rKgOvQ9RXdTZgnLRERY0mD10BRCu2wbKD3+bSsWvvhnwjs+
vuqJUISIV5DbnlLw4Xu+yMRP/YEMPE0yu0eFBklVCX+ZCLYfuadeBXLxizfThIHMGoFiwiyWAf1k
rUcIR3vAg2dstPGXuTKPEWrT6q37a1JcoUxbRxf89X95xI/4qnlXM08OLorzUKYah7nabUCipv6q
e7bHGLfpCe/ELBJaIYET1tbqBttdk+h2/N+JDum7XZzPm8M3fkL4AosxxW/SWRaCYir5uBqdSVGE
fQEfYgOwxh/oOjFtP06xJcy+ockEbNXSl4qfda8w+Lrardzq2j37r3C+ChUT7almymQLk2sJaFVD
FWOYZb0rkliS5czzAY+rGu1UxnkLp3skstsHF2xENTsP9yasYp+tloCHEKNUZ34C4PxnCaQIL73n
177oFHVIWBaz+TO6tOjqpuq7IPBK/deN4WlCMIrb+nmPVKrjeuKbkfe3QSXCMLakpD78w9To42Fl
83E0rygXWIDBriuqkoySfOUqzc2tp8Z5yLhbhhYMXXPQodK464h6BxjjCAbwPEjOTozcmDlMXrJV
nlxymMe9UPlX85Fz4A5OUnx0dUZIhn7yRIMVT77Ve3mVygvkgirYhEWyd0lnF5PbOfRc1Bo/0+mp
F55pfFJVdUN0e03Ipd7nkBC04BDWKexRJrzDoDuMFYzIjQIbT1OzTuscdecnq655+4q5LolWl73C
lt8D4Jv+FxcdAbz7clOYFfBT7adFeGu8CKeAolJFrrbzWQ4gFp1OzldLbr5n8A6aca9x1giuUX+E
VKriKEyyl2tKCZUPNu3mrhaS0v+lB3SER7n1wu+hqrQ3MQMoQVdxwpRX8nW1g1zk4UsAKbC4xzV5
+wpcXcdtr07XoGpM/NFcuy06rnQfg0HceJzsu/Un6yeyZdisHgBp3u1TTpS7SAOC+mgkFWVwohqg
a8d7A7Q6vd4dJfyfEXIzrS2xPZauySXBiMrjXn8NdfpKFKElAUhShRumT69AdG/RncRibjsdC700
8qOhsqxs4mn0MkXijm+2ymRx3+mBsXlrfa8e4FNJaHdaf5pnFLDikGOi7JEb9YqGlQaeMFcneotg
+H8IX+ctNm9k+DPeBHYNqR5J9of9spRECbvuGFbkMK9H/2mfGRrM+lMtUyAh772DzgNjmk/1Ol0b
gOQ8SymCV9s/c4QFxz2l8vJD8Z0e20ND+MscoHJQIrvSIBINHxT4CW5wJHhElZmj8VPkM7kD+wTh
qEy8xOBmMnTL8T/ZdbNsI1gEddh/Z9A6ZY96mHGB4rpKNxsIUV/uAPjMNKb7fJZkmzxAGcXDycJg
08mjsmcykGJfglDSHKJHXcTt5dD6t+XV0mb0FEsR4ToiKg9KDAWW/P9wrGI31/NyKaU3QEjFfrhL
0xhrTKD1vq2cCtwXXS0zhh8LNU7Q+PSDnqjRZjXwWig2eqE5N8yw6a9nWQzQm1u4o8hJrK6+ohXT
UtioBRV9rbO5mqI/j0x0kE3w/BVAsVJFVI9Ep4XjxGvJaG6cd96RujmVE+fUKVhIknmaGc3O+0UH
M1K/SzUlzSVlTvGHKDTy7IA8itPBepbSOFaXRw52EKEaOCPdz9bSN4UXYuriNA1srWgertOzzmxk
zAg4OSPwMTT1uBlZwPFT1aBk8Lv8HCZinnqalNXzKKHecQ/DmB3EBwpg57EaSBpth6WN2aORoiek
6k0idYI9Xv0DEjaRizDn/+VlIt2WsInVhpMGJkvl80Q4xVYvgUGqhrXevs2netPtcAMyzrDaSjSK
UaDe3RdugsgFB1dnpxNeeCFY256hP2Zl6Da9qYWy/E847ln0m/yRbvclD8UoCRIo18KY3rNRa6tx
o0f3qOyqswb7Sf+qTCw0BDDg/C9TCyIYpPOZnckEd83DeX9wcpD8lqD4jaMuUzrPFtNtdyHKj3sq
Pw6/gMl+u6snGF7Rolp4Zz3qiC5LblR6WaJvKEvNrlYSGVmFdgVr+htMCD96lUad8grENY8l91MI
xBhHOp2Ld+Qn8rqt69X/cRVizwKZlN6IUpwSSE3VjsIYE0CPk6oxz22GHFm5J2ppxQC2ucUX+e4y
CxHbc4Uc2acz0SaUQ7tNQ6/eB4j+GdjrpCIH85P9SrMpWEsvtex4eLCGs8EULXHl5wngps8vg0NY
+6K72+eEKfi5XTZLuFrk/quqzkTcAD5+NkaP0ZWFMWH20oCbCLs6WDcMrRGegdTl93L8PJAKnJh8
v5l6f2kHGqogARiUEGQ/wiB8Ta1uI9SimjE9lVpk9U7QRPYO6FqggSu8bDUpnR/A73YhsPo3gy+4
q33w77qgONmrksFI0MTP27psLR7R+QtOoVMqx2CoSLreM7LC8OMY/n6yy33anj0pBBUVk7JZOASD
T8nNj3BSN8sEyiV92dTbJXCmucO59FVDoT6UpafXw/5nMy0OCbMLhyMTTf7n7c1Fig9QrIu9IXSV
/kFvfNCAHEFyvsU4She0sMmXOAKmNCFQtQnZ5B8zvQGBMipLD7LUEq/CEXK0VDWwLDAlVd6s4uOU
LheepQFEXVlgzYea1j7V4Lazzpk8o8k1JwWBAi5DNWCxDbGLOuYpkfgSULkDbaI5SzSH0xJGQHW0
mtVhyKrSYzyVmxdKmvflmLMQ2UeuQOKw5ISmL2wMOX8lWTMU8eQI5+wWA7ZSPUD5nOUKJfxYjUfZ
CJWCXzrWDjT2dqFa4OrDo70D4UjGIb9gDwLfvWJN6yaRqVgL4ga4DJK6x5ANUeLA8LtG658UePM4
1c/tHdxTnFeSHkBMrxXN0dZHIWjMUsiSFrOT4fb6yatope7/rwmzzx56NVVidINQZOACsE2P39ss
hTvpWZXlxIZ5MskZtClciUHurR2YkoBeoZQvFbjLhRYvSuoV4zts+m7h0liWO5n80mdhwfbG1FJe
FB60WucRGmC9WfHl8Ui8d8L9la2ZMrn4uYDPGeocRvpb7eYFE04rRZPw1omxJhbNZ29DzvCn/7pl
Un3oFlzW7e4lJGalddGAQy3FfbYGVKn4zm6F6/cB5rf5cRgPdhUCJxyoRIc4S29TBZmpJfMWnE89
Lv54e2vxxw5k6lpkn0BQcXDrPa0jlGkUWccPPiIwMDhduVu96hodmtq5oHNBSib9TTaW1FwhhsOw
tX1AH/ErGlf+yVeFuiB8j1sYPyg+gQYjZQLPYgzifrTxpR/QKfRPpLApMUJ/mVYbE9XIj0Ld8cS1
gk7l5GunJvlC2+s7k7BP94TvaR0ADOvjfWLiXG9AXjkZxL4+pic35O8JuH2ti6SgLy7QNGmGh0+x
/4w7mSbzlH6TFMPA47MKx9dTBf67GRYfvs+tWQ6CdzNnwxVJ4/IPr1sW9K9swsG3riencCFW8f3i
j4jT3ra42uMvBIgVH6Oqmg5R18Y89+SDRVP9LMWgdh6WsUmlCBjzPn4Um/neofV/zmVvmhdKPacu
QSZVkA41D0CS6Af6/pUTg4pu0Pjl8xoB7rVad7Q/KScs+03tcsU5bWoLAioGB1zqHSNV4Ae/ZSaJ
yrEcqfkQ9cRifq1xoxuCpmGaSxnTfhQ8o4hb9cGnZZ//balEPgF/4I+ME8HYdaLGYzgbdYKwmvQm
fxkiJS3GQLN/a3wFvg9+DAV59yXV54a/1hRNEX04kM8tmExZhXEhlZ7xVebZExPv4taS72kJOFtU
k4yEkSj3+Dl2P6ySk59Rlvg99LyYX3440lffHoOWIGFnBjBtDMW18KEH32M/Shg+LQOTXUUREebr
KqYJWgTBClqTCdqoDMtlO63DmMnKMg5MisjdblcRZChft0vrUrFhPYwy/dGsBIRZlWCxVkbUzcVF
KWsJnD63/Zm8DTDlMREYo063DVGwFnARpQ2OdA1DBWmgzIw/ixD+LNYcPh+sYeiIE35gHu0yqA5u
7EAYB6bSTl7dbWvHXwxK6xys5h5xGGwaj/H+cH7dsjAUW19AHntzfzYcHivSi7NbXnvZN/wG2tCN
IJ5SSv1qykWNCnEke2fAyItxTGkCmOL1zNd96JG4Q42tohPzCwKSxSE/HPLL2YJUAlDfOFyxrd6b
ALgXSyBtwaEb+AZFr+Nz2q2SCFDjeeIm2VTi4Rz/ZL8TIb5y4HmcElaejpb+KtUioti6N5KBpw8U
kZQD8K/MFnXOqOz+yROUBwhwhtD54lMUrkuvTRc3qVPMZTrTFY1pMxDz2nc7kj9UwuUn/rx7Hcxt
cJbtPls+nVPLQyxQguhRnGd4PnCAsC+46F/Rl27aJ0Au9FUuU3D8SOeex4EsfQHsO9PfYPe8Lgpn
DgXZiNcbo1QZwsnTfYmHGJq8AWtT9zdQ3uTxWnWZB5C22tzxH6JmOJAsDGwoUYFiPH604B3BLXXW
7rNL5K1/kFud3+8QRPCyDvz9z4qU+Oh00AAQZItyKKL6JmiAMS0bLCIj1a4qm2X2NWK4mlEMaozo
cmSVpLsrJwRDrNEpSm/5XI16dfAXFoxOw5SvXnGWKRqqgn5pHH4r7rtm0Yy0ETgquVTO+erEcYzC
m4DAiAysvSqS7swRQdWTK5NfZgxzfkPdX5J3Ci8gvK5wiMRBwq2lEYV0u9Qjyn9jX9DhDlxRm0Ip
cvpCaUq+NfI620UfYo3qQ3w16c3IR8ZwZmCHJGch5y/pfOAzVHXW7M0CfxzyAiHNzaM1AqiWIfzK
RDcM+su4oxllYmnSNQqF484jINYeYs2St1q4SDCcR8H2mUuf1/ybTJk2QLkVEVR5Y+IVqvMfg7BL
VCjpU3heNbnXDF4lZ9z3KDUbuZHcxve8hUEq1bZ369gm59VcDRlgJogQae8l2XjheKmYtoCgvjKi
7ThLoCqJUF+v8ANgkMAnyOvtBvNboDrXWOuRjBIw/ha2ekH8HPcLyD/PkkBR0KWEzlIM474E+AN3
gTPQ6HVHPw0rLBAjVV72IDbmxR4+PHUc9Gdpt3oJKw0bFY4EyVLhAZ+zAMccHcCw5anbl3SuKujl
GSvfffQY5/q/fWWZbq2XPgkhnulYIaeY/67U1aXPTRJHDg06xfh6LbSf/8YssyUneP+xrdPSHufp
bt8Y5y2gn9W3fdLYPZ6zhsQ+MFHIkz4GrJjvZIzGoy25FIRKBombDmBNE953FmGMC0VQbP7+3Idx
NGoTsBDvm5mbc/bn2egjU14ORPuJAVzwGK18dEMrwyu/okkzJ9WRQ1BkXDVlZhLxfrgZQ9fgQLYP
NOg9ewj2yqsuAWzWC5Pe0AOisElSqPaJ3gXpiLn8COJ0mjLbMsf2N9eWNKQbF9zgObeO1Wuowfio
9ikwocoQQZ0MJZ/9kagm00gCE99jdJlfWQmFu9kIe6jCOMEgXEFWACZgWShweZNJeQEFL99jrU0v
ZSPk7OAzn2MG+suDymQCi/n9Lv7p6SYus039OMwl9wQrAg04gVYqLLA/Cqz6iV1f691hqGCShlR3
FYAbv19ieobtCmIGi0Rz6zxQ4k+kJ5NXYs880zAzik0JoxJ1TudeYrvAvvHminYw+wMF7n4ABxas
PA9/UBm5hYPQH0ZReb70JA4Wcq7lHjr5CPMDlUWCfg/Uwj6QLEiGUxddWDb847e6FNVs2aFqW/Nf
I+mFiewWodIm+3dxq/DJvHbSStCLLB2s09lTqT8nYsa8tpIb2B6sLN7pB/1d2SvhogXF3RQ2YtG4
mMLUFvkOaBEXDN3ANWgrbrTqdPLUjbrJkDPF/Z5iXkN4mCx9FfAWshGymltzEsFqiTz+2y1ywKsP
xEIQ6Vc8wR0IOEfec7QQpltofsC1cGmTeLXaXA46ef4aBQxkYfTkzVPFAxXSVHOFbXCHp3NhxRjp
i3G0PQWy1naRNq53DkzUSUQZuRyx1fgHan4+urw/jc3MnMS+kFSBZeQK9lwiIbasJpAtpKjD51q5
t6YnZWTdvePTwx0PdoLtUcUsUDn6Iz+d/2dSSHYHFoWboOpgSKNNSHpjAMRc/7VaD3UnBtNTTKMU
hzGiqc+6jlQN3ZH8ru3au8tN1Y6qcT7fY6VFVC73FUs+mhQv1FN2upY5/nZdiZDt27E3M/5pNvca
aZ0tEze3tbKERroBDF1tqYIzzmrWgK/ea/YZXzuGy3j44M3m1Cc1cuOaxsyN9l5PL23+gQiYCfxz
L64EVCmSQhFkTHyhkyprmklwiRK+dwhdaFzPqXeV4566AEVIJGAW8rBY0K2VHpkP4gXlElmSDpO8
vsP36M6QP1c240EH9/I2y8vWnklmtgNLMLtFZiuQBSVS6sklnojx2LXrC9BVeZlyDGDeBv8kpUdR
FmhN0F+ZboZK3yQE0eCXcfhRdCZhr9Jt8fsP/LDi/HTBuBs6FP3UqH6kwH1ZWmVFIf1rX9UPEh/M
/eqYcA0wCSYfIIqCQELjMo79ojd+Bopc1drNhekLHClRdE8OO2trxEXJiV2Kwcz02RWAhj5rZ57D
qV6oR5Jkh5tz2QhlFIPVBo/NhPgnbojPlQufJKZKrl5DJq6jJfdZxEmMktJhJceBaPXtBCyLXHne
CxpCmjT19+2lAxioA4OmL8/DwGP+naVU9P9x50Hni59AeEXA7cprvgxO4SHwb4WW0xeIj7MPANVq
cHSPWifHGauj8M/HaMmn+fb+BGohaTo9yjKCShqxX3PS2RpTjMK8zOLmhBUnr+8eUkGXjPqFpbtJ
LIJyrFhmRJhjXdYvXj57R2hknaJuFTyCQeodhF2twNT5xvO5H9/MnxJH9tsxvPmc/iAKDneSk9DX
1XUDNtXC58Cg0AtzzXYm653mtselquuUetA67csiuUg0rI1ld/16NKiYslxOVXySPEVcI4oiSFpb
EV8KiHgDz7I9MSn2afTkfQbxvEZ53q/E2gEitnWZq8/iyicOKgEQkCGEn6ouNhUCmNjDCGU2VPyF
PiY+HkIutNsB1QdV/YORm1lsWrvM8giVtzfsYBWSgmVshR2PK/vYvwBK4NAnLI4UVYwwgFc+vvkX
2XAQnRK48N9vfwZ2dWrzgTexHDHJm2YYvgjrUam5zpqw/8AzoBXHJXwcz9gVeWNZ2+iaue9l7A5k
4ciL+YP+udSvWrPupTGAH47OddDMfyV5J3BatEhYUlkVFdAjRuD7ajvu4LV/DJVhwV40TeAOg7II
WrmRUJzfOi+xnce8gFHOpE5CvrdxQkLqA2GarzgQlLdcdnfEr+2UNPVJ7xEE4oFmuBNDnH9T56yZ
EFJapiZUao58PHEbTT4FRUaqLtUiqTNGTpZf3Wbrfvb2LzgdYThYIZeNd0n+KGHLUhVpfjeSXfIN
zFLsujoTPyZt0xjARnTmBd7QiMXogBegylaZNBDS4npy4Wofilzu1JVET6WOVMhSu4Gi5HcOga75
93/vlwazOQ0aaK0pJJ2HANdRw90sPUDtrnqVAeA2pVYK5UlJXWkxtW7Q22ZkzMPPtWg6ZV+c1M8+
5tF8kKEW+pR7NeLpumfnphG3k0VH6R9rvJsFMpN7NL32P700Jdin7SSANs3Wv44AzEWd3kbEgKiS
yL+hxx6HeRdL7eAP79/gbyNaV5JkVrEa5Xrc6sSj2/l2oATP3ah9sP5fUctaTNpWMgq6hM71di7c
QovekaYnJdu283i0WwiBv7U86RohQ/KUWC5os6SJ6XlDucOLbNZHRcc4C+Ys3Vet814EIOIMIhM2
7a774K3kcAHX+oCTR9d/4Cxb6SCQ7zUhCOJscMuZ58x6SOgtLjincxJMRouYK1NJgZLhABQ+NqJF
JoDbwdyhKonHYhkhRyQ87BmLuAO1R4EAxSFaGQaxpQUzVvYmctBiOqUEKlCE3lINlnNMhL6YQg99
gqXjm6p0YsDSSlrqPNZlra2JeOdi6VZ8GcjQQg0eZdmc5f2PhJHU9T2AOrQU0ejtjKOcXODA6gfK
q4Obh98Rk+sHefnW4PSpnAXKmKey3JI+mfHjYN1TK2SR1bk2qHBTlpUmOCXYZFFXngzXE8E+vErA
NgFzKGNRPMrAaFMZLx7dSXcZF6ofXGW+P8zOHjusGK6xuoePCNphuowp5Wa7ozFJpmf0ReuZyRC8
MCa6tVk0I3vzRJo8blZGbMqoFeSINMnfc0hcDRlM9lWoGXQArBvi7kHOrta213z7UEGH5lpbvc71
8JL7OvaHq6L5rQOHOJE6qBZMlhONS31kqHzcFYKgVYTzK3SglTNXTU5ITpAkwr4MQo7Vrvuyg6pJ
dH2PJ53KCAUbg42BCB9WUZ2/bHRoWxtf83nOCvVLUXZHOi2h5pdWdkYtblJyuvaqAnNjLOzNGbIl
V9L9S6JM/5tBHNISZBoyGwv+np/Qny4SBEDgo3TGRO1xplg92r8ZXcIMzW06y0iMbftxiqFEl8DB
IO7g3VqBlknXohBdAHINxlaiuzQ/3ra5C5IxYIbfQrLeg4vI533mAu8yB1f93PpEJcxMtyBjZM2h
uZqvPrfXIy1RhyVXntyHv6a6tGMlJRjF0mRvDGashDTQEzV9kjaU/bEr+eZjBbmGhA7vUnXux+nx
OJBNY3pOdlaR0MG1vEHdRQbi0CaOBkD78hFux9biSjNWcw/kz0mt8ACsKO0xl978YoWf2jtzTcWN
KgDILEm8e2WCf3RK/ltwoapNugSMnfFJ1E/8YstlBLmNpJfusbPqmajVp+bsY7wvSRs3NEUtigwM
FtoDEGFUx4LvyOOjeSpkP4KGS0snUMCbObENcW28ZCyzxcnDZlrDsydcIIH0+ljt+CyFg8x3gtWS
yAUFjNxwBLR91DXjK27FiL2y9fqiAkl/ZBfQ//hBZs64wTh0s5bxCet0Lve3KOpUhC+iM9PZQhfR
QCcbeuPnFy0FN25CZYBMQ13yKs7CmqlPRGkwblI8qCUxoTjJdLdk8Fzkw2LzXdnazCCfG5QE8alD
rKfAM4rWWgQHwcMdLw3SkPFEadfTZG0KAnKlBBLwQvOJ+RU2AaIn9Z0yqcsvggGnCvEtRyFaoiG6
BmK0F9/FSgoigHur89aI90l+DpZHRLw9bILQrtmnuYFc5CQJUcwG/lF5lV+rk2yGWIEnLdcYUG4Q
Z+JpKX6T0cQZTWTIo+lhs7ZIT816YmeXlIPB3e3ZLlKTKf0E1kDtM01l6hbNdPVn/3JbrEX/WMbJ
IwN/InbbTBA580cmmRRcb4GD9dAh/v1EEMuoBbWI0RPkuUnbuzc8aX3cvLBhEz1fCAdQpCa8CWym
ci4d4WBBWQXJxy2e6zeySAEbMJ5gBIwWX7j9dzgk7tQl3PwJVi047jG/Quk1RKp4dV42kFy3NoMm
P2ytEgTeUWwjkjagdAvxyTSl1rF+05vtcwvDfdfTxhbYKJxYC8AxTc26/bFa7Wd7MOBjp6vfjcF7
QDbjlwIfgakpFf2LprI/wfiLprWTaYMyMntqgM9dPdBkY8cl7lgPbw7wxmHpbYO7gjJHLZX7Tt0W
GG3Z7dsR0BP3CxmqWnP+P+jKxS3bwW7CsnSYHx25gl+whyudsQF8k5ryw8vEoCvEwjOUB7Vg/IdJ
0HGeG5e+c2o18cSNeVJi1OZKVANJSsq0bgA7dVYLoDmxGP3k92l8f/Pjodd5jJRehBrpZHJI9yn4
kMr3pWWodk4s6S/fBuM3br/EoTU1+LU2ByifZ+cL4dB4jdFPskJHjBDjO6bRozTCJap57l4UDGFI
2zqgs00qbrUsupOqtiXBNY6goCB8j9xLphpMU9oepgwZsO1iUaobtvirB80CsMed4u6+3VLwig6k
g0lJGJgkZPrdaLrwKT/dJRF8B7MTMNDacZqKVHmvf+nvmB+1CrEkwwc6cm2jLl4La0tEgNQJAcWb
sXc1U5urnpYJL9RjqRiIJTwHN2+YzFQARvqVzFF9yV8/xCy5j6/XkmfDn5tLjNSp1AoGCxxiNBWo
x7l2xmP1rWBQEkpx/wAhsukpqJ2VO5vmew3XHpSdfxtVdEQX/7T30BnAeTISroc2I9O6aeBAGSHj
Vt7zDTCdK2KUpK6YjEwS9lmBG5WmLuCQSJ5BAQggJPisAhiEQWl1aN9F5c4oVOLjhVgYWSkDF49+
P6zGLjkYT22fMsf7lSzrTkAS3I02FYS44u+28nh3XFhY2GfFLsGZQMhS2MCV+I3LfVcf06ci3Rsp
M2SsGvdjarpBd5c+FtoZUBer6v0Ed6ZwvPrey0/yrTNoQh0oBPmcDPqFSwHWF99kTzQZnHuO24Kv
3NBPTOzGR2SCFygBH2MM+u7s1oq9tIsHAQd8ZAP1U+rRGS9bCtjJ89P+lcHQwFx01vfzD1nra8mN
Z7M2eU6By/Gs8EkgKv3vkTt/wUJhbDdutbc/+s8WJa7O36dUjANq7mUX87UCuC9htbZFsHQEIVzB
veRctGOcXmYmQ92hzN7peD3p+5WU8GHyhjb3bFw+1aFA9D29iZTxFeOTnMDmKZ970vyn8934nN+4
E5sJSL4xG5MyLE82y2qD7ooYHUkaEQUOufuMNTrR6ujMsnT2ihrBjDVQht/IFiqw2Qoezzylr1vs
DoKhDfVI10O7RWdsXvhP1JEVL+8iM8UunFe1MY8zcEedaVg8i98+2jwko/RL9+sdlmB5X/fg6ENG
EgtzqZytuXouN2QG9v73EXJE1UEM3Vr1AMBLk/FpZL7jM/bsU5dAgb5baiUBaTB9pu1F8isUsM6o
tHUhevBG4OmQ2b0MpgSMySarUOZMgIV1++X9/S04+3A+d3hXDSY1G24U2xaKYN4TCkodavgyi7Ke
/RLUWk7a8h7NyWVnuD0y5erC/JTGBPtCpwJJDWPhBmcIzOnW6+2bYLrFnJMoPqH3Syb2OMHUlnRU
rLfoe9Fvn/Tr+7fBLzcujPZ1021EDbnDZUFKL1lk3WJ/2gGRB9GpGkA7AZqRwey7fIRQrtsTOoec
Wcd3pKlFDBQUngQtV2aEv13NJ4NxXaUaRi7BQa2+eVnqVoO9FiiwmKrzhlrqjSFvt1FLBBB3zLFZ
sSqyosCipuiK5VVQ03CNTFtdrpPWJu8NZ+qcAaQ/OmlGtJ/GHhRj5DjBZGkBLYhk1cNr2rDzn07m
1VU2IU+Xh5sY35kQBhmRcb97AjkKu+eO6bEtPbLhzdz8OLwPFmY+TxpkjMeocAG6mGsyU/7JoHMP
HRtFX4es+pvpiPNHr+rPSr/UrkHOgm7fA+iqRRfoV/QNIzaVC58+tdbAH7y2l7dyA6mVKgEna/q0
dTLbwOGZdUB9G2fl/d+8b1tv+T9aYNYMwQF/F7Pc/VcUq79jQxXlCtYvm1S7vXig15zEw7yVcNu4
jLrArgsmDSqqq4QteWtE4Q3wqGRxAaSb/krfykDgetkw4S5vtevv3Qlcv4IMnUVbFj/vxsCx9rwZ
XUH/GHmutUizakIX69JaPcXfW3doEw69uWhnueST/81ST3Yn4mlBWis6Wt9pu/u8KxrsKaXVDZ4j
hikT0RKRi98xFYkikwAPu+/+vbnMrHiORqa1x/048wQwHtl6MnlqVT9BjSdbyA+Z0ClryqbNHjcr
ngGuS0S8ETpwblEkwQxLXS+WZkMuZHdFH6Zlo+irrbFgIl4adcDUJqoVwikYBrWXmdrW1vK8tV2q
XATOLAd1rdB8O9pWyo9KHUZmVk1KDuwr7InIw4WnFY4lVKLk5sFskuY1XbvWnuGmLGJPLpzMg0Cy
CzlkcOsxQk8nmeb6Plenq6mkY3QGhwS4XlKh5yOA82QCU0jZys4fVTCbY8zuqiX8sx2R4LZUabLD
DrrNtvasyzj4VJgmtDxbWm/MAXCyMvk4pzdN9H5a+cc7GNnVZKhcl0+sKqskBtEghNflxtQ23IWS
Qgm0RDEHA0jV2pEzPcmDlcQ7sV1qrz/A5lmK+YWOXBYz5xT49Xz63i3KEeGi3Z8HZ5r5jDklFznC
jc4zbUJTjE0K7BTfeYlYZtAOL1i3nQ1s7MP3JAbrzSdB03fePIqPqa5x2GxeR7fn2828tKQ2Cdz0
96t5IonXYTCuT6zgfwkMxDO7oRNcN316Ru+LhBM3EcxZAOQYiX7chJCtS7LtT0eSR2UWV+aVPiXu
/QGQmbVXU6gRWyJFKfMTsrWW1yqAhmUPcGq3AbUbEmmnG297kEZaNdxa5G81ciZt6LhlXdLz+/uw
9BJtUs9BrX16sOk71csaEU/ZHMisFo9uUR01UQ00C/x8n7u3doR2XyD9ODtnVQS1mnDNQ3eEvOmO
FiOjGW2mveb+QlM7lCN8sgx0sYvD4YxDyza+iStoUYc+6onrgsrFjkmerwxc0SHEd7DrNu46MPv8
RbXH/kc+wFgm3Fnz32xxydbOFARUvgproU3mKjU7DNh5Ap5cQP3oNcGFn48ULcVaSUu3PfhdwP6j
wQKFr9pPHqco7K5ANgLPO8hTN+Ju46RzKN7Y9ziE2MAVTTuoujnelSdOuSvjh0Ma2jAcP9ezLPNW
vsxafsznPGNjsG8vB0NHxIF9pydpXVVK3ID81lkc0O9Oq0h31yi9ZVsNCjZv/HkzySZre2bD+Z3G
38SU3wrbdjvAARgB2IEGrMmqIqQ9ShCkxDUrt7Y6kY4akavKkGuqF6P4FlfGv7rYrSBfuRs1T1CY
5K3xzvJkoSOh15VjV0hI/bSMs9LEAFpTpeFgOvuMAFyuittfnWVBlbcLv2gBrI9xqu2V+4ENEkaO
hSnymdUMBBTymu+J9vNjAbnLeM0q3WbFpTdtZD3HS0ufQpYxhc1WK97q9QoXhYqek2KmQOcJ7A6P
RIKB6xiOsaeTvXJ+Y5MCZSqmghwwvoHSlLqQdaf22KqR0l/IgauclPSnqcrKy308IFIcDuWHs2JF
Q1iRzOxBeh+5eVfrY8cxuGYwm8D9iyLhcZMU5N6ZwXbY1vJGom3j4maiK0FqWJjTPSskLHNbPsSX
6M5YefB/kj4cug5+3D4pm9g1Mi2LdsySv4saUNSq7Qi105oE6Ju2QZd9/zkl3cYfW3XKHZFgyf/n
sfgCu+zL6G6eCjo+UzUg5Igy3V13N5qhULC4r4lG2sRrOh2geGyrQ5YS9k7RyOlx4hA/HwvuQaCi
unc1kvOoMcBqeAZYGu1h41n9h8+rY4kjDD38aU5OLUa86ZPU+XfPIe9Le5fxQxbKOhAkav1C5lfp
l/jeIl6sugjmf4TYAzWelMnOP2QR1G3z4wxIiftaWsTEp2dUv7iB7sZbL+b/DlfPbqfKXQaz885X
wKL8fumYayGr0Z/MZxktOuNuIG1wa1fvtQjP6b8A9ZBWFbRlaO4P3ytQ7JFmkdQx6M2cDoCYyTFt
HJhj176Vnpcs3/yRNpg6FV8OFnUzzevad+xuyYlYBRZg+suBkeq4H3T3UiJizvHzwKem2wzL0N/8
Jz2oftn3Txl3fGZTqk6ZxPgR3yBkYJGasc6CvHveXUOwjOejuq9qHzXtcwwc8cXpRlhzNTFZZP7+
IpMRYbdrzaf97Ego3N/b7oe7dGLcRGhxgsQMfSVEPKFqqBhbHe1KZ8Pg7pkA4hw/QhFaYV0/8kIa
NDnTeBwtun0y+zsFkigQHh8r27iPSBG4rswh9m9qFmivOp6S/85vYEc3ockOI/ODh0WRt5vZrZl6
jBE5oPn+pl1vDK+k2OkJmqWcDu7y7KP2jUteoYN+dx+HJNeMJJ02eJsRiZkxkzhqgs2+VOSJqk4J
23VQw8Ym7DBIBqoP3k/68at9eRvAaeLHJ8qlqT9GBNfTk/BbHmPkw9+a//0PSY9SlZ+Ahk2j7oJR
13jIpIxy0FyxDjZln5RMKnHE/amMrZEdpH6VFmEeAGG06nfWGEllzwKTH3UpMBR3j65BP3b4kyyj
wgGlcEFi31TVB9W89DBy0YInairB1gDlzMvHz8vMmkOoaiwe97nNn5wGnBAkrMmHKeBbDVrlot3r
O2uAkJ+cYNyFdqW6qQzcioA3gKah+Gv4BjN6jsaNcPtkI/yFjMXlF31ZtC+HDFk5tUCpxSNbv+Pj
DnXhNR71vn8ZWrQUCd2/gVn/48zgieXP9JIOjOpNQ+NcqTFLOiIiRjXePX46gSP6gjjxJbNRDRT5
tYPyyka2CcX3eulv/SNMvTg7EUqPl2dNIH3X9Vd8W1ksk7d3xGn80kJenNw9ymt15puolg4hGViB
1y4AEIaGul2jBb3Wk7f4KDWyoQ80yKHQxov1UNPYOhlpq62mNd5bpMfzM3g+nN+9v1GQtt+VRGtY
dvThkJ74mF5vsgKb7XDcE02p2Wch92akEPNvcwPXJBOtKNQ/65OWaQJo2O0tWQfKfC0IfUoseWuR
aBTmvowSU1wl1hM0ewGWggRKp2kIiTK8+0TmvvXXaet4j2Ewmbj0Rw5t5IEc7Obypttpuxz2i27O
MxNa68VIYGIHzfWiiFvrToVB8K+7U3CUlptkZNcv60BGa2l0nvJbZb/sW6P5IEk/jXL+QcnP5kBK
UyQdQuYIwvmVenC6D48kHl+JqxYordAZQ6HDMWRm3ttKJqNaENSLqZ2+vE0xJx7/vTAdiIR3hG5l
WhiMkv7uR9ERk9UExBYKntcOK/CFO5EXN+T+/me8sOIXE6S2EyY2nHsJ7bp75FudBjmxBlKflnQy
y9nCHSAzD39H01QRJu+y7JiFvUIMhrHqslxLXiAeJaDpFogI0jD8SuSqjkrN/tUaK+Tx25MjeAgt
aszVETvRYBtqrUVJ8KHXm6ch1MHYUds9MaZQ47FYhZdnDr6LclC7B11df2ClHI0rGDCI1WVzRNbY
B+R675QpnOZPplhY95QVZ64LjJrnXo2mYYmqhNyGQOwDhcRVX+eztBaH2q1UyImfoOlYZ6e/KVkd
//kV2qrGBa/JWa6uUjJskO/WHRoj4psCGVLX01zf2QSeZaNH50AP9t8CCs/lSelnzoA86CMrwm1R
sW1e5qLWw49T0pfCx7b1xSTcNQ4/X+C5/6RMNI/FSy+e64n3X+HNGNjROUat37PnrNh+jLQNoD8j
mUSCQZzeBVPmyoiJULHdTSVWEaLEP3WK8N75pPS3EF8UXjlgfMLCBR3Wa+5PMeMjAnuvZv0HF559
MpDm80IunSG/Ory4LDnbL/Ez478cRjQYURjcuFoMOHtb4nCEiHGfwYryRlNOAtTQBLng25AINMTP
UJSawrNXHu0lTDQBOQjOvEdefqtjALuVArqXiJqwFWEdJlza+x1UmSW38hCuIZ5xnd6W/m/KGCEJ
8gkBvE19DB+RL2cxoGoN0z2iI9mOd6RYdB6R115jjVSXMN0liDTQuIjGDnDegQrCwf4qYXGm/Q3j
uUqfIVeT1Q6zJRFx887N2Cou3FuEbyFNjpc3f3KFwLrORvYrxvHfGO6gTpqJGuqavtXva6ixq96R
s9dlnWQiziwOHPB9Ox/Qbk1l0mk7IFdOeJvWaXluRT2fusVeSROQY42YgXynCvQzxVVW9AprtRxY
Ir6Z/sL857a2b73OazeynfjUjtzOSWg3TfVQPueSiKTjhJ2q2MAXy674cI9b6oRnVRVZ9RVySrNF
+9AAwGq2YatJ04YDvdonxxmvClfJDkTFj2SceNfRxCQ+7YO+b75K241NPGidQL0a7UzydrZGCAl5
bsmpcGx785/dXGQN4cbxYQ+IQ/HMzALfLmIHLvQ/fvKQOuvFqkcTBIG75B0kyjWrVB+FhvMmRmRe
yhsHRUem3/Thd5ARKjmjUB0o2GI5NrRG7tR6rGNXT3VmXUCYgclM4k3Ck8/9EB5I8rhJKvGcP9Eu
eFPM/QpYtDupycRzKNqUIKuI72s5BaHQbKWNjS+tAQb2K894kt1K0q55lp+8CqzXH31VcVg1FYIF
oT+f4wrhBxD0TfZrTSllFuXa+gbbSFBWgbHxMRYBQ2Du8xbIlgbdON3YQRGiwV6ZyVVnA4jJKhb0
Uh+IPH/EC7BOfoeK/Oy4/1LFENHfOeA7JteCpPxOCNmfEl58tQxzAqaak7zWO0zvfU+LTt4fBSPv
sHb9GSBFFQqrF3l40AuL+cfgLdfT/X9tmyOurCvbhtJsiQjmw+XMvs2KyqMHowd3EY3OpNPN7Vc+
EMsL0WKgW+dnsLoaNVnJPmRjELEKVPUO1dGWRW+D+Bk8UPoMl4yZoUotXigOa1bTly0Ygdpt/49c
nXkLtRMjUq4e4KoOy/u6qiSLIogGduvMavI3RZRnRZu7MQA2DyPFt2HL0HKaxDGHXqUNj726xw3b
MKHL3KbYO0/Yd6g4QFBt0Ov51+vXlbsXT0Zcdr6t5dgTx52JbiqmzWI6hPulK2l1WkAMNYQ4iS9R
2teKcYRl2pFHTA4P4qFClsjnyGOVLb9Th1phbzpi4Xb55F3IyzVxvybzGV3fliuKC4tJwcEI0WQ7
saZ8X6t6AMsgD8KvD2WCUR/7dJeqMF7DLNQo19CoULo2LWw7nhAvO/hnFy3Sa9bdxUunN3swqgd9
YgBu8lIMTt2dTU78QTP8oJyr/dhPXpiiSSolECQ62sy0hPPVv3jbjYOZ5x7iUfR/S6ZQbW78ojFa
h78yslIKRdhgOsR+4zNcfPNaT0JEBnJx4hzouWk21lRFVKzbW0yg+0W91YUAKbXXIvmNyezsNIDR
8QSWRVgAJmi6EMEaBf1Z97OmlCw1FFMLofhN7LRxWC2Ux4eC7WWna81vxb3Ct5uc2WMEiK1GdJxs
uakA525E3BL6PDG7zVr6nXeSW873MPYVBgfGZYuchQJlrOuWO/cTGF8EUFF35MuM0Z6K7g5yCGJm
fwKL0zqLysmMPou7tl1snaYEgdx+MJP4qDaBy7GEPAMdDVjB8rv1kCqBOfiu/ftv1l6nHxT+IO7m
Xa+cLLHY/0p01ihj2tiPw2Eazgnv06Jpnf99oBJTSY2mvLtyxqcN4AoUq2dWJzma6DdEKAZGCttE
VxGUSqDRiCFm00wgAcreI+6T8vtiOw6+eLZOODahqJfSYnWvdYrbnXvL7si+VRN2YFEUSNf1AieP
7EsooR2STabqtOI23/B7Os2lDaBOR5UOQpUc9KUCTQDlrOnLnpAEegNH6mGMGGu00wDgGFo0Uwl+
lw7y0Fc37ngzsItqF6igcoe9ODEtvvO87y8P+dFqlj4V8Om5Mjniz6WYRPpKPZuQz9c4Rmu1/xKu
oiMlEmeS7TVWGwJ1qdYjqXbgU0r/qCYzgKes7oYsCogHala1Aou6ebwBEkcwHnxwwDGk3aOUUgX5
VX0dF/YvYrl114U3K9L+kgA5m/PUTpNjgotlEeWgAX0SGxk4BctWzNau1ZIojMmOXji0Vz3Pq35u
5AbikkyYIG4U9+oOQv3lQCCwmGSUvOMemWfeWZC+avX4db7E8gtyTC8sDwbGr3e7lsWSZsUZhf3Y
C8dgr4zM7vkgulbGaWXN7Uuksftkzmwz+DQT+ll6kHZDhQZ/v4GavousmNS882qTl6HhpBtY47SC
0+9yWu9dpNZ/5uT+JainFKwKV+wU6v8JzUTMQSNHciECIvsSd48GW/Q17I8GB0kiuESjIxQ8OpIJ
C3KA0upSPg4FbKW0CGiPcPUl/vEpHzScC/aiqGo9qIUhtPN1yD6CzsRNrdQh3dahq5PucKKcta6q
yAEB+AkBDMjVG05/AEv79qRAlyIfhu7hMRcH2v0O7v1Ct9gRexNrF8eCIUbh8Kisvpahi1WAs7bk
AEtOo0NvpOFEjC+R1tJEsBiQAanqBrK3M2ovrMT+5PERMu4Oks96xCWK6040h2WR5KVMUY09MdBy
s26swqjmasrwPkCM9h3kK4+320Uxwxv7YFyM7NF1UGzb3tGGtq0xNmQ++OG7DfWXjIDQ9DPsGWou
fmSnXjfkGSDANAwAVefhjj2KV2lsV80LWcp87Hh8PYfUUIiMMf1CGlp2ZNwC6xqMICC3WOOuhVKq
CsulGCaaC67acbBOEeBhvzK2x6RqRcmeXwMuOSezptCiD3gt3MAXnlQeGuUzahnMbGj+xQmGC1c3
jwCX4XVB3yUH6dCpZOc7qCvRcUyU6v71mWOsogwHL69/uvTUEVJexdmEQmIyaZ9actCRQNSUtccB
m+oSIC2B0Oq9sZ0xs+yHCm7uDGPyLTSM+i4d5fWmSjCHQjgb3bx/asUcMoG4nWkXURZ5lXfL6NFl
/EUwDpZsWYW3Pwf2/OkEO5djd1j2kNDur7kapPN9NBrkOrimbIT90NKR5xCbR6lLqp8rlb/93Inx
cYMOqrTxohzFQDubIWsldQtBylQipZuHWDPPI+mdvld7WoMBm5Zb68kv9mP3R3DkecMnEXq0HTDz
PAv/YKijZ4oSOu4Vk/1SVdHRfsHTOWjaBrLmb2FQFyEYZfJ757WoEK7n9ttgpfJA5Oe5OJ6hxN2G
S1wbAvGdaeSe6de7uhOfxp4Ed0kB5RjGNU4yXfjSlttf8DoUroNPMQHa8yLorEzuK3MeSQKYh8i5
fNChLgfp1TNmhdZrn0dWlBIVj+vsJx0gR4lHxltfGs++Drg/bd1kz+/KN0EZ1gJMsfOk9TCnPoFX
57CfKR5Jjx6ggbGO02+xO315pKY1z/feifDSoVYPVZM9P7bRIDBI7SzAaxirmUqRF77MpyLUc4mr
cGA/2Uxhtxc7Bc0RZu8lEIIgwxM32ejBCDIqRulrYhMIfcx9KtTVqiSZRpG7SQFrpDgiOwUvNlXf
g6+XUqz6ysBpLHJpeq4JPBmrx5OYlvqgXiVsQwpocxpleqYrzzA+CBqV2ID7K+oSGI3qsiKKz0S8
rJ2T6bx4t+S4fRPMkliRtKmILHAGI0HoNm4MHzbIYK4+7PdQ6c19Z6fQn03Q34E9uvdq1No5EqNI
/k2vFVGtBqBQr/reA54q8EzRmDg9k53GY5f/6XZGHvpkOgNEn2hkIqXxP9OOzOyZKJRqT5Jhpka1
Jn6C30ejwglWdiinShIw9FBX8iLOD/pYrissRQeL6U2YVhcqdht9oUgCBXRR6lHgNCztkUj8D4Qf
VOERWPxhuDkjyDz99PfwcJ91BAhh6T8t/xjDfaHmdBdbDoQoQ+7Qf7lxrprXQEZSziaDBSimRGK8
/ugG3eplmw4Phi9b4QWunD1VCvpRNmVg0sEVhM2A5xGPCQZ8SKf85BirRD6P0wcA8fvZuBP0PZI9
cn4AAaDS5FRl9GcjEfe5VRm6FFHns6yOFkXawC8tvwQ3utIg/tJmBKwJWRRbAzxBaNrRoP2ohuRp
UXokLU/Z9Tzabn67hw1XqkqHzhYG9mNEf0T93taBcWZDtlcxYqCSHP5MVdo0T+P+oMESUSTtB1xu
cPCauDevG06IA8pvGssWmiWONAlvduGEDSBw8kOeHbOknajEAcLd4DAX8Roh9bSHoq5o4wXAqBSl
lZvyxwxtnKT0M7nP4X5FtdVp6CLAb1cfZC0eQ+PqMEXYwQ7WxjTfnGO26fJIeGljhJdl9O5FwtxO
3vZXdmUQ/YALd/DgK25ODbRuKmQcVVg+nZSOV2kal62GIaN3XnCzb15pyfhtTqeQOFN+RMmwjtda
8KzHhqXPszRiT5/fn6I7veutQDstLg4aoWCrzc48J+30yL+i7oqJ+QdLsJQxUSB4OmooJRa1r/G0
3Tv1vnJxL6VXZYGo64fmmHU+cwOrYkFqEIkUS8W6c6ZVcLzh2EOJdPU/VYuvsi9tou/2Q3UDXSrq
FF5IH6MtKW3HjW3HoA4x4GhwEehDE1sFMj6USF5ngMZEEtYfprxpqyW6yIAnmMAW8DsSyBhyZmZ5
fBJvZMnCgH+lZsSVEB1dG/ixkiMfxs37fdWwM/wq3Hk9TDYfH1Luwah3STHSkRUYysgn2nfTtezR
bWVwfF6piEV1LJU9PEYke38Ee2+3LG69zqPWBjimXqWFc+uCah1QW/p41XVE06u+ZPgylRt0hTYI
kNcTP9qIROtTx6p1sJdOCHqDpVoeJpocX2RolxEPRoSwsRzOzVY3T5Jv4a6KEuIyDgO+xp0mdD/R
01/0kbCMAMKegVMexj+kCTcdrcWUXQ8BSWMwfYpID+wdCznUVPyFRklSFLzR8v4WAHlH+aV58eI0
eASvUr8Imm0Y69GIzf2rJvIjbdcJHB2X2FTX3BDBrldnxrvqE0Cerg1xVt9xCoRADcQwB57VLyJ0
5LERIZQa68DFbxr5E9/9GASJox/2zl053Z+uQudOG+kV3VMn4+WgcQwqVqANWQ7VqbvSqsF0DG/p
r1t6QhuPWnDGqMYod12OzisMMWGUyB13fNGM5r9ur3eMrSEB1uHRYifaJBWo5mi0NNpXwwtfaq1u
6tY/fHHRiJTY4yU1gUdIEliecy96beBAjORvKnnPboJuUvC4l7kfsIjyBbgXMxY+gSoHtGBSSQPw
FV2rfunt7MUkCW4PaLe+ABXSFEMi5BaYtjwaV1cS1AdgkrHU4hHVM7hwOpCvug1OHY61ZdYT8u2x
GwkFh5aMxtycec8E41q4lfMK2IWUDP2wj7Mg/QW5UqYBePBbH4lrJ9YZm7QIJg/2yqNXvV6oQRs2
WAH/6GbeaM/0IDOJveEY+SmJC9ZCrI+/XTu0FblJV643dFztxPHHn5WJjLAlf8ju6URktD9V3zxm
pL0mobqcIIHm3B6tuVCHPluJMxeYNp39Ft6fnJByVXjvGJ6a0nYOaOWinrUwmScOLR2HQcAxGRGK
zvywbkH92/9fYfI7WmHv352yX+IxSBrBYy5tf2OrDXy/8ScBsuPOKGv07Gr+1gVy0XWQ6c04yYvt
fTj5WRij5Uss2sIavZDaXQnBVaI6zd1QXPd1cf0o/hT111LrAbBOu7UhKEmetLk06rsP6Oe7qc+O
UV6dMRM6chJzUom6sdKGY3PnXYbDVSSLAFE4JacDc3FywhZnJJ7QCBPRo0fgClDeIRBMLvcxH+9a
ljHgByZi5hqXz67oT0RozQuzbeGFrO9QT+uSdVRAecBHAtoq5/J71qdMf5pYp+MrbAkcVZ37m0Nb
Wla7hCLSTR0P/0DuWfD8BALU4wlYWotjU5lpDr1x5TB5rWZ2gEfJlmk0xd++rrC/9eM0YFO/T1su
D/l02+hS5vf4+OHo5phDbWGZ7QraFUDKq1AztaatNRvsi1ViUCXVaeeRXiPOaGxaVCyAfaximM/B
2J+7XjLymlCsW3Kl4k6AzGK02IrFttrSIb8CimXLfHyH3Qm8w9WM0Hw5X7AOe+r64LUVg7aYRWOk
UumU07FjMghiNoeUguDVQt/K1tcmGK7Zr5NNzv2ETIpXkBmGotdRTeuq19Y298F0pMcoGQVnGolV
IxzW2nHnFPW3EFECVbW78fNUSqmTmhFUMDSMeKJzSdg085m7cmPilfa3v9xfURF/GwkhBbh/ZFRE
/bpczpWqxdBU8UpmWrYxqJmJ8IQV0zIzUsDqjQ/rj8UpbcCQUAoouLlt9QN8Uhl049rTJh/FT7as
597s0G5E4ZWe4wiFFYXLE/O8kTtfJYU5K1Wm0A5MCb+0GsVSLJhdXy2QERmOH6obQpm2O2+iEiz6
QuCZfS++byfxO+hpxFd/2xeNE0TJQwbqRgDL0Q0onLe2rUgAdmSRFhRoiq7yQsKewTOp6uNEUpU5
G6GNB+xh3wrw3wRIlDPPe6bQ3kjv8oGVNvBvLr4dRHTOuFeMrZz0BfUVlD5sphODY2164V5j/Kh3
0jMSA3WCpu6+KULsdEjpophIAFqbug7HFDRpsEPGWPVk/hplW1wvwTIufNaE8ypJm150AccvL29f
pUIUBus8Y/LB0CuQ0mLz2qgHu/DHq/P+0XGuLfWFI1g4Ea6Jnj//LUMx5XQpF1PGhToF2Ik6UhCd
iBZDErblhzhpzGZnR2Oxauk03EMRIVB93q0+2TfcGSqGs8ZVyeCdFhGnyHZgI6OZIbkpQLzKeuPU
MdQ+1G166XF2Xty8mrluurmxpza7acswNbrIeatj6MNO7FWYAgKsH8nNP8h1wf9VnKCrMRQh50eP
4iK6qVw8HiE8SFWQ0urP38WycbdEGTxrGy9Dcv0EitMeyaC8Dh+pUfzKCbSnaY37OZE1bI1eCU+2
UWyu/p/VckeczF2wOJHjvIg0yovzAfZlcAzbM018/vCAXRPd6NPWhLzyDMcjSWpJS584w7rbd//H
sPZ/ABsAQyCbRmvtXKq1tOR+YsmjWpFnOZx1zP1ndBSIdj7OcbPNvR3ofLfbs1xV74h4LLOjSAee
JXazral3R/SDoLD8XhLpM1Z2hHB9MPw/3xa/B6+CkdevW70czAEXflV20/CnA+jCq8x0tXiwVN5u
aA0nputwBrFqQCwy8lBNxNPt+1tuYmLbCI2kqCx8/BkH0tdKkx86eSqKeTGG/GA6wqLtSMFAvUc9
twlYDZzwlYttFO0ELvYlK4I+XVQY6MpLqPPF4IjyAAgubmIV2rRnuR2DgKp1XBC4FCSYxG1xMo1h
egRN8sWE1TPLmtNeDrQ9gLe1oP9pMq2SbHm7gDEg3gMMmB5TaEiisiSk92a0T8ANypD1jsEfp6SI
oq9JZK4DAT0b16sRyQzkBv1hOLScaqorEbK6rudTpouQpHQJQ/JOJjMjKEJZAgcqetBa41D5c7C+
YtJPF+XF00Q5XqQklHnsXM7vmpaAvZvHMQGBOCLg4P87j8uhkMiGWKYyyghWtYUOaXQSYtqDzAKR
jb2CL5bGwcZb6ZrehYHCkgvouuGoCcF5BvCgry5urgEt4gQogeY3hQQsT6SdOEnV5I/yeKPvp3Er
trAdd3/sRPPqdN9ippvljmImMbHLBhtK15zaeVfuu6iWIlhQuv8JdMafMjM0ghmKJ6AGITvlQmua
/fk3sdQJC1nJ11GpoceUBX6YutVUWJTHeQk/xxk728aPrvsqlOUm88yuqupa0kaPtrB8boeUlkfL
KqQfV3NFUPX49d1pyayrysCNii7X3hCUFaxg9A19fF6UftylzdSA8hV+zOBXdKMug0dstbnMyfQ4
agbWUo2O0hfuuwoHYok/4Gfem3mVbgD4hQmrcayCGByruDrjW1OJCjEyOLQyEMN7EgxQj0cn1ZSA
l1j4eiyGYLQNJn89zCEeLdfhHtQcSrqoqiz7Hvul5g1bIWL7Yx0g2RTv3R72T7tzgEi9JfHyEH1t
Qd2xcJwd+oc20XOKHC/g1gnaCuNtid4zXJ10Zu81a08jQQjYapIoG2Y5Vz2H1r6CX4PXLsG/tVxB
QWMMEo1u4x6cEyQG639jj2ehxEbCLhAt+DRYBFdkhY065zF+BqNocbyoDKLKd1z/a4MgLHE0o5xN
3WKK/pBKoM5BKdgiDzryWXdP1i2Qp6CBbqRJJLlkDxbg/YMT1EnsIvz3o/U+Ot7oF5K+lt5Zzf0s
JzPUlvRTs1Kk03cWonhzoQ64YhclFYNBWGJKTezHij5zP7vEUBtgWGqyjBWa/eGpbbzufYE4VZ/3
SjaKQGjc9NvTieiPL/Snfc3QNPtaXlw74cSjFBuMqtyom+nF7DdnqBL9UC5rN4N2R23xuSLLi1Uy
34JQ8hVozD4lT7jHvmJF9NVzj3fMIZFqANlQXLj+4tN10yEq71H/ahhWz5nb4AE1tDV0Cjc3uFjb
nHke29ePoUjbymSpmZEmUTx049GPfCkea0SCw1eBmtD3aP6kJBmxMh8tP6Ak3HjNFQm1hIqaC+t1
eQhf6+0OUfqrteDExka7FMjcKB2z4wBJjlXZ/f+O74rsMl6NkvbSuAK2UQ9gn8zP6RgyDFqM0nZh
8dYGxaIfcjsLbSVZiMQK0XCdERBUOHX06jzrD65a5ECtuO9hfWh8k/yK8r0d+EOaUg5Jvlk3jgDR
CzQe/luSgzINRyMiBUb/nac+Xl7ZHPFMwvoeTiyfAZI+0ybRxDhRIT2PihT4R7ZRy5HbW6YHQWJo
IjxZFwtGaO5OTw2MsSZhgmjZ8ZPbq87BIVzn3BSDXuBK9/+u2VSGuI4g+TqXxLq3KIGk+U4V9blm
3ZHxyFbprmNIbl3sdy7+sWSKAxYIBm92P9OhcZ9Sd1fOPsctSVA9CyItVXKCzk+DR3qxHMnUEByW
WBxX6RRKhnlVDDuA0Tsvt8X6YrdPhmgNZuyqCU0HF/OvSs/lFF8F7DRv7AmXMWLGNi2s+cAyZFwN
Ml1U+X8Qb8OSPyXtW52GZ5MyhqFasuokdAlB0TDvX3AN01tuu+PO9EIdGNA8vKOHRZf19b93Qbd/
a17SHvq7VX1EwO5xHukJzUhGy0JELiqlxr4ZxO1L6riZoGPmYIuCBNETAT3tKFc36m2ixk3KkfRf
GYOy8MkGr/ioA8LViYB4C3/3e33WwKpfPvgmaMg8IqvzJPwUMD0KR7OQLbOTTyACol4ZV1/DF84K
0j1APZ4h3Zt4KSWFXQyYfha5WAT4zQ4BYRu3GM8rUg86NLzJXlorlMNk/FINSmezr1r+xRsxqKo2
Krp0orb6phtyynYR399fQNu2Cd2yfMVB68eIGUpVZcx+S9wyqZKxCmLAbKuUx77SmT6Do9qR1oSn
7c3RumviA9Jk2CbhBxS6fT/we2vRDPECQTbQU3uwCtRoGthBkk+mUn5dYia1W/pamESX+awB2KUr
DN7fLI1Rwvwr6fBA+EhJvd/Fg5XANrWSZ2thTlYJ6kaS9X1thPjNZY2ySEVM65rvAX90tUi85v60
3vBPS3rlgXEA4Kn/KNU7Wliz6kEuLEUUbxiW+ojM2H/3SuONfGXKnDYwWWOSWqRKBR6tNuGkTuU0
bDajI2FgTSIJsiroK2zmdgCf+gtO5Sc48j3r7nRqaOQtIkLiODAZarWqrnYvn9BJ68QwP98pJ96o
yl7160B6oHrUP/aMPRNe6RxCURbSgVLbVKq9ufm+fC4sRqCOMXfxpq8dh4zyEehDcUU4vOmudlsG
2+T0h11npV3v9tlXUzgLRFYyxYNAz5fxrr0/Mgd2BmDwYnulH+LaaMMSc0QO4zJzfe+iEzQyjRlR
UAy97GVFe62XbynRNZksm4O3gAm0CQF/jzPQO3uCbHVhLQH8ZVIoThHSRr8+NXPDbQsVuI8ZMgCI
Ef+53n55qQsLA32eGfRrbyR5p+WA1i0MVP2GBWnKCvzU7qyUmvdZOhd0QMl6YA1tcJ2tMH+Y1nok
jdCrzMa8s1CNQwPpLzMaPqmfpaD85k6GKzuNdRm12VVYUuevVQ+vKoY6clk1CbNGXlTawTui4n7g
zwns4nuRRGaWOqiEjQQuKqKsS8pdFCXx0IhkA7WkRscHhWz2ptNM32YhwD4xq9oSOTksCYSfLrU4
+J3CcpkIww5AtTEY7/eRigSFxeuZ3FPn4vthdQvakr11dhCqyEp6ZLCfVKcSnsXi6L01BGDxlqg0
NtDBtAOnl3yQGDZUUVXd1XdQUqfd95XBj+nO3i27yt/n0fYIbbTaijDWRa20OzuxzUMW1Qw1z8Rk
VXSDxHVgV+d4wLshY6foeC3K7Zlh0aliwRExT0UuqDecaF8kQO1mPiBwAHNsh+SmqBtDWe5STy7M
UnaKXxWC3LILK0lBUxM+l2IAxXJNOjkmJb+ri3vhjurvv1lV00xsY0GWnM3lyKPx6hv/WlKD5L8d
KjATvU1FtFILURGY2Vl5J1tRVA8JkVgW22UCPuLnbGe6E90k9mhnTzbcDQ0r2TxPKOuqmSkDgNE1
Hk5s+HxwD0Fiv4W+cNYEa5icN1Iqd8sfYeW9Pdf9ETVB4moJaNxPQYsz0oCRnsZSypDWHa0lko3Y
5/7ViJyGmQFqOphu6nKRxi9EbO7bUeTsOCjIbJlUZMeqr+dj8jA8ENt3Pv5Yjn3O2LGNZ2SFO9xm
rB+sq/3IbgxljjfLY9jF0F627X2ByI9wmk5rbVKazJqspo1E0NqVpyNkeJQiZZxmwhP1RYcUnq+j
bbJj0M4zOMxjS3ManwA1cSY5ap79MpZrKT+WKDeTGg9bboib8z8thxsN2mY0SNKgijbhUGo9mk2P
Nu4Vd7js7r78V/WQsrraL1E90NIOVfQ5e0tbLW9Vg5N117tpS+ZafyZN2+9JCMdiIwthWc6d4/U3
V3wNEhZHSPoHm7hYN6XuLkFakvZjxQ7jJx5YZ099DFZIP3VGHHNHoW33xpKwtrIY6zELSnBKoHX3
yWfSGf0VJgK7DrTNlC0mUUA/avyMA5k/x4WgeGYvXYVTE0Fj0oh+1Xwk3j0m36BYFgMjFWOWBOgE
IGuhFK4K6QYx2XCImiaETLGGmBK4LiW7Ay60gEVU6wAW3oOI7uXZLAFI42TBTSBYeuo6EQDtRozD
uVl3mo5j4oWXR9P6mB6CIbSqsZUpQdoQHVOpkQR9eImKmMTjxlevlHeqWo/uV090NWybFnwMCrfo
IEhVIpbrkZjusSx0bI3NQeL3QzblRoPW/qbkXxhnbpIMSrQaEM4IUvUqegtRmtPDP3DZ2Q5m4fSU
4zrmiAECGtSXda6fTPrgM4WAm7iEMBUHNxx4QOXwmR6Tc4nsTyiwekBoIh8koOIyFPx8QCsQqTcs
SQdciEGNAILfesxSK2PnNkbCUT84qYoSRt0PEnpV1qgpmtI+T7XeNngEuqPRHmnEGbH+r24t13qf
eiXyiTlKDdlC+cnejAy4KX7wjDs7snRxr0Lh/LfRpL0NtdZRnIPyi5C9B3+A8BJr1B5AsQ4hJcMO
Ed9+xRnRoB58+umitLiDrCE+WHScyHSSrljTlo+jpqyl0Cvt35hnugQSqewJSn0jCg6UU2+d4Xts
lfnm5tEXtiPj2bRZD2XnsRktABvOk0JJaEJx3XujhoolpFnUXoD2u8RJ3FArrPD1gC+QMvjZby20
2fNWq3hXPcauqnjQedqQ449s6DH4aoLzypnH6ym/VKQqF/uJ7vkQLe6LuKPr87ne1dNJzL+VFUrF
87HMZZuS/HjChaMig8mNmyWNz9xdjntK4IOsbC3Jy04QCgMCp02hpJ4Vg1MWNG4LQcXXhmz5w/en
JOlIDD3ZX2LCXqfaAls1FHjDTS/MiTl4py50bzWSfZhhocxc7sOBBdRNEUjVqqEBDo7mhjqG4h5C
5FRMySwBPdH3NPWKH/mf9JACw3VQx2FOmD9HsYU1aLqE2iWwZeyR3DEucXgG2t3WYbLY+DrrDPIC
Xmt8rws+765Xxntrz20HKUTWWEkaAynl+fMDibA5VC19n/hN2PmdudNKZFAYeWCgOlH47Bz5nbw7
xTG1L3bOth7rkg8QEfTT3xwN6iKGwNRNg2qlV+ZQqrEjVYVwFuxqQN8rdTMWToiM12x56FdtZVQe
xLv3I19D4uexyjD4JZC014ZbrF4HqhymhmOIkEoe/vzWE9vcJU4K48KQ5hjWf6mcYu/NA4NZAg5p
ZRb2c2FpaPRP4o1xuo6FRlcOA0G00x95IGdrTGxoCQvLx1DYkhIDQ3c0rHKch6KUMFyOem3ztAK5
SmhSa6G0lsfufwwYj96UnUsxMXlyDVpdyTkiWB0MyCVH+uC/Xvivc9UFOKPgACqMK/pwHGqIIKBN
ENGWGvMqcMeCAm5CmII10jrsh5vbkJZphR/+R2uslaZ5UYi96tmVxwOVsrh1szeNdWbRcl8TPtGa
rmJprjqARPt0C8eKgRWkvIOJS5Essn0Mr2YLcVgQrCSW9MKIGFs7VYSxcJpv4ORMATSXVBPYTx2h
2xWDZuGTB0KI94RzreV9P72B61Hz1CmxxTsgTNIaDi9ryphjM6tlL1MMll6fIAkgSKQUOiKSElq5
Dyy3MfD5a2CphnkzrkyhQMzjPX7lbIijKpULS9hgXPrKMHIwRrF4blm4GIBjxRc7bTnqhP4x2xbw
Q4Ty3h7/ykFYcjKIQ1+DS/0ffV/f/h5tHocOlbj6NYgaImWvsWLHvbRYKf1mGjYwMgGh0VpW+Kmc
/GtVgukLBK5yYKhjJ32qkeIPM5f0QTvtwBbL5pzWpqLPtsDxbOK4Eoz2ECLk93DawrTgLifROQQQ
kIq5QJYvW6HKEnLyKquNO3PcxiVk08pmyhcDNfxx+8SMopEM/IEae44kGxt0R06FQZdVQzYbFWRv
/Lq+VTcZ2L5B8+qlgC1+PFXHq+wDYJ0C7lrTqZSfZyeRLxlCUB8SdsYhO32IGz+vR1L/wpIGHufS
/XQIMuK72RhGJKehh+APi1TMOLiOOWW0HnHG5a379H6OOJxjinRQT2GYRuPZgDLIoIQ66V7Uo4cq
HGvrQBhdnj2XGcLpQYrXtpgJnp1mcRHdr6Dix0IgnYnyK7RWq5Agu0wfE4AW2ACwB+RnHasOfD/t
PJPZ29RMRtqG/h4O8wKtopvDRdzAyU6UVQfkeyQUMdZro53SxTSAOCvSaiKge5UiW+8g6qvexO4Q
jCSmmmTu6xLDayPkDpm797XeJz8lBjNTOVJxbi1hPKZGtTGWdQ/IUeVKwiesbzChkWrQ46hIHcKC
Isi8ohFTIdRyy8OS83JPBlGyG4j0BAY3VblYPyQvUFJ9w9cmch794pEIg1023UVdW0nGQ9N2Xm4e
dcWBjnEZs3Pq6AqB+9RJd5ijK5yuOU+yUoOKw7UH/5CKRa1k7ZuAyMIYhviDWbjfs1mCImJCBCFg
nAl5JOn7IgpmZ23AhWvO6tEzLLds8LLENk6n/8IF0PZhRPEIiZ7TsNZc3S53Roauy4+399VSkDkY
I5wifcyyxG2/8mmv8eJqKDsqSbE+QateGAIDIvtngMwjXmS+f5eUklCJVIa5kQ84/YtFvExTyOgs
mmI5Gk7lJPrYa4jhRzc0W5JZlnBgKM+t6VmFUiSBW52qzBWCdWd6B25/sBRLSmoSLTkzr/9GWp9k
c6sN4AGMT28gNRPbwLMKMN4rxx+OHOJqaNVJ6Ic7GBKQac7yAf2JMsHYqk7/qzjZfCNn/TihFE2p
bjeHtnglS7c3SHOdylr5uJNK3LKQPa1nEnSh6Dbgf/ULBaXjzdhR4R/7Lh6zaMuYrxdP4NEZGoJh
5/1sl2FC2Vf9MxZf0t0R3/jNshiU6RWbwa4Rrk6aIjS7f7Sb6wxgEaY3Ukqed+BBApqsC88jRpLP
Z4yjSSVJQ+N/E/KGMJJvEkmh7EKdhm8Ep+1fJjETtcU6fCJ4fHKWlV19SBUuRwDgNhm5TuCrDBBu
110cSpMe8G4rz6sZ+PRXhQ/Q1JIQGyNU/SoH/pI6bt3Fw/W2GuSxbnd5f6qrLY42/o44NqI5dMDw
pt4Or0f60lxlgeY3sUDdyKZtpurihYSX5yA0JUnCib+tmNhIGt7uPOUYd0ZVFsV1vEDIuKAsQJ/P
4Nw81EFdMYzjHEY521rUkWICppZ5AqqZeB2ehtAIDZuQbfvmp6XI3ru9nBaqWAD1Hlb53tvioWpM
xC8C0RzdK4xghJNuw+PSPchKO8n2mV5fVsMuxXRDA2l1iIT933IbTvSr184Z8L8mPsEZoKFogw2R
42ZcQFqJKYUVj7S6+kYVnW1Dt1gncVpsUwdVfxMmva4Xxc/b/livzLelJ0vbaDfrwRsJcBpluNVv
2NA7x/k36uWha0xY3vH46rOiBJ/CY8i4YhtpfjyDS5+JWYAkhWBQiCFw6aZegmBlhEGIfoAvFHta
Zf3yVAmaCusbh825C5MZgdIYJCbra//qNhf8X8WUrXhBEP7o7qFYMtyv/weUB+paHkGcx4uqrzLO
pYKzJWqbHHwG9qxpwJb1DqZSUDraPjqSgLU7ggSPFGhWjxfjvQ/cyrPBh7e2Lxj4fcGqHlgLldq5
JHFUkzyBty4Rt3xZpRcy46cKXdutnobng7XJdUiYOsjoueQvonp9kNp5z1ZaPHj8kbFyADUiK8tf
T5ewizpvS0CWO71wlj49HDGNPHO6gSSBQfEP2EjCE94ObJqBd06xZm4nkrLqMf9YGcFxDlsbNyBb
aOT0LrNrsFlcU8llwUI+EbtCMWbvDVHLzp3xRWy8Lbos9Ku56me6dNtKv4DT4/nzCm8aOKiuPsui
vMJV2RyKE+DU8ByF2Ok5JRW02B42ozx+xgGFEdgFnj68efNoK/kB3zI1SE0rn65QlugPcuyICNfV
Hv7OXuyHUjU5X76dRKuQLSOYhbMtqmI4IghvsSW8OUrV231d87RHJRTSVYZzvQrYBm/bzrTUDt32
Xm2jI5VESSPdbkJJTKJFVV76rwezzNGDi1uY2Rpb0kE2Aq8AVpHv77/6wZ+jJrzGPSaSDvq7WwtG
OEed6dSoCDIH2pT93Pu5fQ6bkg4X5ioy6KuYM8fNg/1FVeAWRyJuNOA12YXeUANjtlRazmpvLCsg
iAnv85NB8ESamauQV0G2dckZktroU9jx61he5c8/WbU/wxxog1EYy8n1Dyr0twaZUfllsG51uz9U
sGgAX5LuTfGVp3cr2+c3hihNJUIdEQnzZNmifVDu3n7YX1irhax4X0qdnxYXmJuDJizqdNj7DCUT
yw40nRzy8r3p2tfDhmFbHw/b+uPNi/snginXy16ywnjKRc/1P4bssDjz/nyl/0X0aKNRWj/+rCq5
shEvFpVwSk8GfOpVQM9J1qgI2nZaQXKOyTMz1G8iM1JNtV1kjpCi94aNMx+ZPKtvk5DEnEeuIm6Z
X1obtSyNfejKFU8wcZen9p7GQ5judxVZ5pxF3teVWOsCpKI0E79OhlHIBZN7ZbK2nPZbJ3USKCv4
3agCRmMJUyVmFF2klYP289PdysQ+DuAWPh6rIcPwf/NfRkVTg1N3HCpPi6RcebiAutNk6QUQ/Rk0
dlKwUUI61RgZPiTzxkNmLmfWkN418hoXN7I+ziL0+vxnrnVknDB9dLJaza+UlYs9qWckvD2HrweY
Pk5PU8g+KKAmngOZb+YyJbNNhzpO9C09NgBrtEK8ia3yqWFh9EsSLU8QKWBlvaZ5WETrjsuEUM30
yzUewBigMC8/Nz2CEihx7qdjzo3RYK+ZZtfa5GIRy/Enc7MQoj+kL10W93EXSXKDC/Bza4PVkmCI
lex74mFlYmmNiwnrZVlUgoFYmK5INme5G+/g2CwE9+tT5xNn9e9iUl+jHfk4pOKsQYMOI578n8IN
BBHIt1cT/h9lT+d8U7EddkUR4t/msOl2zrBt02xDgXYL89dflXYbee+r8mTRBEroVbZp/HqGnAgb
XNI4wugpq8WuUVUxAuam9j05tQO4H2GAURYCs5fEHX8DhmWyWECovOIJD70ryc4ovSTYJDGQGIi3
/JyGpgeTWx5HWA7g59SJTHBBz0+CkBqMbDA8npeMbrx3pm2TRDphaZX3DOBBQZ8s9B4fS+mxKYwX
7FJEL4PernCARZqapuAqzzlPqLX1gtcYTWfTqQfSfeIb/+oNb5RYt+KSezqTZ9lhiMJK/3tyDF26
1faifrCJX+gRYtyvQJm2OweqQofF0nOD9TOlhwCjbRq4sbziXyPHTC15ujJgaZaYyfcxrDyAKyDk
ldn0V9Hpk/5A1gOEfeEi9icZYNHaWK7zbOE8s/llqLqPjgE6tAWBP11pjZexoTukyOnU26ZZdtdw
f+9ZPiRH2hogc6tTkcHgcBheJmMGQHcN2cq5HmNLXkuMKuQYZdEgU6nAXKdRMp20H9yhdd8KAyAi
fDFcS67zfsXQsUE9NeRQwVP3B1jd0vbBGavfpc6bBboD59HH8z93X0+qRyLsE0ot+G09jmptOdpx
7D7J2gB0Px1xAwuN/41+HsRKlhC6zXayNP39SO29dSwFQ5TvJskNG2PyUaTBx5xKi6697S7jkOfD
DtariLGjX676Gr+OZkSVrSz7JvAIjmYGghRthVAl5EDh6n3rVFZTUjNAWJnPLpnWXNy2xQcaCF4K
nyRP0l+GVYxa3lNUa1AGKda/rxM+qhIQNRlrqZcF+ScCSUPORZq2ETx76obkT0w+mTKodXD3V0V7
G5bwXbgxIi/zNgPyXmI95IWWIn8aAPlYxJCGEQ4/h1pxZ4RzDT7hjkb/Q+NLCUqCCTKjItNnMis5
oNjIRIfeJcLDLQtbOq8SMBvwbJ+T4p6qWQ29c5gDutdsE09bSOLs9kS9UlUq5wV+bJ4xm0HaFkkU
tCPpWRD43yGVPfUWIKSR0G55Jjs7zH3CZDdGmYThqESkJiH32scoSW4zhDjFU00R2dOO88tVCIZd
qM89Fev1e3j5Rv9u585+QvlASvfoICXEPzj5yQU4iQaOIRDlYZ4/oEMSIY5Vfi2oKsc8WtYzmBW7
3/nPLpDgBxKkrwAICBzWcYecxbCUhGfOAFBWyrXjoI1YJhIWpxreDq8zRR0rlUHRp6i6eNQuFJ0Z
OyA3L8HKTpPUFGFPMK1xpiWAKQW/ju/mVJX4Tcnmoo1TrqjWA2v1KmTF5nYorIcxtQT8D7Wjaq5q
El6UiSRN7xn42wEsV5DGCgl7cIT2Zd2mDqJ1nMzTfnGU8v0tidr9aEwBHjFdmURPotT0koCwLRhZ
wvkPsPgaAxSsKT3vDg2zxoDL6Zbt8NTSR+LA4QHlBbmyHSuiRW4oIbdqB22KdseXEDxfCuiGITRL
yLmjGSM9/d25SU8LeQ5XwNaUHkKN4STSXzzcY1KPVPVU7HZi/I/DBmgEiyw+K/iuTvpS2L+Pb8tx
Yqv5eihpMv3HktnLqvVeaZwG0d+056iXS7gB0zTKheSJBK4lCKTM60xP3OrmFJ14UCUrTVEjZNg1
fAeFMeYDoWh49XvUzL5GbXTcwC2w3f4aNKHsTJev50328IwleaTB+rvj5/eqUumNTgj4666B1fXX
sjJIiMRMbUCuUrIDH2VWnQ09/sjRgwTfhkAljWXs4Ij6yRgwoCoUyBRnzp/+6BSkIRO0Xd0crTwX
95EkTEXoIqUMqTewznj7vdspcsbrr80M8xBp33ZbAAVPMtF7TYkqVIMqGTRSJRHdjPEADrnra7DM
vv0TbBiuT3dq8UmsmHnIcp+4qRlCVq9uQYiZGDmdyE9Tn1fCzcmbto4Q4a4ovZRoJnmPX/VWUJLq
2bIKmhMN23RK3U5Wv7CE0ZqY8CL6NaABal2aVJZWgGZoAJStvLUSWZZPm8CSYYvjCmf5XK0p/zoj
ZLqb/JxoW9Q091nlUczWOEN6z+oepNeuhMxJ/nhfAKn8n15N2EIV9s9bGUN77de2oR6dmBQL0+Ua
w2ZLah9UCFXphWYGYvy81v0xL4L+9yBO8JbwP9iOA6BCZ5EnJKeljzpl78QacJyAWJV06VtX8uYW
pe0zynvCNrVOXmMw1TGKECOOwCio4QzLoGUE3eN5o03Jur+D/hCjdJzrWVUWaqFh0uWL1GV5NUTd
kRhx6OgobmqVMKP9VUptxnarY7kGYtFNujz2wr5bEjo4dySOXhHUl2U8Thf2odH1zv5agvtdL1EX
HnT0+OG2Wq7w2i+2w06Batx8DNqwJCnTuP5gHnD7TqBlAW6CBG42M7PLVCSUAvzzJeLF3a9TGMoC
XonLPSL29vPDiN1M0/DXfCEGtUcVLMDkKrSZzpR7LoB4p2YUPNPiKzCw5WBg2nd7b/lvciMkouII
PQavwVe2kLZkvqrG3DiTBNLlhoDxR1X2zkeMsMAbuF0dQmVWBSUvOEka4z3lR6FZOIZXqMNmORze
vlHS+IzkZ3WgZXwFsW+a4fS/74M4EvSMfN0Cw3jgj92vPFElgctSwPiEZXFqFbmvMD9f1743TsCX
nRW7ALEVNFuACLnGUwU0PhSRgu8pH/4sh++xUG7IMMUtGFhgX7rMTRleGwVCB9epyyfkhotyQiUa
brJKVWDa1mmnA3tSYW6IxacVoVcIVnN8LUmrTQW7o8RnZbsA5NQ4xpd/UlNYMP7UtyBdLAfr4zJI
5U+4FxGQne9Swp4UkHmF2mMaucBedy3bgjPBdpXZBDp6nsxEeUQhL/FcDlfOu7/Ukv44r+0S9llv
NMHO41h52K5nk0ErVUUBmF2FFdzV2BmigvDZKgicrqs0GkUerZr+J8d7Lldfsf1AzayX7Fdtrvqy
b7EQqFdiUKinIWVmWGta/qothSZeuHKygr1iIuEx/rJX/6bXsEHOBvI2XQ2CR7/0jYzo+c5opyYY
tKYfN7Vphpjlb3BJihG5jjE0fIHv6upHZxRxOd833DuC6koKGgFvgqBpZBWP2p7BDRdh5PkK7x7B
NuvnHO9ZbbQn3mUFIo6VQhznaIrpihP0aZihRV1gPszWmbNwWS4oO9FIhi8bO2puhQQtDXG1mq7r
rpYlPWTXMBRbKQIRuY9b2+gJcjY+3pF4OCtL9ZzCEZzQuErL4gjVFmmjvVx22e6/3Q0TZ7knFN6w
cV6Q3CNZ7C1dzAv1oPJXcIRoFDEa80ZyPQskaMkygFg2yK12+N0JTMOGqdjOkpTIoHx/biegWegp
dIw1iwVoJOO6ljRSsk3vPEejF919sc9cyCxfAaiTJod8kAjeobkjDngFdr8L2e/qo7bts6jnmoJO
RZvFiUjFNmKPekVPR+iYDmjVhNEiiAX6N7Re77akxwP67nbRZapQQHwkSDy7HZp6MpARIWLyyb40
fLz4CxTfSEW4gCLC+Obqg2ISuCeI4ftgco4demAQGfdcMLuItzNn3JbP3lCaCKiRBLaWMB2uK+bj
5C3U8+HL1En2bpNLtYHMUOZd0stfYk3JCf+u9KXO/RCgC7TCPsMWmOGMY3vY9EB4/QGbvaCxv3a7
BJuMPTCg32mJ0JlQ9BI7CKkZRKTcOmAzDRwO6eAXe5yMO0/zVA5Rr7ChNpt+iJRqYSmo6HGp5CfW
ixxLfRr6P2qDYH2rNnll66wFXIZQxVS8qLp3MhILHvnORL9A6O6h5hYc7lQ9qfI01Lu+LlKIcNld
ne/GLTlVPANKpFnXt4E91EnUxEClEimnLIH9Pw1ux/ht3hLasupYUNJXeoVEQh6vBZ+wpV4G3mQt
S2FrdWU49bsRio4ne6LNhfbR7JGk0Zb0rJiz7Yzt3L6rLu5vblGgdedfvFIB5k+3oVPuvGX7UVAn
VoetVx09335WKIM3nXw/IGpMb4ZXq80UFsedijPAPJ8CDPw7GYk/iCtQyaZ1xVhC0SCMfDZJ8uWz
U6Hf6Z/2T01SZcUudOFI/w5ZJltQPx4mHvtpKzZamCYt3LXNK0akY1HIWI7yM65SBbwx5g/SlsbY
dDAxUDWoYf+aQsAO142GsDlxcB5+60o4bhHd1C0KL0BFYEjBUI004vVpcn4zl3fdpX/fXAwAzn4p
twaY8MM78eXM03Hu55nN0r6LjdU3dKw5e2grYy1lwQABYVfLci0M4s1I8cPfsuoJ1uAuJb3tEGqV
zM6gBWB29YUZaSxVeuAA5RP1dQtidKQDcudQXDV2/M3vTko2Fge5nOoef2x1468H+LcZNqtgFY79
hMUcmMbaQFKmaZjTRPPI+xM/LP/aKCMi6bkukh5JhdhhyRMs0bjffWarNGqKxsh2LlkCJ0uC285c
dJfpCcZrI7uKUqD5xiyy2sXDzEvRcUAYOdTTRrhaTCGcK8Ggw7hXLNEUX9lYaj0oySMiooLFBiga
O2jQy/kK2dtaU171QufIAIljlOPBD1hFKpyjJwX2qofx69RaAR/aKVD6V6HZ1DBraVllyjYQxuxp
IVvsQmVv8XxK5cQTEIDOPkiUwDsJafNfqphQHAgnmoV5+4VUdaQpkZpx0+PgsvJppKQlqhREhxa4
q1+j+/Nb1fwsZpuDpfRXPt+HtiB/m6NnXM/MaJZdxI45mIAz9Nccvq0g35tMr68hDH2E6OdPK3Gh
O4FtC9xcjAi5xY1cjR0wLjBzMnwmZyMuwH1UjnH928r9qNLLhSUBNygGCyptggM2N2ll9hk4Tw0P
SORUcgcVkTvLFyPjAQcTHC/flLETb1cTr25qx5TOe7wxSAPBiY1Otpku5rCNSJQ8lr+QNMrhfEII
5bGnNoqHXGN8lOXomqC8wse+b2PMfbVteCYaeDRa3cbinYpeKjEbKTRA5zsFzcJR5pr/db4Qo1sC
z2TOC+FnL4GrahJtX47KLyGCQum9RzpUnG/DL6p/GOq3YNaLjXdIqbb049407+4e4JO0qmSjC/Lm
Zumzpns58G6G3StgjPvKpvFsJxXjfSjqHF5RVrMJnyD7Apy/p/ARedobdMHGgs5mIuMgrXiB/Uv2
JnM3Wnz9e2pKTJT96mZ8QfUA97ZWPyFfeOlg/ZWBu8fCIm94xEswUh2/riyyeHWkshxox4McCXXi
rmuGujwaXMHeHf/A8A5sBaUbdGoUfHJbX0N7yhr5gtZ5HSRLEeZAfQRVzsX2o7f0yfRkthBqdEfc
LQVauZr1nY5H10Mg6safvCn701fsRRhaBTfAiQxcGWzPmSxByT7sbJRjy+DqjkHc/ylw2cMI7e+I
Y2ANg3H8krBbKoYgaeBZNOcBSKBEqDSY1zFLAlViahJ8vVmA+LdQ/uNPKV+yfso7JzIDjs0Oqqa+
ssG0ET3rd68WjwkA4b7GWBLIWEr3mBL3wMuKD4wyocR3iyI5T9cpFM5LvD//M8ueMpf1f8muirUG
9o6xukWG89LJjU9kl/QTYXP6s+8bNd6g3gsZ17U2eVHK4sFRpIGe/fo6vYmNY8bLrPkXkM9RegR1
GFiEqj18OO5vup1jKdQTy0dHZ0lXHOKpojinl+nymHeyMPUyjGK5bWilSoX0SF8FTrledVBrwL9a
5gP9Olg2aANdIBeMw0KrXCGQvy5r6vQtbuUtfsZu3Ie4K1YuwWwyhvfXCTsZf+xUAaxzYELdDien
AOSd6YKppiiT5L/FwqEr0sVreUUNSLlHxDkDLEfqNJyDwVFVGWQ5B+JGXLZSIQtR1sWTxXbq9v89
CaIWV/V86ZtUmimeZxxh11FWGJawyNkCdm82CcKslbntEqSNXRiwN/BXRzZmrwAh3xspD4ovpvt8
uYv1j8Z3WJsOMJjSn/gymw+vU+24aJoQu5ptHHNDKca+Y72ZLKFqwoYN9d651/RBgK1HyQg8t7Ab
v5PXZs4iTbBaAGNOaONRjpl3ox+DheJ6jHCry980dDzCLtLQGRsq3WNCPkY7D8Tat/LpqokAnfGy
lwH76u2fZmp6JeoCZJzD5sjA5aaRvfWwIaqMGVbjngraQJi2u2mJhxWmV82vLULbZJ8XIOK1VOvb
aanDDT170dt1WbZGgBb83efxp2P87LBtoutNqya1j58VyJC2f6vOdMfbys+Xtm/cPKY/FT9FpgHo
mVJO8TeTsH7oJQ2HlyctNeWqI+BT9kUQAWDziXvG7aEgtPfjllqSxz0yCKv+u0kZiIhCLa5RtyVz
nHnK4wXwGIfQzF5qxZtdVm0IbqEaTM1Hldu7h52HS/vh1ufY6eLpLYZVheCTOpLINfatxPJ+dKv6
c4Wds75QdgMqa6RF9eWoYXS/joen8QhwTEJjIdNu0GDRCMIXbEYYK9d99RX2J6ezRErKndUVJrM1
KiCvotItqsKCeMfOuiZ7kjhP9wnZ53GYmoqFqvfbXOOCt9CawReQlkbXwYZtlTEtFfsilutWtPgh
vXauuxku1VYHIxBKxFXbd0qwxiuuHjmujNjT4ZQoqyjYKaxEWBScatbAFZX+0ymds8HHY9FAo+/x
piRjjgAEIly0uPtj57VlIkmiO9+M5t4sNXBGo7dZR+SL/HdBpbU46ob9yLbaw6U/Cxl8FHKUstlx
wETuuSyUEY7A9RQyXs4HFxei+VU6DBHwkGe4ZkMZVy1VW2u3o/IjSuHTtdChBH1ASEIeOh9FNvh7
ELHnWz08YrGyYYr3NOQ26Y3o5IcwIZ5g14elh5P2FDKnlm5xCFhyHDO+9Xu9w5NmobR8Re9jBu4s
ErTP/Wy1Qk22LUNvGtMchNgypNxkMNrIz45aplMmRYK2bjWaj7y8GB01E7KKdhUOo+k4irTGbUD4
6+q871N33zxV6d80dam4z5H+KbIzHOkJSog/uiVXv3CVxkkP10QmLYm+FX3CjZejCxT8ocST0wEf
9u+2374XZCX7meNK+G9PTzuwCR1JFt5WJUNfjLQNnMFC2osWpRHB8ixTdOS5D4y6VvSQJzNrja43
B7jQYVJw1zNNjAeuMJHUEDNstV7WZcWV22MT/sTegJ3amgi31SH2c3XMzk3RsK5NoM0o1xu6FJXC
qJbPBr08Fvn1xzZitHyBMfg0F5iXBRkCx2H4y0QM5coMjY46ewKqlCIszMJ3HQkKnFfj62RtNJHS
52nwIocF1xyGHYi67q1nDavkWGf4g+/DIFVxxVqBDcE32HRdWIoNnLaK9rHvHhgznb9yiBVD2uiE
i4KwBn9lsGGzZoTg4UiFyfBm002NLyo+GRMAtiaBHKXG79xp4zVipvrxpYFF9DmwOzJwi5uC6R33
Ngu+LxzO/n8e+aT4xYYA/G+qpuyGzwO0w/mYJwMZYrGnynm4JhAwMxDbQ0XPULoQeb5ndtJJwWhs
FmnyUSF+9S1n9fgsrR+ynijl53ylj8AdRJysiFOGO4S/h4oSHLEuz695rNvIuRz4keFaDg7rDqdY
7J3LdtbRVld6knF5XgcEZnX+Wqy0JUPYBpuz8rfgs0D6Q6YtszD0AAD1yTWTko+uotibGzjA564S
aLJPJ4f9FFVanj9J3TkGc1kdLf/J9giYVe44W/9lh3gqb6VJGQEIed155/1Gwg8BapdTraAEPIAF
9oWN8ioHw/kfrDJd/xiLc8vIvKaNDeRQJmN/mMpVluyaxvVkJOXp3Y2mlFdC5iAWpQkf4U4xck9M
oZ57xuxCkYnBfuJB/VDaLRuwpn6Py5+3VM5nPGzTxddMViSUWkaTJNBR0qqCNYlkd1judH1LB33M
+7Kt3li/PHeTSxUGe2RAn9thIKZMzJr8uTIuE0AoG7lOdzUhkL7+cT4Sww7hNCTf7JwsK6R6WHtP
RytD+D8SWITR2zH3wUoeSfU21onw1YMwki+JH03NlQCdpwNdP1olpq3m2w1nkAewgx4Y+qM7G8s8
ggXuPkwmXTdrMwTID9XWfWLIrR5JpHVLNV6i0y9BQEXfVU23xV4WCRpUZ1iM7BGaQIhrOM0SXq4X
a9gSCc3UsUB2WVnMgagzdSq3liQCQQgBWMCLQuvFiUuKQQbcCqx9i8HmZSqxtyMnZuF5rLwEc8fO
jv/W28O7SQkSjiO34Cs4ge7zyj3/z5zRa9pDXqOd+PS1rpmhdcFpsoNYKUyahI22g3g3wUNnt7RN
KeHRVUqTT7KQ/XlaIM9DmQvYSldePBYbWF5hymxbMmrDAIc7SGmbJ/k9qDgJ2lNMgdUntTEL2pK3
5UdT3YIN1pI7Lgjn95KuJWpj/UpZjPc7Ti7moOTN/wKplD5pgK2t2GGkI8Z0Sx8KrTColf+ZUFH3
u1gD964xbg6c4rsOXuxe5lQl/oSkoVH1CTs57vboCSgdJm3XMCQabCpfEJbC2sulZhXPf+iKB2kM
Z20jGbemSbHWhF0AABarxB22CRz3Dk9oReeLox7t4sI+P1HeJMCOypDTZBWHa3biQGG63BGbERNT
Igvl1cV2zNw12QUHyNBDC15f+5ZZa0NiqUNqG9H7yMJVICW8Cpi0fUU3zqEY+r0CcoK6sszkcoCg
ii5XBqsajLekLr9znUUBh/GpdXd+bLD4xBj7nQxZAiD0u67hzqe9SM8a+zMNaUOoBp/LnnguPy8L
B+uMEcsXSWzq9SM1elZzcAWfc3r0zaCg1F+vvW1mWZPNMi1Hc5+LBBQerWNr1jrmZRv0CowcX8ve
C0rYGSw23ZjyauHZU83pY1slhs0I2tbzB4CB6Z3WqQTcRVdT+hFn8G/K/ZcWzbFd7FlP2L+bsAv2
p2lVe/rzdoGRailRO4dPZZPLdY4HLDWbAPBBShfsjFmwZPPWLpQs9VcZtJgcY6pd9VgBz7y9WVMQ
pK7241ixOzu/DGkWDmsC8+NsiNiYLgE0TeTW7Stq3LV6uzOjCCxcHDRkJZOTwjJPrQlJnzNaYTuX
yNhlb/OSSMNN5vRV/jNlrZaZ+naztw2dFGadarkhJ7I4U5xNyDMd/JbBbjHCXfHkooc3V1+pvbSP
qYLumHCjgxmdjQCexNDQL9vMaG0ePZD81v+Lnds9Fc0dtxpd2OUK/IA09rnOcVIE0qg3pwlRwSWp
yFpA0ZZm2qe7YV+9iQlEKKsbz7YtBm9vSy9St+Is6n3uf/rbbW1StCbNR7TyosKgoFcQ08z0Va9V
ZxbaxUshEkqbtOF9cf25mX4f+MAar7CaQym7F59irywE41iRplswT82BJPHAIokqpg/iBJ92Xnt2
cqisC8zqzPDku/z8YRWJ2lUWrxHN6ix7yZwJy4hvJ7NwdVMjppM0O4uU/O6Jgujd0YG1PF5tUI/q
0J3gvp+pjPB8lpqXYE2yIg590oiXpVwUfs5ONfD6aUd5faXjHDGXuUmC8IQgtU51jNaIhB8K/x7z
cv4LLjJyh9GRw2Rg325nfYNjLorNHxwrLTN3lnw2Dn6Ge5vkKr6HFzOfLObcsh/ujRwy/J5AjeyF
59d16BHH6tTyTd7ZexnVt33koCuMwd6pOhleAx+7MBly3ShUIBgzeqWbtrrwZcDttIdsIyCOW4Sf
XwXwgE6Jksu190INgoGcPRKqsu3lqePfC3fV4jeKBL1UwOFnTVeN3wrmXBCHIkEJwyxAl21lQ3Fg
5ALK/8OAMPE+RWDT+V08E3AqgsLm6sKxZ51z4Aoh8AkYAJD+bFW2qtXOlDuTArougtVXQRRwYjsw
wBlwMXHYi3rz62NNvozUvxCftIWko1xZPdK5P1duL+FKV9PjlnF3DQRlwgbX5aWWfW4bpaObeuee
tB8WNFGMqDvgYTuoJNyltdhCIOOo94ud4mbtNp/Z7SM0tW4ud8nzZoTq6Sxfa6HPj/l2KaT4Auqg
+iOtJ/fUhfe10AQEeWqLQFoC0JL9bGaLR1PMJWTcycH5mBTo0w4/6csus+ZPTcevwNSYB1mTuhaL
BqphAllJ+q1TvbJSPMEI/phCgOZ+3xMpahQ6KttDkJoc6/USD3/LVVkLQYzhmWs/RFQCSHKqkYi4
HJfsh+SBcN9t6UrtzXamXIGfr6EpA6o4po4y4woF12MASSd6vTgDLJJY3zKJy/JKIAJOBaOKUbTF
utL3/LidsiZHSqjMW4/oQtVSYFvp94Fm8Y5GGUpa3QVRVDpHzJqN0pH8NsMPsNtK5I43uutvh09z
aJx2jHjktn1wYUTT8qvhr51WBiX1yetbU6sh6tgorK1I0bgc8qx2VBrird6G6iRTxxvt9BzQTiOc
J2BsylrI+TQjBD3G7on3ZmHoLUPpISwAmV0XCahHvJj6zLTh48BO98vScKT5eijOv8IE3Fh1tMuZ
FaqGyHSAVJOMrSpU273hqDYrMzqC+aMQlHxivj6L+CwihDGNtDf5s2OGs+rf+qB7095oUwdWDYk4
VuKT4DoETBHDUIBQvEl9g8iSflhvVBYJEawiDObf4itLHfQQs9re0SuK5bSeRir/bzA7Fq3Klk+M
G633w2u+XQTFS8n/zl6Ln2/rfPC+lcfPziQb/msNYJj/aR7iwrN/Jc5H4vNcOuWCCOGF/1M8XU3E
CAT1x3xk3RWUxomd0e+c+HH3fk32u3xdTwWpuZPPU7jJ7z8P/Bcljjr5nTGYbm7ffMAtGfrdmjUU
0q8j6KeIgk8F0gIjvYou57ZuVn9ER6Vtrj/3aDcQKyBRvzgdOcCfWje6UHJXgwFDe/kKARbgkWHX
2mMlNPOkmdXktrk5T/ey3CV5MWm0TRP3uJjUTwJX7bn5MxOFniYgliVJqkBgXNJzcfpZFAwq9PJ5
zMJM3YGV9SAozjOVSwi586m096JQyIAS9Hb3/kWoGPnkWC+x9ZTth1VN+RW5DB5M1AUyedEZlfGG
7J7/wfR41HJHB6Qr7Mkrhc5TMxmY8sEDATjs/+LzhClfpcpKNIovh7UiFUdl94ZW5x/GBEPvJ679
EWu6TXOSnXYMpl+P6HZ/kLmoPm/ZX/3fnwindmaJsnBmh7QFT+aCTkwzP9VSgZB/b0w5CnK6QbGh
TlcZXTCp4dDRe//B0fUswIVuOKCtG3jezDQfGN7XJaFjREz/if1T+NH567rAnzP5t3IIOyC8PgaA
SCAHHOX+1aoAtLdxOSe0g6B07FZkWooXFdbPJphJNN16u7cHJluGvfuIzf5iWKw7HQbnpN/MP3ka
uGPERCYzA5hXrkQrlOf/JfIrIdPI/EElAPKJdigQEaKDSbXy7yAncnOudndKVxVPqwJhL5kNPbKx
OP9sJgbHC+pwL+S+6YWvr7+npDsf+PpAXnxB6+/Do9EGjv+PkEqfATjCGpJdBXGZzGF/RqmZ+AxZ
9IbvB3nVyr+Pa5lPL2tlbM6zUEqpkebV22c/pwLF/z3t/P3iYtF8GNIf2YdqA+Of+ltDk08sK7gS
GXQ6k/+dlJyAtxxSmHVruBWN1BjiSjE/NThxRCkzJlpjep8Z9wUf+Ubc8qTX/423CXo/Q4JaJORA
IQHO9VhlyFL9SMnsi7Il3QXv0YuLFUO52/jYrUjClwNbpMSdHfxjmHKgCY+DPuLq0RWXDm2xYspn
0vId/oxM2TrsCBoQW+x7DuEdwmpQ64J6Ji6bWygdQvgVi9UFvJmu981EJkPj7Y//n1JPfZQ2x/ic
JwMyHPKyti2EAEaB7oEwtqNHjlHfulgaS9c6sLxJxmKrRjJka4TERmvxX6aJUMhwyU7GwJBk1gNW
vMS1BGAn5zJqHWV+o7NVHgTJKSZMs/e3m9DbtpUpVo5l4CBOuBrQnZ4WSnyxXgsgIbo3GjVgNJKL
x6LBMtW9zyqdVHmDA5Q3uCVW+v6fU6AXsgMLX6+nKHpZBSPnmAAZY2G3HDauqPQ6a+upKZxiDnPB
BeRF8KeJ7Lb0LSDEWphMcPKbqBcGNU1YNDjq0B73CPi+7mRho5BxrbdzwSUGmCdZ4MqsQXYcW3Kx
zuoUniS8XU2pYKgtq4pZdMTWxIme/3EeO41OMLfJmZmH1hWKAxAPev83YbTKIMQq17plkPd3XdcG
GLKScyGdR/s9p7ZEPAZFwuIBLnxVsKH4GYeHO7+8qgbnnUVAGYk6jw65b110C0wL7FTI7ZpkURPi
4Th+dtgg5LFFQ8HL7j5Cd83NM/55UIXSMSXGfHGcXXcylL8kjrMchJ9ndVUg+LaG3gZ6MTSjMl/X
cOGcFt+sflWSvOnBrdT96q8Qyg+L9rXpE22hd5PpKESmI+HgkX8LtBPBepYhCQbB8akc7mKIRA46
7vaegHq0XR01XZiuR8DBASMhIQa3qvevgE4LbXj8ItokO9fNWZhS0sL8I/yK5AfTip/QAId9E+uL
Q7eHLh/v+rh1jissCxPSDmaxLjR2gaKaqd79SVii/uKraCVpLYVOTJBdd8wDuho1XdiqNqW5GdIf
DhPTiXJOQAi0728mW0rSC4nyFw7tyCb73vrjdH5/FFYh3+vnDvcbq1z4qjlcUYn5RxKsOEIVQSdH
pGzNB03rk6U/xqE3/nf3+7WSQdwkiWjubIS1ewcSEKZ2HbIA4itayI8LpoLkj6JJAwgmyLLtr1y4
/0fRolFIWUTrsUJZM3r3D7QRAj0Crwluqcz6msRXMh5ehSvjPuv5kEjgqMJquJ+z2nUVDIqx3os5
PhubLTygRPVyCbSMhA39jdwPE1cPq8/xjcfOL79WHQJ4hohHQcBAS/2jM979HIFzguL8g0kQDEeM
TOEzVzEkn0OfrdBetpdxPyE8egelCosuvvDNh4M2tY5kPKCLP2If7SI40i7bAvRfjwc9M3ZikzYW
0kMHR6GeWiuWptpAobIw4skZnS4Bf9vO1AeUNpdkMNmK+4ArKyFUAtOf77gpcKiKGzOo/iM4DwkG
WrURj5Q6vTs7zZWeTDqHuw/gO8ApzdI2V1Cy6gXAcLc+sIeHD4quMCpPDF9d7UorzfFlbvSsRqLe
V9PDETpfSne4uTPJVP/003OyWxtxf6IUpkw/XD2TSF4gQcVG+NKA+GCyDWuJasvgd33KOMj6yezR
JTEGjODW505IKa/m/IXm0cdlmpghBmlyfDXqsbZXOKntmUoh7X9f+aw+zanF8wJJTRqfc9oZVrYM
Du7Uuv+LXrTBTky8QwcnLwTOUOb1IFEbWhGK6mP+wFdcis5/WXjuS/ffjcaSKMgl9aeLHFLJdF9K
+iqMp55Aq+VYWli+PNYLIo11swsNj513CSg4+sa/SfTuq6DAmLRDlOmLDEuHkZHOOvEJlepOSK6Z
6UDpK7asWylUZLJHHC1+pgZW5aZPL0yhuxjdDC1xOm50mkzRXZ8AjAfIPvuOd382XCDvAR1Zm7Nb
2uP8PDZ0klMozHxqAlS2kstHh0JBPnW6OTPwnIlAo5Zd2b7AMKKSF7AupcMGAPF+bJz3+Wx6DFLw
QnSQTAp5fQQ80k6K6fvzuzrIWXIYR8BqUyDFPjelx5mtWY2Qcj+DSW5qp7CEgLLyWqbD40O0DAZq
KQ+J5f4YdhmtOz+tNf8L7F6B5alJPpgh4z26nE2tmvdHkoI5Pf+0jXXdbIMtsbk2ovBwlu/hMyeH
pANGBHwI+IzbZ2LfHaIbQ2XtCsbCwVS4y2gCbmpsPLRzguUczgk0CKfAvELiNHYKI11r6xWrtLtQ
K5mVvUE8G4hr0Y8Zdn/VOEz7KBXfJsgRt7y/Om2vENDYNRH83OjuAfb6mRcPvHUYWjx4HxK4ezpl
F+1vXyHSs+GjSPqXj2fzHnZDzFGyMB385oEkv0n49u995V2U31lMsvN4vwBLbIofyq/Q07qEkFG+
yrT8dJffi5VyfVyMuFqbIUArf3lGHvI5SgPbxbdWYAH6GmDSBGCPzzSZen/ElW6aVfC8G9tjwxKg
HYI1nfJG0+OK/B3j2Di59/P9W6Gj1YHNY/W10J9AxiBdos2kWng+Lq23pnL1rVIU+3Gs1vtz8/dt
faYm/3xiSYejpCN8J15p+2h5nuDW6HRVBQSF8M8TGpYZMdOLfwvzCmlhbhPTbK17vhCmGlvJTMbv
0MWnw1VN6RzOeCD1HN6NvIvEysB28yKJUQEwjtltq0WlAii4gc8ykQYb4jB+Zs7Gqx3bLAOv+xJs
bD9VsQ5+kD6kVU7iEyTPkPStFXc5iz9g5KJ+yuWpqncGpU+I4eyeMIQs0GkawESyQ2R/RRamL/5N
rWmpM8b9iv5bvigEXxWNyU5oGpbSbYexGroWxry2XbXOEmpWxg4Cj6I99biPZhG3y94F5dgvaWtr
V+AQr0vu1+L+MJVgRsQ0xb460DClfEiPXvQcDevW5DSUQYFB+dMMvzAaXgMGcBajUeRxtwW3FTV3
MfgnXGBQFMMCDRH8WY6YwvANdL34T+wL0nuMEBaUiM8uoQ74kkeolHrezSyq+WYPJ2rbi1iWocet
isLMymjIq9bU4hG4ZIOo6OYrnFoOD8yevB/YUrEDcVZaItA4sD0SJiBPHnW40RwoH2hJCNUs7JWE
UvyJlkm6z1u/SdsYj3vTrBmVYMCv97tk0TKbeGeVaG5pV8LoZZcW4qn8S2e+dy+uN+Lagh36AVBl
QBG59htLgGDxh38le+eW2Z3TXi8pZL8NGvnQue70o7es80PwSr2CDqCdmdAnNhSm5k8ZqcAJmTOp
eIZtgdnHVGn8vUsfU2agFaOEr6701Z5DaEF54aLAwH7gnUjnJrq0QxU95UrK4SKI9WcbmtpjpDME
Fe1TIFYjW7cVjCEQmPpat/fgPNzRJ5YteyZge6Zn6LYVfycPQCqs1PnEh+257RzJ6YfnsS1RO5kT
4lx6ZKFHJfDjyrYb/OEFEIWml361WPnVhwvoLsoOgzoqkymVfvuOxB7ZZwa8JZyYJMnepkd2Mfly
1HZhwaoS8qixb2BhlyEu9QU8/CEzGpJex+1AKHFzUn8P+6QM5kwH6XgXHugvakEFFbisTtmfbD2v
XSWg2YpwKeV0O12qbjw5raQZJjLNpZ0lUPTYElJRtx+m7HtCOXqM7l45kI/ZQFzwjhpTjT2DVG/X
ztOb9ZWNF7Cxd0h90alWaews65kOxZjjeqox/tCYHkNwu5q2MGP/RSi6yhlOE7T4g5HLCbn+Vzvp
yceKHAGYq3q+ANbN1JofuzLaOFPnkyczrN2I2NG72DbkvOs+u9kGdA64gRzuzXZu+t/pi553iFPK
3CyjXeodtxM2qFG86uk82GIHKKJopDDkr4DG+XYDi7UsahvlPwqz7S1vTM0hUQa26QHeiPtYpqB/
xHoylsLBOCpeZLgZbu/+47TnPMWh9qmxE/7U6Bf3KJyd4FBSiZnkCJcwZwwd7zUcZ+ZrhpvOtOpR
Jyayqp69obbSgMOODbbHt0ewX9nhgkBqi5VTxZ6GnRr1vkaLRHpvNdQDEVspFIpttTo2oP/Gc3vW
jyoNlq9X/1V8Uk3/GPz0RpOwNf1yeh3tMxFYk4/lTk3Q78IEGQMxPufKG8hWE1siiV9q8opsTVHE
sO+q+fENPOsdHzBiC6XRmK+r1yjGpe1JC6dV8794GQz0OWsHeDg91cwS7F7phEqp0UOXli4ViycF
+DtUeWIjizMcbuDCSMvXKDIBFJ+YIZ2iYL8VC4SaaAiCzxaliY4nnKfodwKyQ4S68K0x8rvctIJS
13kQFvDBhwRWXF87CTgUEqkQktGjGilz2gK3/6DM6AFIYk0FUlvuGbEpo3HxGBWVWve276wvyrmP
F0Lg2aIQpp3+KkrJXRQlQ2D0ceAlwb5rIXGHMPoEqUa8niewKk2jdCV3gTF22fpFp5Wbi1dw9oSP
1wGWeEStuDVxccN7aMCJJYR4FfecRouZbLi2S2+vwbxy2Ai+BfO4LPF1YKpwdKmhJER2SHKSvb8O
6S3qMC8Qp6rVpFYnB1GaE43XzIspiJ+kBVCb0aPyazk8sqBiKFadrbaxPg+O87PA80E3MWHWFQUd
3+RiHSLR3aRq2JRji3gPUVHpJlnL2AGqKlfwY+HbayCUg5TFl+rx2hhU76M+5wtMYyRCAIJgsXux
mHYBFAxqEzFUi6LgjO9f2V1CQsenLWH6VDIceAgbbQZmctkcKw0XcMuKuA+1T7yKPuYMtxJstVLr
lawlY0SIkMItBVFWgALe3nNH6Wu3HvPPvHigg9vrnC6+MxKVRMSV/4U44E1fd1DvSQB4TtTkSiXb
zvmIBRfoSFgV9JfgJl6mvqRNDoiBYkgWWrwA31so2Op+OBFk7jpaOEC8qY5YB6mIA+F8gU/i/rBJ
OlUd9D8b+Wkp7n9y+eHLj0oFyhGNC0pPka7TITnNh5TfQvAQNX6+tJ9FDuzyE96HTzEs93MgmevB
AsmZ6fYkw9P5kQtA7R6FF9a0dALfOCaE23OvMR3RR7qLdSDx/9bxf1s1rW785e1lQjHdujobqjfh
hT9Q/a2sNwGDqnxiu/zmHtjrQKnJgU8veyT8ANa112G5YEn/fKHzk6Vc1aRt3y+ENgeQRaraMe7g
dO3qmBrvjlOmvudizdoGEXTpBNfk8PQU6FbInlDcFF/nVLCEYXDjKU70Lalgkbe5QrdWRO1kP+Fb
NTQ//KAdkswV4dTMy39ncBpswxrA/kYwCShHb4mBOi7XPFTfHlrpUmdk3ZuQ65TcdOivyanHdeR1
JAf5ORfpt1vPvuhIYtKurCeZPZhbUwAnZT0xjJs2KmMOm8WMR/DEaKoWUTYrqG2OA0MCHqs0Ru1i
75M5ImjrLGAjVDEs1yp3U34YeTBTrTP+iiRUEksF2MzVS5W490SK6I+RNjf8M5M8nkkT2alqmrXq
odiUb9Fzdp0LZ/kpCt9g+o21lJ4n2/jGUYR9Kkte5wo30exKFXhqLPZahafZNi54jdIwq7Oos/Vc
VLpWf1ACDabu2XwarXuX9kV0KJGJ6sVhrOaqgPyuI+eDkYFQN/ajs9gMWWqOmrTy+d8l2w6G+5lz
pZu0eT82u7cSrTDXj+GTbitQ99gnBM0sEGx6o6f+1eUAedpiyZG/RZSXKS1Rx9dGv4pn/LJwboWj
qrdpW2vschTDGrjzZeHdat/Fxx8KBKe7TQpicchw7gHgIwyD/Ong4Sl+uErEAMHRaXrM5gRLOFxu
NpqyPTkrHtvTmMXXghbjUpbPfOV2zHQnMfJI5GKpTX9swhOPAQq70z9KHIWE/JkCp69/1+We7ZXn
O+mMuMmlvjMlodoFHT3skNm5DZ/MW0zSH56qd9N4XiImIPlBBepRGrdImtCJWtk2gTlPC47NFJeI
MKoGiD+CdyAeGKVifRxArh/BjXV+pw6GrA+RMWtRk6v0et3jU1Jq8Qw7NyacTBSP22I5CgKml+9G
omoyADirMiIw/jQZkwU0FGrrbD1zzqbzbXwSPtcTVkO4KpnrXLCAoDETP5hDxBJwGvudzrj2Xvmv
mg6qVaTHA06hRq8EVxtvB/N7EZrqtnAsTsYMWTEYlBzuxyvsaG6IqwkeXhRifs6D3KfEAtvJ1tPa
zyxqCMel/7Qj5sUSIddpFu0MkiMCBfNeCisuRd346UrFvv7ec/DF5eJQEIFef42DQDGJPgx1hIw4
k6mR6RJ+yrRqQUtg6S/XrBRJulS+w8xLXztWOCXaZHIQwqGzyMIQoXQmvjrx35NoQXjaWleJsxFj
d1mB0HR7t8pxepnf2HHwcBlF3vEL84KQdmoX9UycqITQ8R1VKtB9k+BhUF9NwT9a9MtEQd/UXmRO
uLUPqZapWHHbbEHXZCV8RHlzr2jW353MtVal+xd48AfOxa6foQ79iIKKXdMOK+IV943Gvuonygb7
+lCrcPN9QLkzrB38D7QfU5M089gpQ0Fri2ZiigNXpRYwrUM8SFLjJyAfw4oIf9C5xd2Rg8gL7p0I
d7Je/pJMOUftHEK0jvedPFznGeoLZ0ZnR6DNexwEFZ6MP5+Uuua7Zrf/GMe214Ww5MIrKhgj+Bf7
96JMG6d5PRyozQk53nDR67KNoczBaYzzBTnDmiGyOf408SKBCf0P97Ga7s7HlotRNsCfgSd4b3Lb
beWUP7t4A720KRP96KvhB2f6/YABvKvSF5iHsqgYsL5vkM+i7ObNS70eHDuOzKOVJqKG2VeQhaR9
tZ8lnzM0qw5HmZueNddpcN28CwJ20Jgg/zhUz/c4Bg/uqDjyc4miFkdkHeLElQuV4UbSZN/bztvB
LRKnwBHgR0iFctEQupobZPUPgByv/KawiaE307dlzjzV2kOfR0NaBHX5ymJiwIiVyr7dUQaXDKSr
QPPdsRl/NWk5Vse2P3sJ/Gkml6dA0pvBEt/sWCWeChZUk25hJFP5/tgm0USvqL+6g2WaOam9udvU
NtORUL7/11yK7fFgOlFQ4/erUxhtauIcFKYMYEu7KfaaS4Z0mBuyLKoqyuRrQLU+2CS2MK58Z/h3
Lb/nneLUsY/mHiobcOdx3x7VSFKTpcPIVQ57mTCVitl0tWjWL+hjbbic0MUKO68VoZ8L09/p7jEa
X7xsXdQmHX3flkd/ET8DHq5eO/BpHqyi1Y4HMgvXD/Xij8lo8+CzhYU8wGdQbuFUQ7Q1+L9oiBwd
CzBPfbkTwBt77FJWV0mrOHTsTmRb3zQXFkd+K1bD32ZVQ4JrnIGsDw92LNkkzTjGGxOfclOGeipS
rXucAhA3q2b2HfMQc62vSHkqRpNWhLOgrLRUIFBg9n2IYa0v5gr7jWgA2/vSjxdjOyxlPAM3pbsL
Fq5k7xhvgLF5Clls7eFps/V18ajmn2bGlgrJVZQqkw2H+C8XPIHd0zBI7IhnGG1WEFodp/WBD9dG
wTA4NlQ6cs/IC5OPNkshpjRwM2x7XE3tDHbYwstBwkPC7riHCMeeujq9+zZu3UT1mtOzEmGTxoAX
qdaq3MWzpuJm2GjYJxkbXYNfwXDFuBaRvjbj3OW8W6wdkr16yGMatEsKkrbUQ2RpfXlJ+PsflyOL
RFVFodBPU2d+tn/Hc2KzKO4KQvhjJfqyK+7wDuixc/49+LeTM0dxZ8YCukDlF9SS4t704hozztOC
oHeqVH64Z2ZswuaGeNleSCGm1psCjTGkvYiuw43ihdf/wzVz6VkFYD8hzCEmnZN/Mc4W1O2+6Dbj
IIlA6vFCNH0ohmD+358JD2Q8097ysjCHJt/8RbC2h0XRlaGg0j2XRAQZR4fcToy5Jd1rPK1Bhzi5
h0fNRt0y3Jt3rQvfAfR9yMwj7MQBKzyy8csM68Os53QwpX9tuQamd4i5kWnzOgtBwgnaqCpvI96D
u/2WHYRiv0W/oRz9otissBVAXlLDW5+t4Irihms2Qx575ctaCTezc59JJas4uefy1Yd0XG7BxSta
CKtJCPkGuACWHInLINt81q0vBttBNt6MjTjruxUHDw2VdvOTFPhHMtxOxji7oKQoMfKtMztzdURs
A6babduZAGNCwSgEGKs7YvT5KtqgroB7G1aEpjJzSXz6yPGvAQgwXiiDYsGTxF8RKVi0JVDUAAw1
+SZnBfwygopE4GLbxorUqEAobuitg3Zm9lDa4ynLaqpJB3jELlDVuIEGKKDwcXTbhzJ5J4/mDDya
MSr1ZDm60DtupTZg54XU6sq1maxB8cablxhaOOU+9nqhNjqFPcIeyxsMh6YaNKP4hbcINIwcp4Rf
jR1U8v/TppR2b6pjG1JY4Qul/46ZSojIV8Thu2uwu+HiZuq+Re/2mQIMwEFjZJ2nlS0Nxe+8c5o5
3Hh0g0nTiWMdpiWUd/bn7Dflng/ioSQABM/TLNzAM7Z5BHkHPQNZoWR9qqfe2wZsuqxZmv/e2xCq
Cox9d1Afqa41Anr1l3hslwfTA+cVdEpLzxtIORZDaBii9U7JTV/07++95ryjt0S5E8uFSxxZaMt8
E+dPqER6/uJ/aahviAOIl4BOH4fs26EoMnMjW+Uc8KmZbfli7wbdk2/Or8el9UKpxAj/RyumXST1
7UDNRoH/miH6H2Entas2ZUI/aj0Mk8T8eJugfj8WredLMNRh+6HicwmE78pzlhst12y2UOTvExlv
E7++3x3sh/i/7a9xuD8wKUW4E0m0z9T2A+AerWGc2ot2GIKBZHnn8EHh88pCXLaGQYcpC0HtIs08
vsBf7b5RiuNjhtcfZ7rHCNtr+5dDp0Sbj1DAZQv5yVZqn86eG0lj5e4QzEaZpQE0lWkVioQZ5grb
8njpueAGPeViIPtEgvHAjVImpzS2H2+qEOi89nNIm3+H/XKF8R+XZUgi07RwVPB+0K6sWFp4jq8/
udOkyVCIT4epxKKEjcKu2Ki9nA0KQP/rSOV6liFLllpDD0SohY4BvdTsjamwFGuqnm9b6xaStzvh
xt3AhqgWcGRtswr8eD3b9MHaXO4iorncB+XuDAWqv1cmBwcj0IwKZtZCQIyClU5PrnYWKpe4tRqg
jpuLnyWEoLzo8ZUu7i+50PvbpdKEb3LEBrb5dGHKchFLIEqyomnRy32c0YwVPS5RcyS6zUDiOQGl
PFu5GcTf3EKBwBFjcsLRMNgGOqXh9fQffLJKMCUUULkOWqITZKzwVHvC3Frs6jtCjciVJDhz8ZUw
N0tcpWbzUffI9oID18i84UlXzG8MQ02saSadi02u2D5qPkpAbHYR5OYFdJR+9N+x+4Cwpg+x7FGk
jUx95WZmk9FmHevfgQFEDTr6+xnxUT1JXkT7rlXi3gVRoLdQY9sYf0V8BweTC+8oxdErLoaEar4Y
7ZzHKTRuyqJoZ0494Z4+Mvrc8otR811gUlp+y1ejNdZhYxlKPa7Czxa3T4PNwD+2cZoUnIbQXmgG
kPDYaWlrGT2oYcvbTE1pKV8TlVXweBQC9fkystnOoVc1tLIj4Il9dRxcWpJDMzijM5mHLqtateUV
KbyFvoLpLNNF2rXLtr+xS3B/qkRzAf3g+e7MoeGjnMcwmNrR0oLHQ5ODV5t/BbRMUalPb/W93TAf
a73KIO0BQUVxdlrfAWSpV+m48i62RtsX07f9mzPLxf25SmUVUrtrGiHrjXoLLJc+xUaZdpCNLbLy
KF2B9BkBnC4TR/QTmEN+ayypUVpO8qX39NtUUr3HVdh1qIqu8j6EeXv7obj6jO2NKZtodvR5c2dR
AulYVAnxJsZRgBylTLOCzjKpsvf1VNUBiu0rDACPPIMVPvVRP3GONICeHR7JqTlQM06gvtRGA9tm
1Q01nCAJh8J2RtnJR3WeOu9Lc3Epk/HiKRHMbV9yXw8+h/N0wJWXIdOKaTWMRYpLuEiIe0KyjrsK
PvNH82POstc5hhP7fPlY9nNFpkzybhEbBS/y26Mb1VfyGgIMcjz0NfB8w/XVX22yAj861XVaKLPT
Q8xfEaZjglz/9ZnNw7/wq+XQia8Witg8S47y2ZILs13mN6kjLSJUNogr1WUodNZVtyTv5xefKxPw
MJhDDEtPEn5X7XC/x/uHKkJjAi2cSK7FJIt3eaQjeFK44R116k8JVHnRgUGErSdVdGv5v485kGFr
OcswRDiVsZBwhMjHb1+BXicd4x7GCh4stkT/sdkW4FKaRE5bL4/OHFBqRFyuPqTRnatgjhRaDz1H
5OBOgwPPdEXZh7jgmOHIx5+lyKBzA/CHnx5GulJGFuI4vKyRZY6+aTpTt+1J9kyeXQLH4+yjEB/t
d6OsHuZj8156aUSq6x5wXcaf7iXr+fbo+BMC6jB6KwZ32F/56aS0m7LaxUl2Pjm+eZwN75v713C9
F/OZnNuNtPn4IaXjMR4a/AvRpOXSrlSd4CrvSia9dCbSDDFgUYHgwb6LC51pSzdJm/jhZBTrjIWE
eIg6KJETqp5TVVaUDNFl/HK9N4V+TbzVOtilULrAaXa9umhx7TMQU87GU4ADWyuxiokM0txJrNRn
L5d9UFaLHiGpUcLRhge9I2RQc4sL7lD3qsmJjNzxBA2pMpPs02ljm6H7jDkqEabNwn4RI5Bmo23N
DT2B8247lcBOTmjY6l8o8Bo3qox1WPZ0L4YzpoDI2jbm+YywtEDvV4aBeJbFDvnk9Q4kF9lW1/LH
H9WSHa7YcF9FtvjL2Sv1ZKNNpzpaJGD7SLn7J2mRdJxpaQgYOGG7ht/ScOdbsW9lB6GULcERGqTn
R4qqSojipFkjXE4CblPHWqXgzt7zWv0C4FD9yL2TFHfexwhxO093SYDX2BN3Hfcst+BA9U3p3P/z
xUOViKugEg0TNvCYXnd0vfbom11+ylCwtWrqPUjAhSNoJJ7HWw2rHjaEJidFuqKwHW7dUOOxtHiq
hnIy3FXzNbsbXW0jndVL+uAl35xU8tY5Xg4c2kJCTJgYrcVzKzcIqSIAu1iliNR3UAOH2g/eXnts
9Go74L6kTgkrfUavSUuq2K3Nw+RX/8Vj4v9B9bxWu2z62+iKoZo6ITtpGgSrraEAAXuPffWcfkMe
05Hgyf+uJ7j3iSz6iRj2AeR8USmi4GhnYvwZ6KzSscTbYPnHYZyp26ZzewII4/CDbPwbRyDa9xsp
btbud6/iguT6n9Y98gm4gqunhrUogo/J1Us9u42VXNON/oi1rV82Z5jTTZTPtx52G0a8sQi9lDs/
CaxruptEjruTR+OC4Pcrv1fKHdCq99InQjpfNMI//nFSpAieFG4XEBMBO5Sushrfa2kfvd6ySc87
4qatAXwP7lxmaWxlmiqxBhj0F1lxalN95oL8oX76EYLKLUQ/TNVZhbJp7H5tnZOp8rd8I/VQqn4R
SG4mYKbB+gJ2wggUENUneZxRO8YY46s6i+BQK/IrnK6th3UXclNDPF0kAjGrxewBx3/t/DjCCp/W
cczoQ5fzKFLrnzWZ5+UW4x6Ysj9No/LiEOY0nZVwksZmKHH4YIio1Q/C34Zh8RsbdI7j9iRueuiE
RwvZlmoBPvEQCJQSFpYzAawskWSchp1IA3hDoF3t294f6YjbBO4NtZCnLs9Lg4w0kbASld7/Y5gU
5iDHGOpPQgavBeiLucJ4/02BU6O3bSey2MgfLC5TzFW46SaOpYS3TkwlayOnJGZ01vwt9hlfLCbP
0hhsqz20cIBQNe5eGA4o+aTUAjPmXDYzaCmlfBgP7RDxvO6rVvwXodJThOthO+YhxjdHK8QjLWaL
ppKrTdxhZzkBee3ICMBtTmHJBtq2sB3So2L103M1KZtmmsiQZOHoZP310Py/f2ygqrx3fxZ6ThTo
a89JkcVbylKn03ifN0nR18RwB8WKACnMFECfKkmkX6+j6fJty1RDNazxcvdayrhuJCZh07kVYzWL
QpWmR2CufoqjudcZCwi681sX7NXWawqkAxN8Fi4fUhLGno6Hsl84cuH6MBcDUsdCTdN2UecmHm80
Xu4yKPS1PwsxDwnN2iiCIv/gdAg216I8TIiBJ8eHRbqYo/rNYByRYyxhjbYrDoT4Oa7sPPB+Ieus
GkcXOlMVCMlXNgjshbIaJuDed0IMqpSrjtwxwEsGVaLYWdc5PBeMzx7CB4HQoQWL3jNpb4OinzXf
WssIqxkC/Uxv0GXQzW05xhMheY/MZdSTmm3/4dngeOBMPA327gOTObP0jeYl2qQn+gzH6WJORJpb
XVtwQJpdZvuP7vkdK0/EB6D3ZiNrBSaFdAzeLmTOHQgcVUx0ggFd1d9VIqnJCytfiEi4ywHqY4e8
joLokN8tz/QEvongdISPjq4Ee0+ikWPUEWMr94A0mdawwoKqw7awR0Shpn560yEYauwbgapo8MvJ
9DXfbVEWE+OEyM4GpBg7ogAn6sGsL3BGOZ2103/qXxCpImsN6GbqfXSdIAHiJWY66AHFW99qcGrV
Da0w7HnfkW5tXjn8FEMt9L0C2GmRiCaPQnT2ndhUDGkRvDlytt5BCwnLpUw8Ax6znPvTii/Oruyp
7ofqMAxtau/+9Yp+0F3BUbxImlbrkDDroK8/VLheZfQGN593fTvDWxp+mUS1g4mv1ge9Y2dNVyB8
ujAR/MoqhIzC0kIFg6O+EHp43l0VBdgVYgsfKSGOw/yaVmugZMz1YqEAAv8h0Qt11GeepfEIhiY6
nQ0xcgwdzgo0EKS3B1goh6dyeuv5+SDJ2uZ8JsE+V6V3sroOjpMZWqZz1uL+Fik2J74HMRGO6eYh
VlMLl81Liqa4aRLWOggkgEUfCWFHAgyNTfFveA/vZMUfvB/aJkL+wk5c84TEnO8PXAY0FDE1uqPr
2xsFsm0p7c6gesRuC8KmbV2IA+krNvGGFc8hMUqyPdVKkP1vYpOL6h63QwOLZSLm+RaW2Out3NVX
M3/GLppH79LXKgSvtqbLtkJIsmSJBPrB4KjCKhkVruVDmpXfATgHIxvWYZVWYnjNwhRQErj6SvJ7
Ws/RbbreBR6i+ClTcQHbMgaTxlSrnjCpjPuR4svv1+fpY5tIEN9R2jJpeDHPxQKrRAEWaGGuarh6
uzD2htZPsgte71QhI3TZknKfS7CmXFK6OdRwRvYsULBkP629HoTlYVjmr5osmkBtZyQ/dLD337u0
adlz/D1TqJRpx0adqrUvHtaaShMkpaUjre6sQSs7rQzaLmfwjFPeyDBHd604qOVMdvRP93NfJ1IB
CtvdlrswAX2hEsKFRwvYLAolFjkpUSiaDFiRj0acHj8uRwjHE5mMAOr3h7wLeMbLjMVrp+37DDBc
bdHVKqK4CKzeGsMa4sFU69ANcXze728s8ytViN3az3dy9c+/hRh/RdTvsls9w3fuLwgX6e4hGBZL
plsXkI6HWy3HVICuVJ8GfI5OUNnRyuw94KRbGLantD9PvkQKsv7vZpYkPzWcCdD1DEhE7SNp2XYi
Q+WWh8B3WAv8NlrOXkTgNJQgqfbhUR19ImvaUkO3kxICHw1TcMrvkT/JmNO6X5UMplbam7LGonpE
OvWsRUDGSw0hwrvS7yYrpjhKkHJaZaroltFAY7Zh31hdO8eZWdZqi9g8v0Xh22rZhPJ7nBQKACir
5sqdK6ijD0xdgXcbxjNgPD+7vjPvDToN/nMKimKRVD5ye9hXSEYinNsIktGwOulk4yYtheraR6uZ
lG6dbvP4A3vrbICaSEkavAx5o8ZED2kdMeN2sJI7Pngmbm4iD4vNkc2lgtaOb5OartGpmp9h3jFP
uqqS5xcnWc2vVTHrzmzqh8tCZnhV/OLyIPXjU1EpBfhRTqEEuZsaYZSQehHc7Ps3d/QVSsXdrvmT
CmVpDflGhXfZrJtSmacPUiqrxnTBpEDyDudm6EktxX3JziXCx+zPTzLFdekHrUPNv2mDAAH1yo2c
D+L+m6esgf8RwZbf6Vsj4avc00mdypSz8Kb2VoaFFl/d2o4szWK4Hd0MgPArJSeiCobvmMT+S4Wd
bPQWeIRyayNO+s9y1k3YuSXpfxbxfRh3mfHKU+2MyciEwu1+emSo+BxV9gWe29TXJdeXcVDwcHX4
QcGEVd75HJV/uSx8R0Gb273bcVUsGJAQuY3nDlhy2mtKhiBOjhA+C2ueMq1mYjwr1AjvA83gy5tj
5640jMbDbM+K9Fev2c8UCI+CNMB+qre4qsYE6zpz3IHY/BP2hgewvsG3hWXW6uOr+zMXCIM5TmPu
LNGp0roJO1A7Dwrx4bnxbndTp6wvqXEwhtxaM50Kh6W9edlA++/sgnimGOHJEm+WQ2U98wgjEBKT
Bb/LFgqi9HkcVhjrjtPfhZ4MF5BSYD+zK7+T1SgxzY5Mw0uqWKuw6sNsBCydJvtuyplGrfvInAr/
DwaCY/P/ofFX3lm3jirC7WtNY9ikyLXEhxbdJPgt7Ruvi4ZU8NPOtJdZvL4x7lRtEkuRCKeSeFQh
LsRPuCXgs7N4bXfro0XTTtrwM9UM1UyzjcW0STyMZwb956Fw0cBnpBFl5Vr4gkoZGxkwQS2EQUo+
OTBolJGRqq1kOiyjyRUJzNdyh7eKjYeqSplL9Vy+9ujtkML7PX6ilfr2akjc73rydT7tLqWXgdV8
Fv0ZRrOh/TL6sh7waYperOmdLDNZ7KW6uc5MOyZMs4XU7Zkcm2pcUToa8qOsAUwUgu23VvRzszXy
ny0NuBr92VZvjh4XU2JQ6wmXABfPSBasmwnLDgXzDpXSPEgxeMB7+YR38t4DGt78Tc/qQuoE+Njz
+qRbceeH5lYdnDrAhqAWik8OF802jjn/p0hXD3VntsfM0OGtbFDGMXcDHumFNH+D516qa8HabuMS
l2IUCXINu9YafMSm6NFm30EVNg9IMPbEgUVdQfsFnK3JAMj7ewYANJdUCO1hPsctC1ENT62y7on3
4dHHBHijHf3Ue7cZfhr/kh45QxP0Nv7xUW76SCzmH2xqE7vMY5cY2qFFi1zA+iyzf3VBJThUA7jr
eOX0P+W755t6ag8vYpB3Xumd12jGMkF8Ecm13njAUeDdSm1vSecCcEHyAa8ZRiwJwM7w25DeDrwF
wcdjimobeFvIrFu/ssIknGrX5C7SFg9ZuzLYYA5qQViuOygbf5ao8CNYqUjVFIfCG8ziJCyJWLIC
ayrrPZZLsSMir0p1dnvLE1MFd8YiUOuzbKnRcU0BoKw1NbLIYJkIeSmjLH0Xu67S5BN9lb7MGctP
rzHyohMb4ztyX7pCv+gyxyFPT7vVNGw40Jf73vI5N21BFFsiisqd/8D7S69Y0sZ/hDcRYdNpC0oV
m0tK3/7pN+0mkjCvFGiwU2njuc0M2mhi9gBuuPyUs0Be+PGcxOAwdsSsN0QJZyvFEF03KhXqQoGY
pgjFXcJFki4q7tuYpiu9e2HbSTQzOXapjDU4H2Wdt7d2Asg2qCq0VsRD3ZLkT4ahdi//A1zKIX8V
lb6EKBTKfCo+51dxNypDjE4krCRYGBNMSS9RBjDcOjYrIKPHA117DGbsHoBcuLUaRfpq6BDqC6dT
H09DNEl6Nf3De9Oa+ve5UQHMUKI88TEYNPj2Zf1a8NSY9TguHfu73g7MX9//NjTaK+5b/pnjr266
611ptl8SzV340+a6Zu1BRd9WfDNlQj9R7bm5BLaaTW3NkZQ/xLWj7/EWYa7AmceRf0aAOdSAWKUi
6y4DQHuEc9YYpC0etysnpPgsfWaBuhwqouEeczM0RgOzZEYcTnLz2HS/A08109xcVTDMJzZPOBh7
Y+cutDfKd4Yj+XLccYv3IcE3zfT8z+GLmNF8Gbdf+tkaHhMSrzNcrn9hxF4OBRNT7DghMkj2/k5f
TwXNZl6uyBqrYjScLiAmvNLhTtfsUEzBFYsLUS0JN4PnyU+916o0AVJ3kxnQpCqnw6+Z2B6Myxg/
xWdovj09s/p+FJ5XVhMSCj8pKsGGCZuyAlYIdkyzPK3bdMmF44VmSb8ZZzfpFnlBUXTBc178R/zI
UFKwcf/ODkAX0KBHUtNCUWSVYRVNyeoKADmTyvQqfFMXWCIw+y6Z4OFHB8MhTeLOjLOYSKrkKVoR
37GC8Wv0Y2jugNBZIIohm2iwsEDpHoF5tE/BJaG1k/qM3X2c68vhUdlK4jaj3ws6wAlwQJ/jHD/F
rgCdbCNV5DRhMZ6ue44/deSeUGxN6eypRUm7J184p3cumlSQcEtVfQAWR4AhIZGNbZdYRYmtCpE+
a3efvZIB13BlqxHU1lqwosUvz/ONumFI22zwZi9j6t7NSEuqlVRGMWyet+yVG8ziVXRde1Zc8/pY
QbhS+qwstR7t5h5bHlduBNB5Jw2updyXIFU54EDRV0/Gt3hc94iBYN3k0f+VB672eBb3GWIX7ycS
DLj0MAOIsuvgnOK015/VvRrXbpIMW2UZ/vMhgdpBzSIo8BaYWfvKQ3MOYiBpOcAmF8XXz0TBGt5m
mSXbf49Rm9euwIQtcD0453bmqB4OIP4FRKc2GWzNyfn1OHaDFGNCwg9+ozJrD72ivsrlf94fF/Gg
RFJFoKKYpCNcCuUo1X+jV4BwrNPrXErGB0I3PD90halhwQNDDOfonpPIW2WLh3ovakyBHUWAmrEn
77LoKk9bc7eXGlJK11aC8/EJ7YyB6LJo9CPXnpAaq+xsUZqjMiZDeGkOy22FuCmIoCqxK81qicgH
WoBZcW2ANL/VDu2Hv9qYGHWT3hIneSIpV6M2VKN0vdm0vOAPe4Pg2oYMfGVDhW+mSPjq2gKd9S5c
bHvIpUs4RheBbVYAYmAu6xFmFwUQD//FpeSTBNTwbGME8D0rQDK/mtJaRcs1Q1fYFpRNay43bMM8
l9t0hslvgrc+fNuAwh5OY8NgTcw1BRhw0eiXHpEu8F3X7BTNJSgauRFNN5yrt2rq4NUAaVUqdi2l
5PnYNUk5jhn7vo6/k9E12uy4k9829E2sfYxdJJPYNiSuYekjyNLXB7XIxHUHm5TotnA11pJj/+n0
Y4n/mVz8O/SN+EAPmkQFVeCMf6IEAnTzMLXM6EM5iZ667YlfAtC74UHRnHvUbfgQo5yW5vJK8ea9
qJYw7Tkc/4da0KrjqyMU+tPp8KqjzA1Vz80KQfvLUsvgW/uxA6MLXy7YB2fpQiL3DqRpXuzVY/In
kgqEiJRZVcACG8rpJOq9iW34pch4KqHrjp6FShIL2VsKEmzMCvtH0+uEcNytmkgbLm5lIW881/qK
mUxdD5N5G2LO28V9XeasnlK75J8pg/20be/j8izGdj62vvdk02xPkFVs0sO1LnadAtl0tnLrPJf3
BRNgKHHBSFpSDT9Fq6WwWLlpy5OTuXWKJyLGMxuKbEsirTbEP1zxreBYdyLYCi5vd12JT+59o3M2
87BPPMA7FwXHyVyn6Wvv8S+YB51c22J0RqfqpE0J7uXxxfcSLSqcmZlD/aQqaZg/41IZuXbKKFP0
6h88q9c7oBbs3mlZGIDCiyVWp1gWBLNzykMB+njPhgedcidJ3UvCzLfp6n96///tvGYwVCIXzObz
JZCZmu/ygGAjYWGlnwCwuF4bqVl3Ud0kT1/rO6w4XcNZrX+i2u1bZp3GKF7EwPA1ynE4hevHGNbl
ZGFNdGAC8DUqk2t0xKyZTyGFBhhsLa928cu2Um5bZrxDI7CTGmqsAVA3rUSs8xdF82t9yLfOqr+r
m5XstTkvYJbr6XHj95l2eibt96lVagLm7rfooxMy2zFrhDoBSYmCpVw7rOX3gz18wF0fj60rE8lG
HlXst/neulTFZAoFUXB+UVokVoifHdqUegSnWT2RZzVt7JgXz1CPDBXiG7+cJE2WxwYhdGyNPlAy
njC/mBgah0DwQRFebn+Bm4nLzfq0P8VLIoES1bksHk/j8yzEHPdCkqk0JZlMIw+leSlWotD92KEr
IwmyRPdYFCWfq++L48vN9ZhRxvWVshOM6tISYoy2tq5swsClc2tCrWxNvCN+SDuSNbxT6tCIvALU
i+F9JbHMKHpw8JB0nKDe5KiaapeWLmKD3Hby+fWcVlvSzxzmzeRbo3zumQhgV8bf+C2S8wmn+AKR
NugdE5aCNCZN15rIzlzuCnC94WO4mg2+llVUih0vx2GyH9QPfkUDBecxXURVtD2HY/XJrqeeUXnn
6KiY6uZe5yitv0Ykcw54oq4OIxJocO9DqecoAVfp9nclTEAa81JP1RrBDGGbpX4HLnVPG1Dk2WRW
dSsvlwD1+HkEuYg+YlWh20VzxqUbfNl60Pr7Qj4klsdVTkAiOm6AoSIfhNuqsnjzQ+IlgKhTPcei
05H8t1b4zSkN8vr09juO9PM3s5ss9DYlQ+uxiWprRPtCAQYpJ8YfNBt6RpTHSSvQTD5ryx2tE7SR
pFjQp0SI5EBvL2jziPGTBlcQnNkDQBVUuEinfIJDcppA8ecozKI9pHCVunJjDTwBcZj00tmC/SSz
WoEA+D58rYjCZ7WgB0Zkh9bRNR05wfT9P2Pg5X7MLv3FZlSt75LD6buHAWqDcic0VAUjmsEoC8/X
P7+axKggFl4iO5eVn8y5J01Vmums5fot2UO51R9EdjufHpAEBAZhTboc2oomYZwVDrAO/OBUqvlh
SWwR3CCS9kRG30t24VskJA1yIfD72S+BB9JdcFuOd1u7B31QjFes0fpj7FpXyvCQNTGIqTCN8D2p
EZFy5Dwyz11zFqKZc/yAGkoqURT63g8/8kzb00OWgurmDOtzyRLcOvFBRWImWJTfJDUtJ3I80U9T
+wFG3lr0GDd+lC4tUmXiPleyeNpG5hhPX/JZcnf+vG6oG9LuNSMLvAwlDBex44L5NpJ3gqeoGN13
zPLR85fqhr7fehi9mEGpIlOs4VG2KiE/MG5ReHcEYamvwCFP9uoNB/+ydMDxzC2eSY9mhIuQypoU
4HXDE4xv36XXzeLMVTN4BkP/Cgof6hw9lWA0+uka8B6/zJmKBq19PyH01dSMqtNANvnBKyxZiptI
9m1Qdok2WwrltLykWEN6pGsyy8ZnRO0LV/tvdCTHhf4q2nV7qFIRATbacSG775kxo7KJH3/9M6f7
ev1XJyRHXM40rtnUBFgVM/G99lytan15r9+N3/sXmvDdB6A3taVMDKdJ397vR/Q0B8pmjQQ1hd1I
VTuh3tH58XYUP4omwCiifdw7svACBeIpvuD5/TYOd1a2S7ky+wjXcrovdHFyB/WKmsgj/fQxYmxC
bOE+APVc4emXIBcPw2wUoTe92foFyDBDMHNECwRQ7+VQA/fSh9lxD42/o6XnRViLDuWfXGJ4l6X6
jdkBAv0e3SdXUiY/oo5POk5ap04xYUwL77KZlAwVF9kZ2wmCOxrQPF/NdFSQZVR1Ju9new3WR5wp
9wqsdKeqZM9gDsu/nx+fOEBhsMAw+A/FcaYKHMWhFVSdgGG7KZbFgNLURJzkaZ4r5TOIGPR5FDw4
ky91uP9Pix6ba42P0JWmiVU0UvkcjNkgbQW9ldiy1YTemaW9FitDgBMDKwwt3SqLaj2FbctjiLJ1
zernMKE918ARoqZLrhPVe2oe8KzWWgP6P5yA1CEDh4D/UmLrw6qwg0S1vuTDaLmYHJuyODK+WvN5
yZYz+6aKhvXUdOhnf33HYDnTeAZV1WpSjf2BBROUPECBp0aQo9jtxS+3Re5m9Gc2WEGuOa+8D2Xc
sc2lj0wDXamGKQbouzvHxPEKuBzrSd5UqySJtVMKqqTbLsHBQ7tO0PfpYt/oBwCa/DXIi3lM9I20
0AaFalqyk+wArSb/NCem3f+yGCpxdZa8OgwMnwvShBrFgoA+TuE9LA3eDvjvxNeOPaA2cLrcoEyA
NP5z0bYekAVDKKYlcM/qmXOVVj4WTuQ2KHYyfszwpxCHO//KaBcBL1CyPaOOhdza4EbAPL/aoiHX
50wZAoyGQkWQfLGRR1hv8AqMfNFGE4LZsrEzc/sSyckWS0FuQBCSR3nuSSfNcxh+fiCoX/GZQDpc
U8e7LxZZGO9MyXmWvZQ7RgganTgCJPcR6M8Iq+/pZLJ/m+tjxrOET6rZrYvW4H8C29h1q1bWRqir
1VayLzHN8EEJk3TUimG7zUsrXzJDTO2HjUpEUlD2ILwH9C+TkL7GR6pu9EZBhx7195E19phw+99e
h9wnmAukFxXKCxsnypHW+WHMCS89uvOzJHtEIG+QDuWeJMNs3ICkTXXEAG6z3AtKRp039wf+RDL2
TZP6iNnu+JsqlvvHRT5XhUXt4xoZC1I9fRZr2UaV6fn2BVX/yoxmmNjCX9rEHIfvy/ZP2ZiOnQ8W
u01KvJ8dnV9WJreUOLwqwqRBLbkbX6c5bl3rsB+9DhN6vU6ktiN9quGv21Fd2pXllpE5nuKif+vJ
/9Pf375BZ/Tg48IIS/cgkylmqjBYr3g6qH4BzWECWKRdd0jnG8G8tDQsNspzdYvDPXH8Q5e83nNP
GOeulbg+xLwfgHH530XrHHfMRX07YuxKz3ShtAo6MeguQhfFVWLQiTeT9FqmXOkjI3Cri3gh94Rv
jyTxA4cTjBmPJ6wOk4r78hd84uEDrOKvs8dpj6yu+00JOjT7zg6Xd7LsBVDJUBOAy2y0Yec8HAVy
BNsJVwFhU0FJ8kO6apSsifHLN7PM8mX0HYG8tSz8hOt2DbKr1mBKxbOYHItgMeU4jmNPtiDxNiAP
ZMpMqSdDxEiJS73G54XIwNQj8pQkpXr1SkZqIIutFTQHPJukDUrbu4nvtD41zwgybPwTuXlpOa3i
WXriv/EY+KzS7g5VlyomfLzxnW4ONyhzIxAvPl+RW18Qi3sxRdaawoKV1n67AKfY++OjzXsHnYn/
U2p5A4DwZwZrbeW7GoD3SanHym7UWwVqxzhaP37PIBNB7lUyOAgg13aSdGLmQohJMvSAGt/bgmW7
LWh1qKBEX7qq45BI4v0Cc3hsCEogjpLsNqMTBkt+yNWhCJwwpzFbA4Ow0UDrNIZAze0p+3UmLG2Q
Oa51deS5rRmvK/oWk5KQr06LnTd5SOyEqjM3zDuoXwhwOjKDdBjEWHQox502KsMsxZwXJlIZXzeY
acjjulRL3RVEe7RYXJws2JbwNIFRybp2kl7EPKTbVPRR9Kmx0vx4ujg9KMAGpwYmQuatVCjNQitu
bwJ9bkRdjOTryziUjwkTZp/haa+I1fgqNx2dptRPx+GMARZtT5ZaVtDjWWsrSNJrbmrTqbzyvarF
P7AjuEAOlGoqkMYmybSV5ouvABPvs60JNOZ6r/lc7wPyDLWEKhfpTOUAU6MP5bX5zkK3G4zChY7q
rVruqbwOg3YzqN+XWca4IM6mPlPo4/zbHT5LTPKp0pgRgbel4KSWk3+2NvAAZuWDdbNFq2CAXBIY
mathHOER/BxIeGdS3h7MdvzAc/d1N00qk0z9zsgHSnM2bX5MxMfaT08PRta6i60xeupyc7oIUeaH
BZM8Ttp6xhvlholtpmJtDeBsC851i3Xw7ihLK9kC9ujcvMM5hfM37Vfh4Pb3QNb2w1KZiSG47Yix
8fb18DGJrNnYpMOuOqqX+FsmNcuIV933rNx65nQ0jDKaRr6JQa8sb0Jfwq3rVAlHmI2/1HBCU23F
5rW1Qqu4b/47M2NZnZk1xyelgURG5H/zxb9r1aAIs+Yykx8auuNBKdMT9uJsIRQ+oYWwgCHEbfyH
gGqkHZ12mJbdGD2NB6o63sBHf9Q7QZrceR0drXrQBda8QhY6R0LRPQjUSWDVP80FzRhAou/OB5r0
XJj3NAcFGVm7WT4rVQDpgv0rhv5YPksRGHuFXIvzVOqYPC2F3qSYoHckoTY1bVZxuT6SHe2LJC41
bl4HLybgzEfgoAe/TM6JIj2p626NaQvNSEMW01fMJT0NcX2r8SC7XUr8TqgpoYbien5RIGY2KLBR
dcB8CyGqBRAJbdGA2O0e0k40zNKtb1OwplGLwLF8zF+NArvVJFWCCrrlXZ9VPgymvOp2xkZ/2+0Q
u3c2qyVRsfUxz5iw4/kf9rw9gB/Dm/erYNe+sPFi1fJ/MHuPbAoFJujP/UdQSF5kSZzekEperpFF
EfDAwUi2qAeKBNlXKZNGOF+mRYHTJP3tshQrIxIeiPYVvBK+igS9VcnLzpgp1kYqgJuAkmvToPl+
CM5YMm++QI8kTu8XuNqX23TodSofrNBT8mj5KpXRhvy5cdpgQlQ30g52c8yVb+aFRWPV2iwYTfKm
Dum/PhywaLZvNasbC4x+dc/DR/8Urv4UHij/IiGoKUNWY4S0yB9vE1zcG4V0t9EIulSYVcembRzB
QLfs85fEDFdNjPU5X4Cgtn/bRAvNA8TnhBCyKdbLqZ8n0FGBvhlX+DqEtxjeEJUNp3EtPC5NUrM3
VJYTlrZbrviH5ebw08k0X5Xwl1izKJz4jbmOhcgmJtWfJPi9uMahutq53aniAgfVKAGBF0u0+p/S
5kLPb49bf0ueMbgEQD/W0CC3cp7y25lVP8rHWxNkUiJ/Xuroz5RW1bMiuGv+cwPlmrK8idwfgLRP
InTe15PRGouwhYDMOQEWqXOsd0wLswJ6doFJ0lkn+p1jy+zP1nH2S9Mvxt+FrsRybMlZkn/1YFE5
XPLj6JhdpDVnxF67p0fhDsGCsRJ4wH4qIitJCVptewgrW2pXbJPm3OjUbken+oZwC6Vyp/4B5XwY
b6xhBwNGeKRvzTo5D1TEkPrScyGFg7fgfgqtdIg9rKHzcOKbmpbMlCIi6gJmjWNw7pjTblWHFuf1
v2LBVfhZHa1cTjekqc+6Z+9YH9vJm4mu377aGKDS0yo6DtXESWTGCI9qd2GyCQJ8mwua9kCGyjAt
NiAuZ6mPnr8W1HYO8i6EO1d/RQmxFWXHoAVuBAYZXWi78RAV0Kj/GqonoTiv+OxDXk98lhmd99tM
pcMdMVIdJeeYanPMgFzook/TPOSk3PTNsFyIvil35tlM5/lSEyEk7Qs7YJ37w0GUg6bKjYrP1ckG
I7uCEQV1sxfBILAv3wxzPpOXPnuuHNDDmKGAe0SPXH7fIa8SWEGQnwO2jHafSyFEoD4RgjAJdWms
ZQ5/73DTzyXTR6ikg06vw+eNUQpiW/LSwGkM0/D6vNrUeayQTgOH4lwAvClpzfUpMS/+o4V9RwcQ
prKq4k0yQz83/qPlkSiipHTWMwulF7y9Fcew8hmKCVBP8BwVBG3l2kzSpZv04Z2aoG0Ds8G8c8bu
9mwqggSShBK/0PN7pCwapCh5pFaRQy13rdOWrZIN2g0FJSU0G47wEbMM6NcKMvDgql8o4s99kDTO
08f45ARvLv9HjLluOYMXu3V/dPZBANg/T+OsAUu9y6e6O2KDiXSNq9vMQeVzEFY6Bowh3PMNs+5B
Tqn/rBSEKaVDTdoiO/qshVSqadb7aV0JwwywSH7MO3GzSpeqKuObOBYocMNcsmrCYvqA33ljG8D9
CPP/2dafaz5x8UTQIm0Jh8+FltNLkS0YShkKccjKn25ZDbHATTjxp5GFCHwAA7Cg8xjwTFNhjXvV
E+PoanKdOxiSQ8FEJYGDS4VXRAE03Jo1dTpMOrAz3KIpGleozpJHxadBAHGKiTnzyzDLtK2ZbECr
dOCjQjmORXk8RtEKKhmwQndDdMh9AqZualZ06/uTt21DgEY/qot9VKV2jZSSbcTXL7knqhJsRPH/
zUXIboEuG+I5rt5goMywWQmjatzVnEZ2lu74HkuFGvHpACYBUDNaihVHeuFaW0npbFWJSrwfncBe
zxbcRhvwkj+BGQ3ooa0rr0atY7fOuh4MMDFmupiEAFlu3MiuWAtDBqpQCsqwf2aDxX+YCW8CEisQ
XIMIBMxiXdUaBDEvtgJBMNVB4ZZaGV2C+WGJkirk6RcEVSdS3VsV3o93BZ0kKZCyLkMqg31AkOAr
TS96GVaJZ+GvSNQJ7y4Q0tOCdScAsW+8a0LUjOdRCdXoOILx3uC6SJtVFceEe9iVKed7cKhs7hTY
YuXFdlwkUKNQdPpzt+64Xg3USV9W8rIKHwyEiJEpTwdzSvMf6QLzGfo4yF23MACu1lxlIZ6ZZpBt
GH3EgLSBv7Zfzr/tg2NeNL57tcWqvPiGxPhCbhZfW0gI/SwoWJK8wNN237JSAgc0WT1t3XRoQrE5
YmFrvnUAeJp3rS/QssvVyKscM3qfYJqS06BasH2Hejhrmi8wf8X6VVQRgEDEL0x+hoDDGt6CmkSO
IuBzoADm28EmZwbvdJ4JrXYkCh52Bwm6yol9E88OSzUG3E37A9KyZGLkwNQQc8eoarM0apgs2w0i
o//jaz0RifNlkv4T3Ya4tHL64XvlRdN6ERKwOB/onbgOWw5kO4uRwkymvXga+yj0i8WpOVUWgo4f
Oxz3JzorCLsgnvK5uZgybWGwkjKCKsJwYQKUPiRX92ILebHPq0BONNcSpeUIIA2tTrt78OB7EyYN
d7IdHWWUzz/8uYQyerLC0fFv8hjy3D2p0inZqBzg2YEVJHuQIKCvRArfApXFpNyE01pZqxcHL1XX
C0d5YLzEiE72SaRCKKOUFOYzuYnnNZc0bm4GAUEj/aC6mnoihO59M1xm+9/roIpeSgBhbPqBIkUd
G9rv1O7zWg5R9EMefFUd4gsjnIUXcNP0mgG+nBjIhjz7itCPoGMt74ygB69xGIIOdYS+ekmU2RlJ
9yCQa/+iMPac7/5Kp4BcAF+2QDzgVxjtTFv8rQgLdVZFhO9dWd/RAc3pFGsZSmbD3Fh/CiT3jX3d
pZX03BFrgMZmjP8pQndWV5PGYa8waxUJLSwT7ZIY6nhesJzdzUP8j5PUC/6tFXLGKFSg7QSmu91M
U972i4RYiydM2HR14uMj9R7wiF4sX60r2C/oriytlcqe6t728cMV+PU4jfNZ0XCNbKw9lllrSSvn
HQkPDYdGiy7WImoGGXAd7hSnF74rGWbb8TOHZe15RraGpp8DeNIUZSFQSStEpjRkcBMm5BzuPnKi
KJL5a8AQnSx11S7xAY4Kw28F2ECl+vT76ViNl/bh233+LUu/3AGEo09Qll/gL0bBU3ToKeGSrlkQ
9fOmPkmol/RuF+4n8hrLbxfNhtFeSlJihIrGahkJw3RIiS8QV/pPA7EUVbc9YDTus/7G5VmUVOx5
1o4NzMYZXwf8r8u7pnAvld661cZJZtuD/sZ6vrrKnehdArOyovEtE8UJaOkvP14XMUx2ydLWge7Y
RUxy1e4q7L5dchjqTptOH3RT27PiEIc6kGo6pJmrQxqi+YUVmqrqy01g9qbGLtP/tqul1/z30x0l
hFeotbpvnjpjHjYo8oHJUqA38Yw4sYMhgZroaz7oEf32tSC8HDH4+wtLLpwZKtppSUHBbhsNiqp5
/mGYCNVxFd9tDsih31x5spu/FaqPF64P/tjlkcwVGnekns3t1atGPNWOuOmS32eK/sBtrnvdFiqy
YrtXHdF6YUKjFYwxntYF6xpiHhzlscnQUEQjkyMMQ9Jxy6zOEU8RJk5o9MeHoUxyrqxdpym93rD5
YVcdrhpY5Jexvhn7u3hAbMAIlx+Z/ulFhLSlMrYmSNMkDdWTb2m8b9LK5JzYjonWw4rqjn/64LzA
QZkKSE9G+wfhcgkEvcE9vkRsKS1ksg4dlei3C6Xg76FNQV42mm8RV1ObnBcXAgDYqkTW6qrbR/1u
PUqcBV+/Ivk+cYAL6FoeLEhmTmqDLOEatWp0q3i4qcsnubW2FKZkUiEqI5gjYUqlsxvHvqBkQhcd
BglZcH3s7p9llLOmoxcTvUvlQL+z6Sxg/tyIUu/KCutjOoHlsp+D/8gPscLzhzn8or9InTBL3feS
YBiyOEx/deVadXbnaTTFeSYgM5ia+XnWxDc9BDyk3jTbOvV2gXKqTU3/QMzOjKHt106I29Rwoa/y
/qAfGKrgOusOQS1tJoypBI5EyVt5UhAa5Rn94Y9RaJbCRHcbmKsuWVFOWYRFD5f7AydwLqaF7uc8
rOhfTdU4y+VUnSEApNNXEVYIQoXelMa2q4I3L3y0qC7wftUoQ+G86evSHE1gzuedbW1XF2m8pn6+
uEep84OedKtu7A5NpFWMZVZR5sFdNjf9ow9Bo498aqMkjJyBW1BL3AhQCDVBX/rCxu1jWsRUY3Y0
QEtLIKpMDiq6wt6hUA2dtWQ9Zmx+1klayeLagFtcAVr/NxBMbDQJKf/3yzGA8k5j1Rnc8W+Ztcj6
pX2VtJP+K2fHWzqCNM8Jgn3RkzpcToBWR156YAxyma2UDWRX24fnlzLrHGVY4nCx9AjkM/08C48r
FceRjpar6DXJBWhAxMkQ4wodO1ehlN2oX/qODQmNz+x99lOIGO6fevzAovUGURJEupxDF2MfBrsL
BUl2Oe56G2KL3gm4id0VGsbynIbFYO7gRTAu+GA8gjjEYwWkmcyoQzWU4N4eGf+HKakVaNhg7uIx
GtcUWFWQMUKyrR3VA/l3MN1C4UBiELaxOEm8EUqjWVaS260AYRcr9QT471TrxRXQjQtdS7QQvqly
Kn4XwpHYTgifPCS3jzwgTn0XX7t1ev2LlNkD8jzNIZwkkLPkS+ddECZB3nWHbJMr5zE/gf+T07Ga
mGPJ3B3hzZlWFoev1Ydm+/aoyIY0jt2p89HMXT9sD9EU306WUIeqyLEPXS5OwuwXT/4UwoaO9Gim
KR5u8YgMzjx+LgqapgFcdyEwAxGvOR849Qxl+46zlW6XmfMdp/CoZgF8yBasAB2tOBFOUkPVRoXx
IiVPmXV3gm0zeYAPWMjy3VzJ25IwDKSoNyVIJfpvkyccKBGkH3GQsDjFLy3REZ/P014gORH8MnTh
scugxnlmm/MtoBvUd0f00KK/03xvtxvmAGFkJgANbskwt3ZTvvRtsJfc9kAsMcIHsS/olgFVvbVy
SSAzK0zUkZSj+fgRN3k5AkWL4FPUbgNTlUihGMpePEFh7ZhfDJ86rtGv8h2lDYJaj6lwbsLA/J4o
5DpFLoL/Kz62mqQSneVxmm5Yx78h0NVGHhe4PNosTSv61P3wn0CK0tE7nvMGY4GJAmhmoEnB4XXl
qvOfNgQVRhKjS2KgvNHIq167Gwa2z5JPZtKuzj7X3rnMORw/FET+vCCTWeGAHeg9h/7WafdOD6cY
CPCEBOKcbHjf3px98aGdS49/uOkE+PTuvNknYpyNu5mzAes78m/5KNm06t9CHEAA29RImTtyA1Wd
iNF0X0fRIxMgy3Qgh4XJMK02dLctTrDAEtFsgNijWODghCvV5RA2FGbzPyDk5NmC7lE7FUy0F9Oz
7ag7WTrnkrPVmKZalrP4hwqV7enl+LgAqtigOilAZxJ+/W22epsLg96wqQIrvWmrt12bmk5R4jCG
jeClwXHo7akq5F0mELkBqF5KBk1gJnJS02W0vKeK3CuMNtQBYNAR0KbGf/X88wK9PEKyDNEJJlPY
Sy5hHO2bvkntZo8iCBY7WM5QBHl5FmQw0JKvshOMBTIGJW3rvosBZlfbEzj9aYAfguNeUzTNTO/6
zos0sbjKLCfLiGee1xBGMVFfONJb6Wx9d/3H3vs1SP1llZ/RkL1CViDtcaNewZFLaZHivR18vS+W
uCH/XHrCsQBaNqYAL/BFKyDVqLpu/GOjT2WddAUdVWFP3j0qUA0XDCNoJ3f1l/UXtMRMNiAoxJKT
YjW1LceWbwhB5ApH3TdrVHBNJFUkgjdaJz+MDihF3xJp1uLGRoWUgmk6muTSh5IkaxxMyp1G8y3Z
JFlG7kg3iDsVC9krir34sNqyAdDhiK7UQ3MXdPaSYzZrS7zFHgeDjg/G7sS7eggm4QxP40bdZOMz
At+JUCZkhKJMAXmZMzQtjhYV5d+3tIiY3oS0GWzlYd8lTA4GQ8R8oGoLKEbcSRZx6FEkyRYsBm87
AvWDsxZYjkL2UIXadkHS0Z/R0ihP3nKcUkZzWyNOc0tJIl794HHDbgzvLHfo18w6VrGvz1nspgZB
B5ywAgiAoVx5BxaOWDd5dzvFmoIoTTWpTM7oqWXlsrR2w0nWDDyw6ERD0Qvd4JtaD4nj45mjaw/Q
T+pi2pDrD1nY3QLJRjREvPgb1H8crwZETMjvzuBYBPVQi5IzAroEgcV15FYMVN2cJpLck/wtHlNv
rAF68HJnZurhSJ+b38juV1rNUhFPg0lkdbWgNwERMS+q0+jTvoFBrlPZnCVVUEKCPuLmFpDK8iX7
YPjqXATnq2RnZCV81dzwsSwnJ68YQnJ/QKkXDHf408o6QVjcza8bGU9QHf10q3V3Eq2UANOtN7Z7
Uhl3mXAFTzw6eTibCDxXE1cRM2Wxd6PuhEGx1XPmeSirgI9UNdndYvcIdzpS1mRIJJAwL/q0Ugi7
NVteyQmLTeM0t4ax4KF537Gs817bSS3Jx0Fnzm62hNQZtnG09cwzCmC8ATI5wNEP8OJ4q01yiK/2
heZm4jtLlOJ3K/k1IHBiFfLCTvHM0El/jfgiFgufiKU2srR5shH5uZDMczSTJIcYixn46uq/2SaI
XGhax3w2/mKoFxyT60GaLQbUp+s7mX62KCBBJTWxRav/fni+2UtI8QHzk0aruwX2j9C2UkrUisUJ
j8cWqasvDLFtAe140V4U8LqhlvuG/ZG+z/LpoI7h9W4je2a9jBktAJ80Iw1eUO70uyqIJfL4+CBD
tB5ZtCj0S+csFYBFfSZs/YbYUW19eX0iDIY1Hkjq/3QrNF5agTL94BFcqD0bVNXORy6eQ8ntSHZX
8jFmPIk1qgIDHeHUf9FRj+ML4KQDz1JmcG2CONo+E1RX4gKaZJLFsJx1Hq6zM2JIB/Pq2OGxukAf
gBQfwgBw1JgZsqizwKT7E1u7bq4OFhpiQOkpgcqOOpSP5yMiuYmLJhXdDHiMNpYi94Sz4HdZiIut
iuCSIKkvrVRWHjaeEStVTWmkJ2FLZB5mcwsCErvDNfn4rxyEiTyF/x/2kjV+8eIgavL3mLnUbadW
GzPw3q5j1CkHJQVRY0auioYpyVl9KXtxp5wxMkzo1MQ8zrdJIe7EcE8g9xQuySdcmpX+gMeM4fXp
+3KLfwWCoQkrAPYy7jVvUM2EXfXudzHC+z8z72zylBjBCPOPrbp7z22+L/3XS870REyaMpBrbEW6
7b2JSUDKm1h2z+KOPrtECSdlLrxymdQf87GHuwjwVQMYDDrzex9B5YaQWJE4PPgi+qLE4u5TYzru
ZrPjL/8l1FhDMTHOHNr6NxXYc6UVq07GWo1idbyCGRAFspODt5CxSw5AfSFfDfS3V4S98rEsLGZL
oQHSFqESLexjHmyqDYGzFbZM83fyOL0RMmC0riUjjG8ZGSYqxXvlSBEFk07T3yvwD9MUe+Fa9BW2
desyYkh1A5byVUJJUUQ1ywbVol0ouZxhdoq+rkwqix8eSklK5WPXYCQ/potHNigSYI0XDxz7PuHt
ZThneHs2gH3SQqfK95FK+YFBra6AzzoSQKv5+GcBoR8o5a0ei2nWi4i4Xc0YmXloFaouuQE+je/h
Lh1B/5xfEqI9JNOeJQxgMsA1BTB8t0bGaBTgHc6r/G4KpX4r5tfQ+V3+2FBZLadYqw1+nBqFuAQO
TW+4uNiaA4qTXiHEkTrjxgZjM4p7LJ+010QyVPLjndLrhWj//RpdigAdsmD/cZQaRkEQAqHID2Gu
hxx2j+9w4D8OZmCgo4t3CwUAurrmlwY//QBi2J5rVz4nzdczYPEOCV8enU/SAXL3vrHWNwHOGTCP
CGOcLen4PfP79BxY21QXxPOW8ktjQ4OafLFC4da2LeuJ1rpEkb4FIwmRyv8DFaBqjilDYnNzQri9
wPdSza1Sn3PnY5lnw4Fqz8CjgoNbi38A0Juk1AAV3dBYszhiJvO+M45wAxm9xAPsY96VNKlEYNIC
clDk7nJKvJ3U9kjqx1jl+vjrxahBjYVFSmyqIZTe1muJR/7KTPXXOQAylvE1uM10eLrUaVKp7b8m
+RelHFxfrEmqkQ5fJVvLM16rNx2lHkxxRF6L6XOsRAmPr8ciO5RwzQJmeVRPJrp4pkHNmExSr42Z
ULcd7W9pW8cKkxHJc2GmmqwcCHgheMdkbsxpa9CogsZAbUfxFpmaY49P5XJ/4UwRKrIU1lg0XqxE
4xGLwNE96EWyiHqGnBG7SLq/FFRUQjdosuACxTjH73HlZzTnZnCXUNXghZyUynlhNTDP0Uy99BOU
YlG7y9vfOth3/EqEV9Uz+28UxkCljvySjX5kDz5lE3u1hpV4KdIc7cXZxBHpfP2F0/QeQMWh0lfl
WjP3nuCS6SpN4nXz++JHKxzoBOhPfsVHHtNhvmBefLw5DkmH72idJKidADzJsCW6csSCFVcXfYw1
8S4IZDnW6acut4o0l7R+YjfGoSOdQIS4duz8Edluc2cWJKDLuLi+AYnpFkTWki8fYROZJcYaVIqI
LHRleq7E/z5weuFNOEKCR+UQTTKBEs0MY4eEZb8fcqT7uDz1EJFEb8hKf6n0bzW9Hppm0dc8dpV+
uzna0761ldYQfn/Dq9h+HFS88/ZG0NLP7Tep8rsMRXMyOCuH38+Pr2bDZkRN+WCa+bNRR1Bxus5I
RoKt6rGc6Znd1N6iRjXSYPjoVjrgusYpRiHWDsq3N9kKZXXIiELXUmdxKfyNQO6vDNu8sKAI3wlb
o4NiMxZfiyke/9pJPJ1wU06f77lIgyVUC0Li/OAcKwX2C58Y8F8kDxBtsV2kdETg+IWVaQ1aEbZO
NKTLvESijYecv1dhU8orgPJBajz5RU+9U2syqLR/W7Vi6/d53ERzjhMeIu1IxuU0G1MAWGX7sva6
aV6eh5hLIFwdo+qt/IFdRER4j/vlNqhVJNvY7QQeYUYIVZtDnp75XdqUYlgRcYXAtFswPgC8NpFz
zdM2vzC5yE0rfe9CGVTsPjUirb0UlxC8lYdHPRQL4U3m9qB7HGyCLWKwaWjvYbt/a6KqBfL6FKeq
oVfOPR/AF/nI3yuXShYHkzLxUl2ND70upKXDuey0b0TP4oDJlul73EeNqHokn7bDe86YlbmflzzJ
jlxaxsU6xUVsqIcsngezGTinK+XZfBkkFSpKkdms5HLHl6ASPSNys1OmHoff3NDSGL3fgtUOvGx4
ADs4aV7H4gvufbONv0anHjA/nw11EbBVWVDDHQhCWtnmKDngbLzdbysjhCr44M7KEV746Oh6cU8g
qDILjETww43yTy0prBAovjXHIPi1TBMh23fOtKAsetukZuI21CLNEnDWVvwVuX9qfqyVHi+diIaX
YyudcIu3emiObAQ3QKpO/jOq3sUDpioAPiyrpwMLB3Uu0ke6zx6B9iSdYWvxOC7wOloKWSaM6xDO
Ka4XXTsfF4Cw/tmy79W2f+xDDM/7cHUlbZMRF/ev8ztZ3cuRFWHSpNqFxZdeHM9+TMdEUVnsevXY
9oFqPbzqNBh2KsbLC+oxi8zjJbx/+rx49x6ld9Ymh1mQmS58bTLtLDmpK1fctG4uEHqMUn19qO+V
PnPocNEiLTd6CJtqAwuX6L2UbeVup48Qo+BMgj8eN6kUddtoqbNFX7FHvkL42lr5xlkkcfVEU5U2
FEEXF2FPRdVXzqVaz3HPECJrcbYVPPtTuiLGb+WDLQzr8VbRqxR+DeuC7qm/+Jz7ml8MFNeSia9B
VR/eqH/wZXcrH1vzLbgr6ZsUFQsdt/ldSyY7d3UFkG3wtpg9XphCYE5dxuLIT4LwvP/A83ltlC5V
5BFt5vY/hZJpyanQzKHLOENvHoAkS80kW+FzQYzb9GFwzBaYB+yuwykpIQXU+c5F4capbmbRhVa6
SNP62dJMs6P+CBcL7gmSg3ByEf1kbneLp5oGbOyaJhEOY1ZHBHIdaRv2Kpem9GwlNF5bA4/StziP
U9AbN4TGF4g1PHk++ofYyQc+Q1dM6tpFYyFjGJvlEAoym40JmjLso6m2R2y94IwY3GwJ655nwAOF
+XhHL3Y+YJrClXuSl5PqNwUUoUZK65xDNRIUOhUpooLBh5pX78XdrpmtXEzKDB2DgdvpNZFZzPfN
VeqDBwouah5u6Hw3JEPOaq0A8Q6kLnu265dSf/+R9st4WDn1/ozZB9Y+8/9WarBegn6VrqoUNb7G
6FzyYSca8oqE7sSnOS2GXt/4aBsgvy0xwVST5YUTQl6d5UirRXXcrj0lx7OAg+/pjpOaZpZH+jJ+
+z5XsBJtE4pv1LQ+FwgFGsM5O1z5Fi660QkVxxkBEnTfYOwR4JaLqz4waktHBnAPMuc2aaWn0D5B
iR3uSn3ge7WWKUDe6BB0Tj8KfdMyFGRqaYCLPogQ0OW4m7CHIMweZW/+dCxRgxQ8mDD3Z8YrYN12
+AXrWO3DPp0OvTZV8WqAfkMhJXR/OcL570XIiiOBFNfW6pcQnE1QYEl039NJX8UjVfEgtDED5mr8
/wrTCrOgaHGsjBf95Gl7bT64UGQE673bgXqmkDo61YRd/6HhTMURo+XGVnkjq5XjaI8/KHQW4C2t
SL5cQdf6oP67EpKyZ6J2zx7Y17M+9lAKE9mzANylPfk3N4p0fE4RNkJjA1+G0QaxvCl6U68t9sUG
PBmjbEbBZE5Vx9kmyJXY3ItbVKt3cNYd74L78hTgsKqE2oqCyQEEYbSR2CfOqNkGlw4osqXzXzE1
rI6rARFAN/89+uO3y3wTz/oDwKMR/5LmUfg4mlgCfhGB72UYfrXjct3JBXEXKjYILrasolsPzhva
o7G9Owqsi/+Y3o3tiV5mSgVUFORcN/xsRgfArWyH1MtKxvnlMGc09aSHILgl80nMr1b+KEkHA4qE
lhwQfYSc8lF/mV+7iZrEuD71a00QYpi6+Ru53+nEWS+P487C7C55tYZmS2PsnLWslBEIQtp5ppWw
B5y8A01qHkEZCos7OtncyOTjEt3w3+gW5FY408aD7M7pEHWNwf71Mh7i8N6n6JHhx86lOCWl2Q1+
tAE9nBA3FikfazYvfGCjSUwt4trht3PkB98K6xd0KdqxZMRk5+b0koo1LG4ak4LNi0CPz12ldyUl
DQJzzO/RVOsRA5W9jGB/BwsrPsgtBTcAWxI2B3NhKryMWsMSO2UNTzIYmDJuTvhvkeyLnO6vzI3V
8r3FuxYVIPgE3HpCOhqKB4J4kG3bfD5k7FZXMNBFTITaNXOp4i1fpHF0jh0us4b6hrhoRcRB3Ni+
6NY5TBrTNhSbynRfF5NgBTsz1IVguxMwVXyDhD7K6xC7mB42QVcHt/qtgp1Y/1xfGWiIUkvMqBOS
KRi2P2ZfmW7GDOFBd4xWTkNECPS7jb1yjPe4imbdAvky4dgpn1kqwN5OxkQ5keiPucoJiylFlnHC
bk19PU31lcEy4Uu8IB3zlSrFZ10IZwY8ONFbW9vpH9/cim+CVZC/4pZm/vthOaDg/spapJDm7hXI
WjxOZ/dX6jAZ0nLmdLfmwCMNwv8Nj/d6fABXV6zje10rUvane+mlJCNVzcv/5t7+yAywAJkOpf3z
3MNTSCSDOBThG9c8kKrUfQwrz2R78BQ1ZVmd4puJmrXlGvM2EZA6k7REtK7tJB8CY5eJUYYv15SZ
r4bkFzYzfh++/SU2VCMbp6+kx0FX959JMcTWxMUzb/IbZ3r9yZsTtStQW8kgAi9uMVTjsqJKuQRt
GbNqq9qHX9cUHKYpAFI8Gsye4Yh/NEL845zis8Oe0sMJi/7uEmF8gC1K9+JBdSYggd/V8MmAamWc
vSRYrLuKYd9AH9zZz1C6eMLsNCRHL3TZ966GF2ht8lbXRh7LBkHEMjc+qnyrP/zglgTI8B7N2ywj
0k/Cj8AXmJCUixmTue1S3cfo+TwOtZaaYaV3U7OKHgnMRjj2IDR3tGdZxF9NTBKkhoTbDwO5pryy
/NkY7VRPRr/6+8XX2MKSIp5OAZlpoiBffDJYnHBwGcZN/hPAAbLeDrHmF+PQTBcXHl1bLzjzx+Qs
MKVzG1bTmWcqhEtzjBEdXbpa82cPP6asvCDUD6kYcWedfUCTdAf7vx5bB5NqwXNUDfUG6qUnKbl4
we4mmwQew+ZdY/g1TUKgvoAe20EUNe+bNXkQ8olCER+PtDpuceHY5dm825KfsUfDhjEiGKdma7+2
MC9AIJL1WXLdv9v280b/uYCWfAXT25ksiRB/3EqQWzzf2War5tXZ6LimzwKnMve92FWlCrzEhhVL
DBaluriKxP3X+9npMUBbFI7KugTwDRPmGgXYSgbFPDPUGuHaExClENgHR0O545DSsm1zmduOFEnE
DfNX9N4nZZn4178o+JIHtPR6M/ki++bsH1h6gZtFmyJr0n1dOjQ28mgkkoWqyj6alhM8ShNlT7Ee
QO4Ot4lzZ0yOpszjk6AIwiWgpBBVAK8AN9iZN0Nl4uLvmNh40zJ5bS324NvSiswBJCL9ltZnSBNX
7AbyuwBuaZ4T2UzAh51tXcVHas8seOzpVwenfaJqNaKfaeyI1DZ6eGRXs4Nd9xwh/5vCTZcyZJ/x
gQnZ5l8A2hvRZfZ4IbSMqdbqD+XTC9BMjzjjM7VODhBZJpGOiCXqLb39xHiNGobaZAXRiPGeE3Ue
EoEGTCNRUxgtFCzaES6/aDzYK+ugMP/4gyuXQcPU5aS7gWFKNjNn12eP0vjqZ9+3n3f0Eg6bz0mA
6C3+9/4bKC0gxMKVfO8+cVsr/9dwi6VedPLuLLPZzPOlYwwSj2Pp7o23r+qz0RiCOrY1LGLlw1ub
BO9vwnSlJRshORNmaBn2m2TuizZWs2E+SYD6yL239IWm6xMnJhhJuQdkHWjZV+Yz6lWcwkthcsBy
deihaT2BGA3UWvRu9DQxP2T3uK+fm/yf6a3LR8aXKYntEsUNcMTBoilo6kuJ0KIa90Zx6TGJ1app
pR1D69Pzf+2yozMieYXBz+7hQXRJdOwvGMh7JXqll2y7aI1qhUHuSZ6jzm5zqR4aHCfj9jIsOS3U
ydt3cWfGr86vMtULEoDaQ4GgMKC44y+D1v67DbamIcvFItovBrNWe5uItjKY2FIv6yA7DR+M+QOS
tyFxmPeiKYL45zduOFriYfyZMAWBtgNkkiZgo7cKUbc/ylzCfTUSbfjJml4CJYoQqYEGuoVq/AeB
I1/4WhJltYhBC/AFH95iK8YjG+ifgossFTeQuHxNgv0Axr8GZVJ35WuSAcvIX2ReuyCY6/Z7HHYJ
FR45B5Hsyam0Yoe9Oid/LXvrSMqP9Ctvh7gh93c8mmbkQxWTSWMc/0ReKsftD22ECd8K85RSm/5z
FyYHNTaZLglgqbk+T/9ziMrHBO9wp1ZiX6HDUCHK5t7NHxQk7VgEI+y0goXjk+3cJKFbiSNq5PPa
egx/cBiJts1Xk1iL466uz9hysTQMem8CvNz2ZgFNOYHH/T4E4ADwUsqsbf9cehPZoBP1osGDU3VG
VMjeV4dOLWRNoa8VUJMMXkGIE1Gu2DY1eO/E4b2UM/H7RK8V19APJgbIKpKUDwQdJAkdPawJ4koK
BICrzHbKjUY0QKGs1AuuwDj5b0C2Gne+g03q55fj+ZGDtsmG6d/2aktS9iR7Kdr4c/DGkQZ/C1LH
+bMQrIomsyMFCGEjt3QX4jN3SJe0TY84m8C0H/FRcWdVclMDRJKvi3mz0i4mtz3kWwh/WOnHjTEo
VxJDCG6oD5paBLF+mCwb3VirDRvtjxkeXbKZ96OuQlrH09BT2ZPKkgl3qUZkG9cyI/SvyV4zdDJ0
7OEViDgT7jt+tbcdy+t+UObK9F5G1xqke4zFqXT0vxYv3qScOga9gon/qATwtspd58W4GH0cPtmS
boRmwMpjzEXIUg5mlOodLy/m1kjRWM5Az3hvr+qbQ0YCbPylGgFX2aFmaKHw+9OjmQtnDoCF8DXd
UscpjTAUyuOTBKyRDPXB5+8mQRS3jfpX1LD1G7KZwIgTSoM8YeESs0Ev+YxJil1a4t6cyywxxthw
mTAP5MXDFWslUsWZJRCOk7I51A2lmDUXhMMQExxw5UL7xRHjIopF/6txGzwzTeAFxu349XokR6dI
9NgW5wNdyN5ixl0qfCobq14cmfUNJAf8aFyc4//740D4mLuiF02S0xxjjYkZZ+FnORT4yBvDBiqB
rcroPVYfVs1hlebnvvXnuxf2KplzJ4e5AOxiH63fbKXIFWq85IMiNILUOgV5MZXGKosG9iiHZ1+m
yFT3a2AxnhdtD1oGZUIxXeIIDk2QcNF9XcDPmbs7dvw6l8+nMib0nmVYTEbEsMVUoa4+XFtmB3HZ
PY0Bt3umtF74OSiWPJOpCJkxEzG8baH8BasMVXirmv5KwOD4Z9bt6vrKwzy08iqJDKiwKGb1d7Mp
aP2GIS7vd4Z0L/rlZUikUDoKadaQJVzVszGCYuGkDu0dEY/zpYgvPnUDcDUHpn7kPBLKMnwPCmN4
dwcUJoSDZ5pJ2cXi1uFhRFGOO+AyM6q4cmsJf6obhlu+inkwEwwEmE3kVbIsr57ElQyZTyRgmgu/
2f2Xfji4ZP0WStAUfitAudwGb4wOp9H0DZREF88JOocHcRX7u/+08gyJL3D3J4VU8wmGMlUDLQH6
7wI/Y2Aslxwss9qyrjQQE4UhxbZEConAGTvddX1bWRE4gb0Hjv8tS09o4DQR8tJ8G/IvbHv1Rpcv
Ofv49cg2UP0/XeE2K7zfPpdqoRFGi8cIVKY/lcrzMeFBJ3Ak5aXQfL3B+4rj071aNf/h3pRu1v2Q
Sne2/vpEO9ZNp4xNb7otzzrmFoHl2OBbj3p5+Spbk0EnQopPyP7+HRDioD3iY3bYSFbhdzdQhXL6
V404Ud73gk+GDfE+lriJ26P5IckgzLJkMPffkQ9YPlf8z02wee3beIofYOjEQC7daw3IWeK3DweM
JSH/HTRalyvfMQSDJmb3Q06lt4IEcl8biU/R9GzwY44Ch+RhAECnpS+rBBX6veAilinVEC1lFvvZ
FuFt/Ee5vlrTcaKwb6EaVYyq9+ZiBe06TYyX0UeGvsIPubxtADtIomuikTisKH2hG3ehi0PSkGkA
5rZAHO97rU04TBblrCVZ3xzht353aipnnuYYSJYl8dePas/7NOuvwiW3gZSdh/4qX4wyrlvcYMHR
MsFD2gXmrXAQrSe/PG/B2xRBY3rCFcxVTVavpuOs+cF9TR9+E0LsPb3+MTeBxZguffxFxo18KJCm
tATXXmyNtHpy5pLuA1u9BnSwL6eupCbJQ//R6TCQCfY/pe7o696hAA4boAj32IYwuwLrd4HS1gbb
Wka0vNEl/YG/PpEJwW8C+35eMroGOYcM9qeToAmIjjo6y0oXduP+SjKVWHFJTcvA+/BT2DeSRaYA
JSc/Zq/wJBQiu8bAJ9mM6GMU2SbMNOYn+KAcAGo3sbTagfRemB5PF3fDeBLraFqx/WNHtksomH2O
Nxcqo+i6kMcwJJNqKPMSPmkj2n447fOGPBK69SYpYlj7PkdG/KdA969GmPQAzwuCXL/SLc99SEm0
/UftHwmmq7zLbRXnyRGusgFDJ1ViXXMWeGkM8iCJQ1j7K21AebO0YRkz4aG5K87ONOVdMoBRLjV6
XUcqc690emUlePOd4SSUC4lZvXo+68iUsGfCxa5OuiRpKcEnPPAijliHkcBeEgSv0uBhe5BBAn22
t0xtYTOt+0amOwROLH2+At0LbMLYIxSRQBZ/1Q2qE6qOAtdJvj/NpL4Lh6ayEi1GdZKJFEEUkDB3
MoVNcnMUldjnKa2FNsykyxs/49aiNp5c/zM5xR2o6wtdkrHtyjtsfPudWi7fqPAuFxxQavUG4R12
0mHWhtShoXn5h0uAo4Mwk4nLUjPGNCjk751sm4Hg0YQGBcyLjU7Kw1tjMUxqzqhQa7Sf1ZkllMdy
33unv7hoaFVEiZ3KXFKVpLY+tF1NVzK61EvhYsc0xrYyg/lTrV0DPtltk5HmBTMowo92ISvZWU5V
+zo6H1wWkUkaII1lYs1+jJGT2AzUt8R8Ns7G08XP8hZiHG2zPJQ812PcYo347e5MrYIljdNxLYoF
88HYCWynfhhCQckLVVpTmc8Wjr1DPWDpbsaKSrUogluP4dIkTVRWZN6EJbV7C3FUfaCwswalO7Hn
sF14NaruMBfE3pNutYJE0yu0uyClz/EGK8yehN+4yS40SGMRE7TsvdVdJcb2FRe4OOO8MsJPQsF6
qzyo6Wsx7aHFQnYgbbey+zS28G+nowDvc0xBWZEjQa3JLOQs52USBjK/3rZ2Rf1AhP5o5JB7K3Ap
+eh1234IzSZ9+1ZxN66InxdqShfGyOV+6x/CZ4n5zElA4YT+bGOkVDDFD37krSeRMbt5uuB0pmqb
GfSFktz4hyvp6C7Ex74LUAkU8mFiqv8QyKBn/L88VtLDcq6iww+DvDejplgIMUfDO0nwPnGQjMGy
oGVono9fwnPp/BKx3hZoXKoRCSLKRpVNBnD3J4wXIHYvUjrFFqvroEP6m06BImo3I3byEUaLz7SH
BnOzNzhJi7Gych6/9QLiQfZwSpae7W1OhYjZVLtiaRntkj22zNKYZp430fBCaMOaZP6Vdv912IPa
7Q7L1iqvBNd1MvAg23tXUjrW3IAz/rYwlRKMAdUkuAVxGv23rDllfMA+WFk4T3CAgloD2pzvAYwj
T4pXDKddUd+OLo6Awe13VOHxBPHvtAu2rLLKf2CVd8TR8vRjKmUsaHQY5T8AE8evefYk9C+/pab2
Eue80QxNJq5P8MwOeiR/Zrmrd9lGv005/yHj/eCbgH17dmSq7Wx9jJv1s0ctyYxrthEPj9ylIdMS
sWWGtODCtPzqSPUnXxU79LsdZQa0nfR7hpkwelRi6wGlkyTpKL6fAYdmf8ccMlgR65WkQr7gWiN3
WeBaR2yDEsNbBqs7mYZH3RHk6X2+2WvK+uI0xW/9N9Mt5yhcpbMb/IDkxzPlCIA3klKIngEV5UbD
lEsFm2zdNN8dGpUaAeC7Mlak0K9592FjYGMysmx1Y7Hd9ejgvkxFSSSUA4hzo5rF9jr7t3fcdFHa
QLDWoEnn16RzmFtnvJsHaR0tYMDq81rsS3ebUfyJ0exqxXIDUb/yYl0y+WApoKE0TLHwARzw/5hs
bcTd5MBuw4rr+mIxy3f+VrXRZRll/t0kN+hAvoTKd9b/mQYuEN+EG8FduFGi/pnf2SPFnooN31Pr
6jEnA6dFP1+epIBRMctdahcgvYMu1D+Yr7DQ2m0r2HIEhJi3u3YMIhCSKa257pZjnqstNAajeQ+t
PqGvGgg0gnyRoJ2ulTdkLtH1dOa3+PFwe9hNqykjkJrI2rIbHvcx1rSxAUvdc6s8cHSB0XGDWWTC
G/xcbhZ60n+KYntJoTEvG4dH1W6aByx7pFDNOg4iRzq2/5Sn0dYmcNPakCSpom9H6NsxvC/JQFX9
fSmV5+Qs6Maa8iZi0WDnej+waSXzmfUfhVRGCwgsDplGXmIY4yG4TB2IR4aoyICJJM4UQlfrRWuw
B3ObVyu3W4s3+0k5ZPEe4vBkaXqW2CWaWRoEKzE7tdBBAqitLv9G7gqPmc0LKZHIvU6yERPx1CXv
iIxYU0Ix8J0tysJwgVLucytpdiYSPElkAA5B1WmDYL9OxSlWG/8rQWSxcyKR7ldd6KwsD09EJXkT
jFYwLwGxSErwe4Jjic1I73Mqfw3ns772pQWkO5QjVV0nXlS+bCHfHOA0GcdiQzwltbCmzHyBAIeQ
aaon13LP1G9nnB9oXtay5nlZHwrqb1qpaRFSCibmz7zbFWSQmbb/utpW+1wpJ40rVDiy/RvAfbet
m51GqFPAvXLcPPoGUrKc+9dp0cssV7YF/n2GPxei6g6qQAbFfriuwPaCCZWwE+LoSRJ8ybqeTF6V
CDDbP3z7RncjA0X2cc7DOuOlPoX1aEXPA5iqBlEULXVItQ3uOiQedtkbsvuU0Z9yWAB2tuUEuYI+
eHqQmKygXMAHjuaG85pVdaerebCwsTHLOrttrG4JS9fT+tAQwsMO5YecssEV1gTZvKdn6yUoBvcU
sVD4ZCQtiZ7YpgrDpMLkp7gn/k5LWi/xrEUefG7MvsbAN8+wuuqyKe7xoBn9Eh8fap7kgLRa2W9m
c63pYk+yWaSODeIQJiS7FY7BK5FFbtA3dFsAHyi8zOn+5AMqCEjXdmS1lyBmdgo9CTufzT53SDLi
CxFjqLgvaZ1s3zlj3q58EWsHUZAeuYpPg6rD5ynwHdnv0SsOpZ7vXlE0sijjeERV/w1T1agCJW6a
XybocR9sgTyQ9w2GW/WXWoGIhXlfRSS3v0xxbJOZey6H7fYSAzO2/XiMKQQNFsUftOLeLD28aZag
GZqdDQLd5hL3jHEjZyqNsE8nH7Ttxy7YkE4YLfoDQlOFeijLs4IlUX+SsE6B7j7TY1Qh8X/jfmTM
QFA9W6bLcpQE8+MMRFZD6h8Gz1K56HiKdrIpCUGwnGpfLApJu1l6B4J3Ok478fV1TIVrvhtm1v0U
aW2Nhi7cmR43eOWL8I/h3uQ83GQv/kxEP0JylZHTJzHiJbgd2fu7UHJ3s4fNOLyXpcDbwFHjRmBt
112y1MTGwtBTsk5NbzBuYwGsubeRIztPw3fQdZ61rKXr9G+V3/wyhzzTdH5bdcRXMbr/bgWmUQET
PZ6PKCB1JYeGNmQB3zxBKBkudpWnre6tZ+JWSrLGQhfzi8sNwsLJKnmxZtelKcmxKp8UXbkllF0P
PcPRJWlJTSdMhCBrWUYLZfis466BWZw2uXzTWCPKyw+1EotomXazHWTYqBPKhecWwUhcY9fXlaNL
aJuv0ODkYkCLoBQywTyDif4SVyfOP6fqBE0wAj2r61DRE4cmEof3zK/aXhEs7NjD6hZT5icK4+Ws
n8o1UbUisDBCo6aNf8RaiOG1QJ+XciiA7IePlKLce1pMJygAb8v6uxOrK0McsrCakh2cqCCHVP7s
WfD8htfCDyx0aEvAYykXGJK77YuMjNEk5VVh2ig36v4OY80jazAZfUGy+yEDqRfHBUB0xtwQUmgk
/gs0924vTUPrkGIqZ1cS+YVboMHZZ1dd+cHl5qFLpCFo4H7f4HW9FmNArjEyIk612zEYuggj6B+r
7CtaDC9czuygrx3bEUkbpyjA5zz1Pq80dKIs+AjFBzIHEZAzYfdktizOi07OEfwgVwWWfkP4TRNO
krbJ5vMV2DJk0yYrIn7PdB9DECrpo+PV2lVMedowawN6l/0lPy9Q1PsQJkklCqIzglN11f5rHl05
s+ueaBCrLEOP9Tf7DHcMemCdSV096ai1GJb8dvq6lWbr/Vp2a9HvAg84TMoYdkLGLSALhOpGv8/E
iOpRYqVQNNX9nB0NnfiEPQsQpujgJ1taWTooeXVLoOoDAfmBkscpZaTFAhE1fJzomy5RhY+OyVb5
GOPqUrlepTa1Cn2R5hKvLqyfODY07Y1eZq3WZcbWM2TRil7WOP5YfTmwdNCwiVCjfrps8bbpkOty
Uvnj1qEmr7K87Nh8EcnDXfwljwdOr82AGV7sjb4C4Avv81yWMl6OBTRIkcIKyFrFWDX8che5Fil9
mdQAkuTuaxYPH99uxMpYfSllwuTz82JMijHFeJDKUo34cIkT14TVX7LifPYyFOkps/z9YQV95Vyh
tkt2DHPj2aGNpxntQ2NalDFlF9bbHg1dZjsK/0swTKp4hl/Msnpg2KkP5+QQygXc1TtmzxVwgTJv
z0mnK+71xbJHLJnLI3y2AcYrV/z/ndyU58eoTzCo4s9SesIDZXENSj1rNNIFZjQfqQvtAD0efgI/
UU0xg0nbBGZ1lNsTHeWyPXEJQEkURZuA1LaQxWJ/GGpXAQ+pbbJs0UvkuRKfNVtCSrvuCRTvvv5c
4UG7hKIZNUQMCeAMtOH1vzEZ85Cg7NIFjPTEUkocA8Q5T1T9vcedS3/ztw113a3QJS0KPV4ZeZPT
r9hiZnTxLnfd8C85NC2Ombl/K0vooWuVVD0OCVL4mQc8CbVEKeOT5Zfgbrrmh+sflWzPBHLAwFU8
9ZdFjaOQIeBBuLXFwThgMoH/MwEcy5Zc2+/G+Km98avuwkgFMiUvFd70QomtimPFSE/xP/VEPHb7
ADx3SR8OqdoXXY+yhYoSYma2PZv7VCqJGqLmQOnsCyPlulwYgaUov3EJ16iJcQnpN/C/jwi4yRYN
Ygb8cE5y7qMN4iXaVYjN4ZNWkQogR/M3RUZQNSCo0W5dzDOOOLzAZa9isI12FYrjQBKoI8EkyuMZ
y9wIGXM8P13n68nnW+HrBPCiFZs6ax+te0TMVh5ONZ7skwX9wwt6iKtMdwDshGtZVrs9sAyLEbNA
JCACGUnSgj8ABa5UjgywYCME4xm4Mc2QV62Tx3BJawG36GYsw2Ih+ktNasPtAkEGbintn8YboUfA
4IEeObw8FoSAYlL95ckZo2ITKcZhpmUxcz4cMqeAGvNbDaHfNVA91m/ErrqRVcdIL668xQjV6ArS
Af+EteS7YJbGHBUODgJ/bjFn/Cn9MNcmi0SBfjPO8hJnYl6RZzInLTYQwGhUREZEKaZ8fgN5ySOw
VaFEMhBhX4JwIZ4A+JllEISdflESibc21pHJ6uZ4I6Qr6w9vjDduXQRrEr/kTn9YHH0JHHWLmgrw
zv9JbWEIqbIA070T8ZyP0LAT0hThI9ignjTPLsVbYOhrPxsw+VB3UQks2oplq0zAsn9ngFp9YXUU
GFFY3pWyJQ+7vV4Y9QM1jlIeywDIdqe8I5cduiDnrWqIfzMtT2LGSzAwjtGawa/USs4x15YcNdCp
T1P3N3N+OF+Rz07KRXsnl4q4wUbmKZbr9zLEbxqHpurc/1ylxeZ6Ah4kmxhqwAeJJyS854qg45NO
BW3x8pcwI2Ec7GxggVjXntyNwNwijDdvCgDPWL/Yu6Dx9UWsEUpJ68AN33hXYv6JxK8lDlNFeY+n
7SBsjo1eUDRcy8tlL6FPOHXHfWR37d7mxe22yO/Ed4HdYwGVKCmQfXS47Wi5p8DbIc1c8kte03EA
6pgDzOhHRkcuh+2j0WpJd3un0FEtvHLymesxpCbsyA6ZqHXwBjD2R6vgKexdEduZqJzO17XSy6ZC
3h1e+A856n8EZmI/TSFgXV3RZg/8ETKm4hfec03wCruXtC/ySMCmC33OqLXdweCBkIkMW6Dsog19
Sjh7Xlnzck2OLGuiJnRvGXCCD0auPKzYSJN/xPh0nbxSWsAtNoK2IJFvZgW2E1Ja8PsKWPzdqjCu
vAXqFuf1UgylASKaHcaNLwBhQGYOmMlA23ZE4zj3ggvAERJQ7gI67SnlJVFQC3C+pfe6tzw2hY5t
HbBVzJZFyvq69bxUfctXld992tvWrhB5uXbHqu3OnRPNKAz+af4j/+pDlZzHCpmvIfpU3TuOCdGJ
uEHgFwtMF+o4r33pUlZlLDfloVlaZ0FkA4f6ovpu7pHZReSf4AGI8NQQPrU4/jo1dpP6Cweh5G73
040I9eX0UULqRhw4LMkgz+/9UzGPfVMPjdd+lFEBbg3PCp1Sf+oiCGatghTetNplXUdboLARbQkd
fJFOByiVcbkzGpZf1pT/QIyOgFHIBdM+6Osv8sWK4e3t9CsDjxbEOpu/6z7O3pbtXeHa6DWmejjL
CznN2lYNGD8ty+TFWYvSLW71mYECJV4OAjq7gfmOcRfWPz1KDRwihXjNtKPOcOVHPIX9KQ+G46eG
gz4A7MHo0a6t/eQdguR4HJ2zF4Y8XUoQTvln8RFPHIuWajLTiXXQnOqWUIzM8TbR+5vgxWECyjFM
myGykapyaALrwnLvGU5FMNZemt/KcdsLZN7vh44nm8++fs1J9Zn9qiCVgX3WxIQ9DoS9IAQC0hyL
tyFHSltbT3j2psO38MMhxN0Z27l00LPvQAiXTYNDhbq2xc8RfZkgveb4GSigYvYc/NdkKsK3G930
/Oq0WgKtNMhRRTpHa4hcmAkgbOM7a8/4lVzqZSZ+K4bilFwp+y3SSAwl4zo7QuHSC4FKwgP7j5ls
SZDYKWQ/iOiLbgBiNsnyK+L+ZT050kRn7S/i/ugcIMYxFvykXUPx9O94W+l9YDli4PuVoi8agKwW
85ZQqigJtMNRfBY4Pium6tgLrfymBlWVG11kZE/UEkOOVtKTW4rC/B6zLwJ+bZXFqZsUiei4/w4y
50bG92IZcUhntpZDWXfjWNAcaF7qWYxc5SjIRN1je4hgB2w2SETIHPEnQQgKtWUSeCGCVdqzISNt
q7kOsWcu1W1D4uceRpeGpxitakiwdrHk5nkOAKpEGItssKWGhmBEvLexp4VvHOu36IKVOoKl6uIe
IBFWnouf6C/+mB+ohSQcCDnCOSGUFkxtvp2IU7OtjY9eC739R9j6samO+TtD+w+ZP8slnur/GHpW
l2wOt+6q6CKfWj5SNVA+AbF9+eLQ10kgL7puRr8hrpcCEvxugVRu8snVXNJZkaX1pBK6CAdTSkB4
OJVHlI53oCSZ0hI+Btpo1Xu1Iw9n0ypKUsTIaPgSssVmNg6CGrToXKrfZJEOOMSYA9wol7talykF
fh+wZOk9bLxLBBeuvlqYVD5HC1VZkOeWqMCzGFw1HiEIGSqbA7U6SkGUPLcOqDQ5V4N16G/Z2PDg
1rvpBq3doL2osTxDKAJknDhVUnVWvMN1faQUSOO3/xmMy//889IAzmRDGGH73IaNJwWSGV7DdNx6
nLM763HCJWwxRiSSmMd8egyQiLJnfdtK3P82Yp3ioT+yWBglEGz3rtJSfBNHKUnvpP2gXpzD+kq7
1eIqbAVKORaGJQfkPF0vJ9c6mjS412LTr9k30G1qxUni16cvgJJ657LuM7duASnre5BtJMFmPwC3
jrj26NCjajtEsKVrI2pA1EGbD/ROtkxG6XaLbdi9BJ2oeftIPi5dk9jVy5v6uIth0vTvRfmbLFo0
G2qjwIxE2J54wCc/tKJ0LXGsoTmRAuJ0/MM0toyhnBJz+GpJ+eaTSO+0e7XUVl9y8V8gIEwRWJzz
JHacJcwFB5YxTxIRfdLTgAI/cO0fbuejUcg4oG54wWiNyhV3+h+wdS8u8HJH5+hcWgVJMadkp0SD
Z9mFV1Eb68NC29bXoAbQqzqeLnw70/QOfDSsdMEp0pkair4uKV/sF9Q32XqW8wdOIeNz9OdKozrd
Dxdxl9MdncASStB0+B6EhoBwUe9HpsTOpEJkz+UrpYj3/3zUUSFATwyDTvt1t49bP84PuA0yYjY5
0BkN7Vf+S8o9AeqsiKMimzpkmFHvpaIdBqleA3Hy7k5R8VZPVACfBkGFPSKKQ1uCkc7Hq0THuksj
TCY7V3xlhkGAkLbzx5bN35PO03z5gjy+XYR5thLO4svfEOavjh8GT90pMI3j5Yi3k8r1XGr9/JUv
LQ2IG1e1DrG5HHq3of71i+t1MhLoxawd01uPky7I5mDy+H8hx/Tm6tFPQA4b6h3WO5ek26sowYLX
6SOGWLs6Ma6Nv+lMme2tDMzWiBYgqVSwl/7DumbJamdy0yk7+3Ay7INQAByXf3HqPGpqjR8/7QQb
94/YHKIwFNQ0h1ukDRBdBwxGKeckQzAmjMKt9ESwowIGBZKmt8b7xy1Ye5v51Paa3QFCX5rQjxkh
MbVLQ/+xHBvVlqmWVBIkBm4+HZC+VxlcOoW8IxDcpXZXbZVpuF1vquokI0p0/F1hxP3+78zqe0f5
Y2B2JbeifPFBvyDGCSjI9Pg9Xa/RtADdxXjCYxrOQbBzb5TD0/3elZ66dFUoQIgCM9POgC2PyFpK
g793OvVoMpET+Bc0CCJeKY/Gcco3rpQz8/kUYs7Hmdp4quyn9Pp5F2+89G9/CzozuqbUtdIPfztQ
e4vFMl0E7XKu92NQ7IISQ4Vfioo3+HSj5KqpauYrbQYonJx1L9nv7kuaQc+JBusPyYfa/6A2x2sZ
I3WdWFqyln+Rb+I+dEhnYIY5WYWv8TafzPS0fbghaEbtzwqDhGdlssbYJuYjUKH0scjzU9Rnj0Wj
OCWi2jM+zzmf/x8llqrXuDwzjiNnwSwMzPVqjsX9E205vOVUoeH8oMcnb/zrWqkJA9h87TKxcAqv
4My/uyP7a5zr5wj/6DBS4mYUTE3vWaEpIlY7w1sFS+jwg9oV3XPBarWse1BdkdEPmwPmUTVTFNiw
3mM9D+fwX7h7djqUh7p4gRcsWSrwFwjISVRIC9CCeJnjuC+BOwM1SCKjpJ/Nr57XAsxwFx/xStQS
vZyHr2uGRvU1DiJxxGzsVN+52opTQyCEO5+crdgXgPnpNFR13kINQxR1R5zJpoeNJR4CelzVFTM4
+NsonzM2a2S5lWn9LJeLmGIPQ+24qxLLfdkorAMiE6wyGqEh3DgNs66u7cpjdCxyj/JMGn0E/XR/
uN2jWX7qZdGUOPESeu96h5MfeaJV45A65pW5NsreHbcc9pVrwYsgQoH3jf/QKRpBoqJ3LQtmuDYo
hTLicqKTLzjxVKSLgayNiztQdljuKRxL23mMmqK+VkWUvtVxy5wDhiZqG6d2PtX1889zNw8guf/e
NE1oav7H4tdkHWijqvm0lc8rByDC6EW6eiRxBDLKtxL96TuGbec8VINrSeT+CIBtRjVw54xBwAdE
TCNLFJXYMI0MDK/VpCH1fP6eczm9Cz5Nj6t5Q3uZEu7j1RXMN0LIOpX/NuwjednYGIauP2aOkJVs
/OuKB6lxY0Y4X0MzykmlxyGD8VZiX5Un97yG8z0zNIihuqjHuVId/gYVlKZOLOMrG7ppB7yc4KgM
bQDoNzizPZEIUZ38Se7yZsbfCqsbzWGs8NV9yp6w5FCp39h3G+ks6WKPsOjlEx/+I7VlpG2t0OOu
4Bju9zC/ADbczDjYAGQEhvz1PhQcfL7002wXiwfPIxS+cHPdQT8Brat6UsVdIgK72zfHUHbKWO9x
zrLJEV0FdiI+5ovvWIbYzViDCXJlXv5hf/THJqBM4FqzYr4poLOuUBcPFFfCz8efBdz0iYQR3irU
exGpIC8+3wQCa3cdqqOixiX6TwmguRlPRM31WiGnt4xCe9VqyWrMbo136jitdD+6tGnUezDiheVQ
S+uJT4DpbtFbCWbgRYlUjwWx11UuBD3UiPWTRnfETdYV3BYrNL9QmhNBXp/D6j+E4d/W/Ik3Idxw
+2Uzu7Ya9nGsfqu8ifSwUycHcL50a2Br0c1XzsEObcOQY2kw4+EHLwCuMmmhRLoIJlo9ilCNWbSH
ehSurrEr7ox48JRGqhPhfaW0V1LV9LFyAbV/7lbzzKd5utfBzs0Lu9WfwoP/00ZpDHYeszgGzj1U
RL6rj5Twa/57j/44CN2UnTgeo5HfZumQBPyrrmYYuK5I0CR4fmkKS335rFd7bmfedEZhqhA7ZfP5
Jyr7ueTVLtETpi2/OzY8tUUKEMY/1DXzorKpbeFaEOvJIXgwg5d+smt/9z8i8FSWA6YVwo60eEGV
Jz5lolUSd++DKWXKn1xqXAK/Mts4K6l1N+wOfw9Pl9b9Tc+lU0X/PgUvTD8B0tKKc1FLt57kdpbK
4X06unWzPRk+aZi/quEVs0xpSrVFOVPoa0AUwXWyE0HRogKV6t885gUBtd3XUgczC9NMe5yBzgMd
nQF9Tkcjv6VlUCi+IZkr8Q86SZNI472evEQAXNz8sW2OF7kL+ARwVzmLMLtKoMKryoyuVbRm2tSM
nt4zjHTaUhA46dVzc+rFTMM4hK3ARvbKYw7coulJp0LabGPGHQuGxVVfX75kS3tDNB7Udf7YWV2E
ShnPTgiS0690kC1OGmDy8+XPih7fIHuCEqI2pNk0XdsPSHauilq8DUtkYu+DQpZwY/EGGD1s9J+J
AkqkIZjAQu54RiobzmeLj19+A9Q/99nOSpannI3OzLGp7vVKUWQETCSMb0ZtZBM1pt0RVhLQIlTm
W6CTXEX169NzoGXny2CGyEtBuwboCcWd12nJUdEj0WXCeCrszOsMSeOWzM0hcN99JExmKEBiGGL2
Xwm/AhW8Sg5C6SDkA1VVTI4CTWHi6v0RGEz9LksCVizVO37TviBWjWUVHMLA5m6iULcPNbWrffTq
UyHbQjMfaGr2xurK0eoteISshJrBSVNc0iw1Tx3xZEe6ylrRRRtEypnfFcfcTSMBUTpwuSkDwggu
3CQbLRvt0maJ9YaFjyp+KbaMkpf5u0dMVx9D0Z5E0SoGWlYCCLxcADhGhz5bPYaAu/aT0dVJ78yg
zg4xvkGizjvJrezN7yizqSOx45g1ZxpYqeHiqXD2HNmNqQAtUcU2REVd2Kb0QVRR8sk1dZNrrXs2
s+JGYXjGLiMmgOTOjIHFE8XAuTWJJ8oa492LoVaIDUNCXKH68hthWPGoKX5nMFUhDh0+ewoMYm4d
DTLdsdkzAjl9SesC7vJJ8YRzzaHFLxbhfmbpLQvK7fQCwlCYU57+fqdUkzMWLmKAKEybpPjJUSPy
z8cq2ha2IJlHojB2hJ+aQlPb8ITn1P24kTY/pVgJcmHb4+HUWYw2cYqLMJcE+w9gMSno1/jPVqN1
4DW0LCSfGV6I7F5+TbsJOrVO8ZtN5Sc3hBhD1TuFJzsfqfjYz1Gd27f8LRn03HRfUZKCC4RYp8oB
VfcupreOAbMzJ5eSV4KTiCYBOiy8oyOBkYJ7Uk9u0DIyIn76kkfa9DL1mS6lTxopqPqMoTej9L6j
FETkqHfXO+hXyT68MXcN6chLqbPxqDmfrwb2lFfZEmydlCL1IrKYbNt5tNhHpMj6fwDC7ROTz6qO
otXj9Gkg+R2hL5iiMdiOGFHb0jEJt3cawkcP12ks0VK75LiP8+IRGJFLBLJXGR7OSojBbAt6rqdZ
Hi6TAdldoAUPI1WolS79TH4LfpG4GD66YPEpFb1WJIspn8l1MffPzC8tqKSasjmmX+iRVqlS0cZF
6VViNbcwlhSlv2FdJT5sVzvPH1GdcXFh5/pMLRqoJhwj4RWx2vOBmTSdEsnMXe/Od3bBRpzJMxQa
UWgdEKZEzPnIiJ95e2GiCRiJ3q7fh3rnzlg+U6IiOSOOGdLa1g68Bos5QVYVmAdB3vJgkFautYVe
sM+2u4pzdf047nPLOJAeg1Qok1sY4zWPnLR0AfULuBN/YUOfalw6IdezScoL43d0qnuRem9MusQl
300uMlAOO8fLS57kuQ/CiFrpbsuNSke/TcvWRBP7w9LAyd+/SiDx5NHwZ0W9VDjyYBPsWK3j4VOT
TpUI9nw82kEvSSatjQwcwQVJ8CtiZmc6xlxNxWEcShkntgMtYBEX5gBjRvEn6bP1NwWhBywcXok0
87eZpkt684jYCt45k+zNEEEAV2DDTdBNp8IwjUCpb9KywxiUVM8d6kx0ghYLsAu9ctl1r9D5+WIm
OYmww+aIuvq57RjI+Kb5DVPJmdTgf5ak+h+liHph/MwcZFXMM+cS1x/CZiVYnZj37tJKXhLwAHKj
KmnfMvKXctbJFINBK5PsE5Z0EKHSLEeRxbthYGf2k1e/mIY8Tix8IRktHsM/kvg4/XqXJvmXTKTE
g5rC7j1E7TwyNCPNz6SDy3P3+eRaM3ipWUzxPYaOOp+0aWz2WKnSC0DdY9P3zXNDYJ3NuJxZhxKB
n+PeEj5GchTxenZQZK9/nM9A+dyua+aC8cIbxyTuJKFQzZEYoIHeodwQUPt+qoE5uTWrSLVFmXYj
J0CB3RgFQLmmosOchJDBtNQKP57TN/IV3RV5pAqWMlTl2GhR4e66la6bgLP4wxoTLOlqddtVvXuI
kxkZa1/2yp5JakRhcx7FgbT/kpdeD9DuEAV26ta+Wb6n0K9RVn6hIJNyv0KF4lutGgjn/4//aAra
adEEwBkpzyUql9orhRLcg23sFk34u+MKNF5cmewXyJ6ZYDZO7zPwkd4I34fRoiYwfskondAYXOei
lrCgBg4AGqRY0TTXlNIk4QdSpxnjvXTv1TGjHBmTg7wmn4C1U32LQ10RujVU2uj++gcD7nxnuA6r
fBCs46DjewyYxbQgTdedg1G4PR+7EEVIaSPCGqI/Y5oBTO1UQLW9vhW3fNMtczb3kVMNQp43S8Ij
3prCKQ4o7UU5Jrkc9xCZvmXgsvZMHSiNGADMwegZRSz99dnOfRYoUvoFVDye8e/xOJ77srnwawku
T4KJvqOYn8w901sC/W/K08nNf0KT592Xy55/GM2kjkXCfA69zeNVuyQTKy/TFbgj7BF01tQutpFJ
TpEfuJBN63irDXdXdbmVybTLXpiqrKXpSfKTaHjMhkZqV/hBRvLsBo6tKHO0xKKfKMdLpOtvyUmI
CLp91OM/9iKQVmYKX8vfBSv6AK5DNh9bhmGIQ/J1R4c7q25O3E8/X6xjScGrtNKiy1m4gHYbofHF
+c3eixVUt6jHArHlQYZNXY+juQr9S2OHnZRTyR8+FKJ7nQ/UoMlqiP6bDFUdEM5sZNioZz5E6q7S
RRjbrTxiR0cJZtdwMcMU6ymLy10CA1ntXiERCYltRFX7bADdGPTby+J85utlpDRVCpTwLZPHoJEn
pIFUhthEqfiJeQM/z64wrxhRP2stATGjhFOTpRtv+7fnnB4DKSLomS8RwfQBOIPy2+9Z3PFJlSoj
dXjB0GJ52IqTPFgSRmhb/YjaBF5Fq/2ZPr6fvetuQrq0v+6B6OzK2UkpKvY3vhImeniNdDeAizwn
Y3rAFtxYYsutrhNg1hF+fIdYx3iiKvIzb0ojTfXknXh8F1Nj86Y8bfyUg5DoC60E8RGOcC+KL7sO
F52zCCaYVp/+maE+VoB6CGMOA2+avXQKEgft2/n9aLC3tyfHf6szpLXwWjyfSHAJ/0ZDRY6Ni1b+
f50trzaQyeQRvdWoPCRpfSCXZghaC99XHSettwwlD09qrZlEUseR5RCCRB0ZdYlvrGAVWyS6bhsH
CjeyCvhOvUo+6x+eEGsmRpVFBMKAqpnL/TaBYiccpOvwIjM5m3Dh9wOEnOT5GMWlJhJ86/FwrlXL
BDdOoVhlPvSlbn3RYTE1bugVamothlaxabrDO3xIpDPrDfnZ6TOtUSOyulT49acGUdyr0j+izZCC
qfyJDBY7N2bfTMsTmxOxOCAk0mnmRUlH7ygjVal4CeBPwHyqPOY0dBic6GJ6vMtnhTFzVysbbs1F
60FHyQZM95nInmDO2lihjZ6ZdDAKFmmorqxQhkkV9e0RPof/lJWrs/t3G7UMLGcipz1XQFy0H3p/
+9dhXim+dYpBKvXCWhalXwffOePhuAZy2bjtonVeneqjhCAe8vg1U1shM+Z2mJS9z7H+AwirRL/I
WcWM/fQ8rrRLi9vMzhgny9vIXmVrrzzob4AM0aGaseminowjf0qwJWFueMqHfz1Z8Z6NjFhKZrRx
T2169Dx9aPr81hBpJBoG2NnKa6UpcAaQrC8j8B/fHN8FR14ncVXhmSmAG69gRNSI64eZrq0hGiRi
Uw9DlN+7i998G7ljJeRgTv41Z0VEF2AgH7oEDH3t5ic4jxl0HmeHfWX3mAGKRAiZzEqLLGHYHNXA
xEV1gNs6JKTs16sfU2cqDTOQRRBh7wvUMx5TexTFFqIT4BqhIvvnzxyHtpwG3zJzRa2SKwfzdU7M
Sp/31IwrV0YsIc7KMF4T4zgbt2OZmrZDMV9fRnLv1TmY+2dFZ02ibEMv8QZMYRhkdl9Q7+gmNkQy
4Np1DZ/uZEVKGRE+Wf+lcLsnuqIq7SbqXWNLxCwf0J6wIfkDyqzOBZfC0Y2Pn8cEZ05mSQg6kmMB
W99CZmrpLmn0MkeAcIKGKcc/ZynAvLmxg4wl7bhVljUpjwzy6hwcoHZCDRfW1wRnXsuBuJ67w55y
oL8VemOKEozZ5YUr2HBKgsLWDTuioOB3FMKKJqM9jybsgF0NEVgGbjrcu5VfVt86X1q3z/gYQu1Q
dzZALm2k+IkyUFC75bQQCO5Egg1epgsNPbe9JhAdVA7wiWj+NNQ7Yq8kvO5hLWyTp59EDWXjsr74
A+GzujLNR59jKqGBR2IsPIsjHBVvTXlDIQQrMVRlV5408AW16GSAbFaSWPGQ+iAILJidqB/f/Yqa
kfbOl1e6JBy13dabjdW0r8Kfz4LgY/shXnpUhh90S8eRYY+G0SBI5hgWqxm0JjzFvlKVG+ZBDwh5
WzqIpHGZ6jMytN53YfWHPaaeniuy8xDNt/EvJ+kSz12LfzW2z2sTYXRsTO5OPyX2fsjUJhgMeRHC
G9j0jGYCGSRvFlbYYS1nIWH0IzeN0VJUnA41E+DI68w+Qe1Gm5Z6Jf7+MZNI3M4cvS2ztMUstf4G
fqb5oWVZC0qdd0CJoABn8cji8wy+HQSMsZViT3fjP1F+Ys/5HRhGbBz1rB9IPFZlv5fVYEVdVw6w
ESOKwZDmd7D0I2SwplUpU29PeNJiqniG1vS1xYg+PkG0VT28mNx+JtYsQZqBvquXqH/ztfIxWV0Q
H1SHcZGT8ey45HuU6fk6R8Dg/DCD/3ht/uAUPCsOdqC+FRTBlEKz3M1DJLZ64Erie3j1lHuwzsMX
jpwDo9d6AHiVjekEJk777GIQE9wslyocPPyu91X7LmVixgwK/aIYblc+D17czWORHnR/rjkjORUn
5Xb9+E93kXBCumJAManINVQVCkuA398oTk9UsQ72hb4jCsQIpVs8H2EQ9FE+M7hni0exvKamO8GU
TR9GYIKdSQQO2AHnrewKdEXQZRqEfWO/apkrOB4R5vMb5x9RrGfcNrZwotCxPO1ha4e/8OcKnfX4
J0BH/VvxOup/qyNNxyW9QfE3lsQOvpWZjFhY79zUd46fQNtkTexMa20R9i7DLSdAPBDDobY2ogG9
ZUvB0ligPrY/fNUmXp/doWfpahaZicRBptXyKLpdCzFSptW8xUST4qNI6eAgJWf/UfbuPa/VlgCW
Jnma6qt6uyCP+jdInBoW2bIjaBDwLi4GJN4HrzC0fVeGHyNMV186vFjda+4IEljhnHCdatVOLfYE
RFl/uR+wdGxKEJzjhPPgExFBXgxfQsl6nBZ4F86bPDHDdJMtpIhJfX5bgxR3l7/uCt5HiXAXg8vy
SFJfv76lAVAbiURMg5qMUHH5AS+Xzx/aKoHg2zEEDr6SM7zzl1ULlWB3h5Fw4SmxdwgoutcIfiyR
Kdx33MAzXk+cuudAnieHnsAuipP2m1ICkB1TTepSL/mIrK4+htAQWZCFRIqTe+FnhscCe2+DTbFH
9B58f/skcvLKE370jBwTmas+8SDL38KsJdwpdhzt5jguE1lun/DTTSZw/btr0raryae4/891Gwxt
2Sjfe+Y+IdnwHrdpm9gsSOzUefZESGO3/j/sGdeFWnw+koPWpOOqTPQVTI60JxFwNDhnYX9eFye0
AVOd3X+e3CZLs5tzUNgnDShtUfHgHGCrvufi5/BAQC6k+aJlPn/0y+fZDO6ODq2QFbGmx5sAYNRz
4weRBzJnWY8ts0AUEH8qRECJpzY6NJBsJTNb29vscYZKiewopJBEyNLGdVTqEcPe3uBjPjjbP8DJ
HctG/l8OyFabWm/dnJrESbm91pyi02LvuQtfl94OwTI4eWXnpWI3JxOkq2H2A19NeCDriFXoH62B
Degs4XOhtvSQAkNNwZw9SMxfb3NfxYJx+36UrkYKDuRppCxh3pT1p1z7jveo5xrPpYp9qzbnXSpy
VFch+EOBfy8Dj0rdbVkSeDZ4y61A21wYKRsvB1DzC1fiN5dWjrrAZNlW7jzGQnRwWx9cANFe0H7u
EgJoUYfZxuMafK43t54Lm2UMEXtyyfravcjD6HUOozpcBPjb/CB1mLKHuqjrgubp9BYo8c9f88h6
/3hrvSW1eGURoc2/ApmTIUSBBoqDbPIq3BFFmqhpGsM2O8ielJPeP9jGlBfspyC1JusqE6K/MRHN
SbiiZ8TpJ8UYHQMwBRI4PEtfJqDdLbYb7UYg3afZj/lCpOCSwHTEFDodW4EZfVX9yHyQvjxC6kBT
AwBfZUzG3kfl+Bnw90sXEdN7rUY5bZ6MCwM7aJ5tjPPz4NOKO5qVqATxLtiqY9ERnVUWy3Mb09TL
g27VFrijavXcqCI0Ldr9WkcP041RqdjKsgq3zrw6bcXnw0M/NxAAX+/NxpMOsT6mVFW6CuZ2Tr/5
Occ/M/AGTb0orGhmH8w6Ds5uoK3QwAJuBMjFCSzLbq2C1c0xRF0LTx8SBu8bDwMslYrHVdwXYK3o
saXGmpifejY9TD4gkz8t2JdiaRC5D93vyVmaiMQ5hf2YWXOylQiTrzMXm4uRHrIEBvrgI0OIKGDK
gQXXLupX4zh3Axr72bwNrfIr2dgEAw57jkwNC/ngNfrewpgswa0bW4H9XrPGKnQltL0Z1jozhqzk
+nx73W2YpheSERDtkY/u2xN96+AnMIIsQ7gGHYteyqDYKVjIRDgj9zwlvAdDaEBh5cS7T2TsEacz
0SjI+gSHB8bSNo257hLTKwiZPevnPll1prZMgkvAoT5dR2met/LzBNxwwRlZDpqhN7pdsVl+e0jo
c5JyQnyokS9ONWZXIBJFncGQgJCo3goCcca8RZ+1/EVq6YTiUOYZbrlX+rjx1Bia1EWJ0VQeP5jL
Poi4Kjrm78vHNhE5nELrfLzzpq97pTL+49/jnGUUUoVG6Fluk38RuZpvzhDL4EeH8Lb+F3jKGzG3
Y1H9UduNHrnCEoFz9A7MXolLSjWEMSPcpPTGbOeORb2J6B3z+b5u250xRbYZwEbcqS9jS2vguNpP
CcVBQ+F5pYmJGodTHKqIYoSo7YgIlA1zTJNxKQh90ytcgJN5+/+6r1S7HdzVONBgVOSu/ydDqK8N
W9X8UbCrX0Bk2hE07lSqbCXOP3w7CikYYyG4YdJVCH1dFGSZAPrDS39ndRDhtdgEmF2LhpNNB4DS
vvwUMtCzGttqyPUWUKZHD4Zy9e8sv39MDaCr8PwSs43XW8KCCjeipYA20xcTCvmTVmPYjVNLqhjl
GuUt28+25bj8ULpm3XaRT30aM5potmvLvOA21ejEm7SBcFnF6VWHOrPaUgKQNlvJsXEb9mAvSksv
t/w2PjZ/JGtI5jrZ5s9J0WAvNBYgcV0fLTH3fgztllI2MWF8SDOotjEYpTe5qDRWcY5SBmfzB7+3
hmXRpPF+4WbGVzYKTm2FliJOrR/d2/G3E/rpXjPyT4fNq0mPs1Re25cduylw89lFj70WSEUi9H22
bp2764xGCr9MwBYNZlUgJfRwIrr7jHxjhZnQd04CXMysleVmFx3bXFUEhtHTI9eNUNIHnbUr+Qrv
ZkKjn5jF/h0N0FrFiUpmCNI6koaj47ncnVpx1yXoPKnvqLAhQF9lOdklsgMbiSJpHxZ1L2Osu4Gk
wj0QIXEyu4ewztGFY2VB4PalZBztGfZpfDItFcxvhB6cKvE3eE6Q0wCuofEsxj2iIi9+13mF1CRQ
iwPLbus+zM/vcSxXnwwfx1t1tHfyyRU+3zmrTtggEDHvDqhbtTCmOaVzMYn1psdyq61AboRXOvfJ
JvdFoa+hSlMqWID/I4TkBFZv6RVRuO3sG3G+A2Pg9uu0n6Yik8L+9CdgzFz88lMpxm8ZrE5UCvA+
jO4Q0oHHCn+Z65enb8i6qEkySigmps2PWYwwtATSm9a7o5FoBBkwGfwazXG8JgHixXHDikA39GO0
ckwvLdOJE4BNhoTdhr5+XQep6IOqZVuOdG/H+wAQLgKVfcluIPxcVz5GuS5t5WAfTdXCLaVTt1LD
WVeN0yqIo8CBfs+XLts/PGbIMHQ7QCXiP2JV+Pg3qNcTiGckpbbz/tpuqg4esx7CK2ByE6usXrkj
ERSFTY5i3inZuYgGC6cSwlcnazHhD9bR/6/2q2RRzBuNShjCXXXXJEFrMZLsC5S50eX+pkRgBFs0
JgbnV+kGqcb5DtrM5YBjASIQpi0j5I6oFDnY207IT1dF7XNTzofnsWN1R38L4C/z4j9Mh+h5Ff6I
2sGfUm1Z3pyjZTaE1eqOXCv4csbdmeVnB4wUBn0G/ATmfS6HF9kmmomPI3omjbCbnDfvGPYXWr8F
Nx7IrbGdJWjchOXywcaRB2Si9CvpIdLIUyvqAECFWVoXsKvdgVoy3i3tzWXwdmJsVFPL3f0ZtKyN
7T5Pvsp3fZkE40vP9UBH6Fpyr5vDKeZKbm/iML4c/qLmxMFIPPX8gEkI7Lw7Wej+8MOdeXAGx0f1
2sby3DMF8ouNzH2mQ+86DTx8SlxirDDBSOBxl3xXP8fr3kEVuyZmGNBzt0UapxZw3XJ30TQZjShu
1rZunzNYIRFK3ViYFfgAaValyMHYiYJwpZvniSjBLpacbxp6BdYbfzlOGaQLruk0fWjM4kb6rUkf
1sdIF2u/r0/ik6n0OnBKmWfibNfKtLd7qKvX4ieUPfXym6MR5mYoIBzikTx2XqRvuIwbL5pd+mFQ
Ukiig61zgjg2wnGl7jZUtO5Abwu6/GtbvsYbj5adIRjk8+zQHjZ0OMd88Wp0P+9AfIntum9LUzX3
GTjlYxD+T76r5oNnD/fOcyzTdJgGK8dRZ0lPKg+7SMyuGfEjGXHDA46Fn0YC5iVHonu/AhXPE4Yk
Hi8ikHS9azyO8Gm/KWiVBi4tS1RS/IIUIXjA5vaW7NcAEQI+Y8p+71bQP9/cgCTb1VpufRpCTFWG
RQbH/oU+Oi2e5CNk3tOatfGPC180sAsTm8cGTjDjSeiCcrRRuGkd9WlclPiS56vBwh2OHFE79PZH
xBJAphDTaC2BWv3CsZgSq/rbIy53aySzf5/8r4cSKAbiyFtoChJ2/7eUgz/01/ZLxV5N1qgGpvrF
tArLSrVKqSI/somMcZyLo79lf+UGjlHWGmEZq5gKYktJS1B6tZ3e1rsPBBQGDfnMElLZT/dkja6X
kEZ8WyOIh5/jG0OYNfQ1p7wE7FqA2c8lyzu+lp7ratLHhTkF0HX7kWLPh5o9TDvbVncAp5VWVIJf
ALl0qvSIbxJxYkfyeBl4TmHuDyTh4BcZ0wG/thbB5wFp4n0QJhqRpGA33JOSHwQXpEgZ2wvSUZHy
jRAu+yZT7UGex1OfkzIKMpAr/+C/ixFWq+0oxqd4mcuwNlAZtdf54BCuft1f7Vhk1HOb5VQsM4l7
KRG2ZdWwOuGdwX7ApejEgdJenBdIqg/fK8H6w5ZQCvEn2tipJH/2IplhmsHoPILJno3usbxwkYqk
qQYWtpOhhcldldsKAxkgWQS1s9Gz2SBmGjXbWZ1dnRCHKVxCcamDEgV/EYidJYa05SmXC+uCwPqa
QN+n3r5C8jHHoWvOOPh+2aOPcoSyA/iYKGg68vVu+JXnH9mRZpBy2/AiO9g8ycdgeVXc+VyLn5L9
PWTTr/goOCjx0HVWri2tZRxcmz2v91zlONtrWc9CgzANMl/bUPPfoTCIS8KZnct0FfbUWrFcdVlc
3s1G4HiL3D1VIa98gYsj81mvhuNWf46+mRAH8ke2A2EWGlSz6Jj7VUPspCwQmTZ6ndPyO9pHpQAk
If9e5XfLwAITHdea9zrte78HEU09n0t+VJA/TbJMcABh91lFkQAteiL+nU8KYMH2ZJmwb4giNg+K
dB9G3izq0zokHLi8D/19Jh5dsj3HYA2w7JbX81jdWm3zcTBHPuQYRtiVSEfyIzhBOPDtlt6Jp/d7
/AdJqLPbcOiiI1mpzrHRiW/TBiejWR4+6yTIbaJUDWiDEZV6gN4/jIQvMx12JOWJeCrmJVK8HVHv
MJh8k5i/WPUofdMlbXzI94Wvz+BiRe9jl89HCQFVrJSdb7FeA3jqdpcQdai8qlqy6u6rQdXRObJA
JBo8y7RQLhBaOlsYDWtzGzB/wMaWp1LnnzvYQDQ7v0wc6HKYLkJGNxvQQ7MGfcfNEHYg3CFq6HgJ
3DnXT6UhQtW9Oozr9M5VVqs5FgewN+fSiXuVUgaeWv3AoDFFnLkOmDxljuiKGMX7j2kRpoz2Cfl8
PV/Ydupm1C3oDsnnfAGrVbTu7LVvFQD1RMMyCHnjh7mhWMABu7LdjGu614tK7a8HSISODG9G0MSP
vOQ7564boJOzyb5kblURve9W37NzeMFm21tv5e7Q3xwqc3jJ1lCSb3vSVp44eOah1vPcmnmbUnZR
dNxkXM1RuMONnp2ue+oFYDoXGeITbVBBDyzix9hMeid+xWardG7+MS+bBPlCF4IoRXG0W1tEIWGl
SwNWzDBy3JRaXKDGDBjkCUemLvBbTfSryjlP/VWP+gKucmL6BE8RSNs28Zx+Dez/+PfMjlgwrMrU
XyCuOOt3OjKAXd3NMRpbPURgUlDzc27YTLJer/sbO/O/9PpcEU8fd6AVD4OhU7e49mskZBJDTwyM
LQ0jE90JuXFc3OTsW7cjRfIiTUKqpaIoj0wHun5hGNUX8OEaf+rToQJbSUnUgcEMbT5n42xQIvlM
dnvwBYC6YQS/UX2ZYACpGCy16jIr9hc/hLu0d6cbV1Z6ag/B/h++ceu9IW9N4ZZldueqCmGAWTI4
6vQtvvGOSgZkECZnhY46NghZGjqBlIsDDqkkhw/eKFN+w2hPoyqV9NEJ2XdFl1aV1+01epChwmo3
3q/FkHwUxPzLPYgRs2NpKrg6KAbK2le5wVWN6tIuZtliZLbxBZAkLGvF2dkYEKI3QEQeATUn+rwG
nehI1C07c7YRkTfRsWF/L5Lw0sflOA5V8Nm8eI3mzC1QwhvMxv50Okkxqt5dsri+TZS/fnaqbbUj
CZTwB1teYe+GF4eeKV54s1WcI35WD2vM0hG9ikCpa2L0bDufb+20Hqh/6NLLFrTZZ9Zp1uQIX3d8
n7235Ic//Fp72vWbX7bm5oRMEELsp4aeBg2kZA7npKIiUs8hQuvJlE68VSnVyC1N4wQwQ0BT3LGD
w1coDbbCf4VnL9hS1j4aIhQO23S1D78D+RWkfrQcnnZdGTG2uhYCjt2VPchjsTS0r+/ezbPjM5uh
ezDlZBq6jjsd/3+OfEnHVjPvzur7d5QseK+xMrNLqzFEzXcio64sK5qfWu/msy62PfzeIp4C4566
2aGluKnMEUtgdeBpTuujc6B8eXiEvqMf/nF+t0zDvwRFVNk7cWwS3rUTyXAq//jBOgUwlsqPy5EX
oGl580jEz6GFndOD/CWWQ/DWrKe5lDNT+eWsgj1qvpr68X3zm6fU0lTJZw17nf2WQsmf7Nr0Ihe/
BklxABZISHJFzvUXrlu1cj85xKiv1ZBjcAMS4hGVYS4/999olRwxE6eNoNs2vT0t2ft9+mVBGOle
ZAUUch4Oguo3ofcLqbi2PfgDDKiV80SNOtpBG3vzI6SXHwq0ddjgKmcmoqfLTiNR+jtHoVUdGanD
zA5WIL+bo540x51fFNPy8X5LG57BcdlMLLHNslummeRJ2jKL7Ir9HL6A0JOXLnH3fF5ZApYLNQAn
6hJd0geJSRggQhqEf54bpsoudl0MhMopGSgeWFde2T67niZyavfxQ3vDkIgZoKSn0if7m3JK++H1
89v55+YsY1W3gzbiuVF5j3NtG8PyDxpXrr3YHdmuuiDuFfa5UGj16FVkNjJzcrC8GzUFqF6H6PJD
Q5DIQDRrb33CDRNVyXXqdHeMmu4uUEFi6VyryPiwVC6/ycN3VascV8nh6fCnGYT3CQV6xvyMTBPQ
qQ5YJqPSsuwSE4msVSzp1ooHdMIqzWRX8OISH8QyqYQ8GqaP9wy6T+NEiJSMw0s26WTa7pCw/FRe
buqPJzN566Xwp+D6ajrNW4OEktXEYhSUhGpOM3yImO0tc/M1bI4YTZqNZ6mSnHxzgF0pzdBtsq7z
qjpvWSCyxJUYUvX7UyT87YcqX51cIFe8y7HeCxspSVZx7YY0vRvfzuotksXV1b0cttrtHpHf7Ep8
3Ifnba1tUN7eOV7QdXHUyJzcyqkkL0bPdcUlO0tBZoPXeydY6PNZYeiilgkwjNJYa2Pw/+vgI07F
E9tp4hgL5sMP021Cb8Q21beI3Qi3pEkn4smMaOrCqKlJTZMTFZiNQ71q7nTPC1+cOf2vpyjFF036
KsYQhs4WwjFd4GfmP5GKmH2HBLHGsSlX8a8XmbwrHfe3uXvMj/x98SPxqhVBQkiMjhIKYhsWHohc
T1LD0MCn4qHGBSmNSWN6zi4krLGixgSomxjtR2tNismtWNwmb25SdBVePO/df+eCrQP9QuOjJkwm
ok6k2gdoq4hG4x2iculGf/+E5xouE/eXT2GrgeuSjxr3p7VusxOONfTrkWDiFomQbJG9bpKKGHIh
LGrZofv+fFZyw04B2nOGzllWzLeKH8MMU6crS0QLy32BCLaeAdvwaKSCxpB3pz/Ij9hj5iX835ws
uCLshrMl6YPRFgncavhfQV4vyzYyGnRpyZsNEPyauXADBz2FLjs7b5jjJWiN4Rs98T2Q8n4cgYPu
b/bvtbdp8RDaLxHczf2kSDqTbyr77WVn8nwoNpIUIn88k+nN/g3Vy3wY/XMZGRBpjVv2Gj7G3C+Z
DOA1aDIJsR8hqQIdPw3OKaxaHYkRiDgB9NF/Wz7kj6oJTkc1cvN9hNjOb3c3U9eM/6BgYmMdKMkR
FC6HodULEuNnb6xc9jlUt/U6vKku6gM34O5McEkVUpY6sYhmk8XRtl8ogs0CxW8FJa7BRTIQvWgz
cCi0RHY0nL15G/IT5UcRXMRn/fwq+mH5zt/hDEQePzgtO5v7jwkrZ+YDBL5ZxiY2RqdHVoTEhwiz
VI7dQdQ8EgDKpp96zIhFCTFsYe5UPNV0dDuS+Lo67td9Bt7QGhA9YDQHo+xu8xYxeqzkOlFw8qXY
Wkmxlagdt+todTPqz1dpJzWWsfzTxXWHq/Vq2WoUf89zz/dOwc93pimChY3bv4y70qhWFzImswLv
Ou7Y7icTCMVfyzZHHVsKunQ2kleHu/3YTr2kBK0u7slAzlmHC9fUciUayIkNGIXlj9s/W89SK3PV
FQNkVtMxY4GqZcko4YWaCpxAkwDXYWnPT3PSqJyihnQtb8j2d+HhdHaiU7XlmeY5ZiV+e4jWVgsh
u8DSAo/Ms9sBYaaJLMlCfcrBXO3ukjMqPgjZEQlHGyDR0iHY9hm0JXF7UcDPvQF+dk1zHVfEGr4I
/9Tu95rReht3bGbJhFM4xWoJZ/qzciSqbmtyLC6R/KOu/rnTpL+1mJiWd02BInlUDAB3mQnZeXGj
1dNi1/XyGq7NQG8oRRy4Ci09ydIZJ0pjXQA8bS3b+UYLcvModkwt8rX+k9QlClf2b35tG1SSQsSy
0XDfd8URf2tnQeZjhYIZ6zDV9osmetZuofc8oOjR6lmtxzrBN0o1qlRoQ1cFNwSqbFRHN8m2bmqb
v77deuRh3aI9QBK7+gRus+y+tpSnCGdqf+q+t05OkO+x0nQZ4NlY/8B7FqiGUBNfbdeGF9YfxvWJ
rFEDkHFM9Y+F5XTZ8lbi0a1tt6iATXGjCxwenZyGfnzSfWjd1CCpYB6Tfrbr/xC5SaKVHBRu1g2W
udZgWgYYohBXFjdj85/SpPfTp3Ni1JseifnRhfhwKpEzhksLAiJpgZeLZp6B+FRGtwTjnFO+GzMG
YTEzjHD8nH9/zEQqibp/Z4twimW+GXznhKpHhGaKRvfmmx/rbIU5a7KQnrQqAmC9Y/TtHa89Qcnv
/3ukDl3mwjbkXI+WNj6OXBv2kYE74PtXk6vHC4Yp09uKU3TtNBtBpg55g3UpyIqhkB7Py2HehuCr
gWnmVUMtfgE9sUEA1s8+LjI2Su6vMgGqqhB22BjJ5GX2G8LKmwkozTTylhMy8DyUcsyMo1QGECnX
GfOiQVccRFsT3k97zvGpfoWQvpAtgBfLSSfTbkUFtbFpCY64C2u3AKDOgxqU2L2U1plcFMuQeVpL
dlsnj/c1cihGJhHSTIgbxEBEYmMvud+2+m5eo29401TyYd6rRvcZd1JNeuk8LoXLV2epKBWPVi8z
1wREEAhGKe+FCCguwhVRPlbfBNJ8QVTdIOugxD1romWZWHaThRYZYoucO3IrS4K/fsIuZuhkSPxr
I99hNb8NYYR1uZLf4yoZR6UBBW0iS9mS2kjCiOShayN5jaQJfxtiVzbCPj404n5SQThYoPjIxrSv
QKnBHK6X5WhVMpZcaXDO6zCUaawIePsJczNLdKXov3KmtYcc/YJyvGryu7kC0phkCE29LBfWPXl+
FQXTKIosvlGWm9TBhrnHg4sakI0bruDer3ISV2FZJOHOAR4jX7HWuJRb79K07n0ACc2nUB34aIaT
KIrJ8PMDJAVCPua5Km7UPPrHHdyIHHhw19neKTcj5lM6dtzKEXdUp2IHIKap4mVVmUwag+GaPupt
tUZ0gYMMRgCgZgexJLKLZwPncIcQox30hjGN1QiwffqbR6ZjhOWH+fzsTK5OJeE3smYj0cJVQn6W
nKnbR1joLMx6ok+jM6kMfwCHS4E9lw4TGEfKOt4r6eJYAiW6VEW+mPQAgL7o83eftl27rOGWFX3Y
ErQPiyNmDywPo6z28bXbo4J4Wdg1t4ED7K1epY6yw94iak33c9jRljvIFWgYEutkbophcL0S+ZP6
Hz6lOGfe/Q3tQ/LDjrQEb5gMKWRgSdhMRAKtDfNDnPU12YHGZEmI/GQT6INBchCYsYDOzW8E16yn
l0Bgz9KinRNtu/inh351qSBXP0kwm3fvKzpGfMyzHwZgCoq/RlOwHTnQEfdUjbfy/T7L3muAC//F
cfemq1FLx+A+SPvL9NwWI1a1yLh5aAwSnWom099/vxVXJQtnYA3XegoMbNMUKhwb5dYP7XVGNXYi
Q3MHRNYYXfwznWPOVUA+DDMAboWyuwydTQNX2erJI5x/Bzz6rGU5lKCIGoWAacmeTNnfZgjd7+dq
LFusoh7ubpCdjl/DBn8qaZc1Ajx66T3wnfXuQHblgslbeXHJsCLzMG8IU7qXDgk+WYsPd5lVYKgW
lvjch+PgSh4uBWArR5phv1xMnLdiEzfgJgxVTRz0Is7T4y4tClTpDFIitApwif1FEeOwv/PVXo6f
HhxRO5LEks/TYXlP36KFCl4NMIOEx/DPGj04YYnEizDp1LKvIJVk6rL8vOqv/SyvaPEDWXwWC2bS
U6E1LMrQ3flxNC1h45rPxt7V/7dbLt8Ni1RpA0tdyfiRw/cokEY1WfEk5XCE++Kbuo67vfIuyGC8
3DVuEPOQM2+t/FdwKy+qaKL8SMgTyiWhJN1l4KDXEZtyX+u5rywNkCsm7k9sh1magc0pXlbtdM/r
QQ03z/lw2G1qtH7ZRE0JwlqxKPBmFx5YsaNN1USlOYJ2h9zbVyek3J12psSHQevnL0T5Cvp3PmnV
gD6v/ObYbdeQ15CKnfmgueuiKX/qL2yIC6WgjlbXSKi1UOhASEuUUp9pbRr1UxyUwiUNol9flhZ9
GqP/aW3jzwgj0p/8aoghAa8+1qfbrhbhiVVGNgN71mA6Qyf7QbJV1tTDx6cgMSnsEwLdX/FGbBet
y4K0sYVcNnoF8exiCoJ/MhxpHJqad7UEbC8cKj25RGDcqHpnSIo2Es+RMrs5cqjTHMibIxSKoGOG
v43TD9GEptGYwdXtUpjHRY9Fw6i0JTnNMe2BTFSerP0Wk+pxYGmeQ92mN0duaOcU2WCorX4gRVJE
Y/jmc7wW8I2YFFQOvvesGU6QW9t5JAWkfNI6tHpxepfSAx1WNPET6l9WECgADlltNDdDQtI8eCav
v8x/KbaUUmbHzAovZvi6d+Sy0ZoZ7Yx5YNsKPURYHcIJ74JdQeZkpWHxS6q2xr9b/J2yiO1MjhF4
MUiKGZqDzytK+Hs77aHbtMRFMqjOQuk7EvHKNYMiJ9fwiKu5qFOUg1YZPSFoAE3/lwWVBLD85RJp
koeU1ppZFod/+xE8pYYoLLFIGyaK8fSDC8IuaU1gW0ABEckpLQj6dwtbIBo7fYGp/OAxiSExj8b7
SE8TU3tLncDLDdxOmjpuBt99O34gDefz9N3RCNpAmUqUKgXUuFs9QhHWx3DqJV8HgcoJEH77o2Vb
9Jtf3s7dWyw/wstHlbV87W3gSVDXyKRDEozd1TbKItbethSfejhH8o+E+x7J7oqxx+K7Wo/J7Kt/
xOS7dVwG9X5tNmi2ogDuzzdXn0tluDnuO4FeL67yH6mba884cDzR9zNKKEzX5xbyBM8ly7h1iq4U
ss/vJTqYqzdDi6xO8YePLjcTj0bmMsf/UwBAJSdEzykxoOhSiYRfeBLrN3srFqsR5wkWoCrpgKtx
0uohAfWEBDLrwl9ynr7K1tIyKARK0mnswBJlT8JErVfdA8zl3/Fb0DOJk26gKsT9CQJ65+2PUA1B
04tlJwjneBodEFo2OH3je0sWv9n/4ksYmqE9JHEY2w/v6jQVwgkRinKKw4TENCQxS59qfK95LZOe
vAP4WThTgLYRK/ebPmuLdNpbDAKFA4J2iHpSScZrWgC1R5IvANTowSQzZpWFsGeqCo46mN56Y0Sk
Zz3cAyqOChk7dATv/RS4Coq0tHx+de+qt9TMuIAGcOdHn/CrSbKL5n4X6lKCqAdbkraqkzJg07oi
t+Rtzj+l6sfFRslxIfE2YZBF7MeUXGs293iNaVZIy9yCItJ1b7lyExjreiEyikQcMSFqJy4RborQ
/QZI+aELrNSvrVY9ycV3TgaujSpTgPwtBfHhYwCrgvC3yd0G2dottS0MsN/TAUExpQGEUqE5Pet7
I+2CRGTdnVnlwkgT5qc9e5rNn4RlLvPbwhwrtbcbnS7bPvxzNeq54lULbrmQzirunsZwK2U78Zah
4pPo9EeoeBwqNMwVSJf/O/9O18p4iq+4kUmCxEihSMW2zKno1cVbuskkwjYWEO/dkxUxtNH4KtrK
5SGx5RCCOEFp7CUnbtVN1Gg8+beWSNflmOxkz7V2//IRrMO21RnQ/y2g2iU4Wyqk3hdQu7Z3p2Xv
0nqNN2ZQOly5o/gPRKabP7ONPOLa1VA4WOxSX/nut2REvElKytXj1nq2TfDfh3D5Tv9/rRXm0CEv
joeWgugVPCeIGd6LnIPVeH8HNOe1LBs1A4joZsQwXPM4XvXS+DshRsLn44oFcDbYAm0UM4YRzqzS
UJz/WzceY1lQFbrZZDroTVz/EXQHp0R6i6FkjK6Hyd9v5Ld6DBAKTf26IzepQ4inHydm7+9PdhSQ
uvNchr0UJwckG1XB4xgFC1jDYSoWGAq0Q3VspwTwtY+U0H7v+6lwkjTAcjxaasIYCgB3EjUWbMJJ
q8nXy7iRABCz2rvqg6Qs5JfJra2MYO5RsNdGihpOC+KA/YvzmQLBWGUNefwsBRX2DE5+0IQStNH8
YUSEDhywQ9EFld1iV9w50nS1hdTdp+2q3s74OQeiO6L7auyeHBCmytLWJsTuY5NoJH7qFB70aGg3
XXLN6V4d8k/LHQDdQzUm6+Pe4M7cDl0ISDPxh/oTIT7ka8Ap/kUOHOi7mBw5bGkq3oiTYC3V5OP8
9tmwED3CS1sX4+BoBXBDFhgoNAMmcwAS/4lOftYYQAemoqBfkXNsUyc4Zv1LgvwO3nPdOHP111/S
U9VODo1fnKlMBgVZkG35OQrDytwTEjdgb6OGVjH0qUah6hNPaxGn8HkpTodSUFDrCVmkXyWJhX+O
NKzA6IEoxqGT5zN47Da6uaEmnwsuGj24HENkGtg5nWGo5nxYMc6JPzvD2xP5jWiodnnkb+48k0E8
rL2D9yHe9E3FPpzTq73hi52NXXOcS1mcprfnwNrbpBA0FJ8LOucskhrWrwMYw8LPDFqaIY1RRA6R
uNeMqTgBmJY9/g1A6UnF+LpxpUd4TG77ghN7TBP2bOrvqz7SUDhw56o0YSjQW2SSL4fbeeTln/oe
6rYHn+AwdapWcSnaPcRodcx4iFZVl+qbdEV/c6bWGEsB2ZGZcPy6K0+DonIr4QPhgeVt8GLhHWjV
cxvp5m0ZQLZ+84JTVGcc+Af0gNYG6CnZvHxfDFP0Ktg2gt/xePjraUA0qDofxXQVUhVjC8toR+wK
w82yH+KIgxGVaO3HEXgxtpFS5TN77KEVdhBGkNq6vFT+4luYNz1AkL0Iuqszvt0rCbhFV9qRtvP+
qXiF106KC9i2V/UX6puaUOH5PHFbGEYzqnYf25KIPWsjfDf9zA8vaFuOAujlZKQFQ2ADXqCE0oAN
0aYrdgFc97AdHcQbqxtMclsH12PYhX4ged+871sJn129Q9R8wNnYYvegrjmxH4VVc54QZuXFBLtJ
1KQGmX4n0qr7KTFmUP3zM7i3cpqYdbkgJImnX1x9c7/eoBU41fHxwBGSy6fO02hnhdlulaxDcwED
4DLAKEAK34oiXq9JPMQ+U2L30lSzDQ/kGhwrQxoWo5I76Pe3pru1kexJEpVFH7zd2ls25dOSYC/D
+HkTo6qgNucVqoPJTUtTLW0vpRhAr1LcQYh/hsVbF5TYpSYtI8ykodYlgLSYak42/BiLYEKHUmFC
+O8QMZiOuZggGec36KhPRxdZK2IMMhJ1oailbwiggbEqKHNjyD1tOuBY5PF7ICIuDEDWIFVSBjh7
ShcN4yx5Cso3bXy6ILDgy65q8cHwltwd8fkvkBKnPrEKI3UOwUBf9ktccjyTLla0G6oE8Sq/R/Io
cgNYuEZoKe7Oa8I/y3KYp7TUeydpM0yL5j/E7aEYDiKh11/SmZLhBC0HrXZ3UfYmWNh613OsvVvt
zIzFD4MO9YJ9huhfbB69RNs2H3R5S/9GHtMxTtawyTDuULnroFEuQyZ2lE5zQxWiqawSg5ssAes7
cpJOtzBBqgHp36nDe8y46JfhHqvyTx/pfb5lvdIYgXz5yiL8SXPmfWNePVr/9iyw+KI3hxj4bT6j
BWxEoxKCo1kIwTnfNOBkxYKkL0yi3DcQ7hxRYFQJ34HgzX8D5cqCm+IgoiKqGtTiQ/YktE5WiurS
6o3j+7g9xBA/fgWSXYw11fThRAtcJI4i2aF85yWrCprRGgE9fM0yvf8KOpwgA+k9tww4vWXvlJFs
XgVklyPkLtrmQLlIQFJCaQZHsRqFrZk1Yk1T5hWL6pKvmK1p5IeIWQD1ll/c6U3DVuvoOQn3Xg4F
lnas1XuuZ895p8v2fvqCXg8NA//MrQbreSprOem7xQyjRyT92sMMH1xsx31yM6pN2jkaHKjZ8YPi
tLdEhxveRtY1VNzXnN1Ze9vHyU/lH5WQ9TbgcOf87oTO3DHUN2THIjGL7+TqpmiGITaUOKkH9PUx
G+bg5Ucu4kCxX2E40509lWolk5bo0NcnV8G82maWnwts83fV4VveZZbIV3Q9E7QLSBImOontq/EV
ag67u5SG9+lUgWHkBeZOPNcm4lvzvyOys9t+AqSiGjgGziM0TQUuSUXU6K/TGgqQLjKpMD4s0+CC
WzHjVIKh4rjA/tOLp0CMULAHajtkVkBQkoOuQrYk7UYY74GnxcJjfm88B/S7sYNg5S5E2vs8OUxF
pfAtpiszNMItPVjKp8jPqmQ0XwUBXMrZ2HnngJqjVmx1gF375gU8oGmwlbRoOaQ7N0o4cqNdprrK
lcKR4k+h141aUrUQkbPakFwLfIqHJ0mM0EfCREx1+NIXhUbRuF1EgNOfoFWqLC4M9dM4aXNXJFHn
EoD71rV55T6+r6aDW6k8dbyKIdNsaLnTnEVcMM/eidmxaxzm1lbAP1nN8vi2sBDLuxTc/wDla27v
+ylTZ7rFu8qwSuhLcTPTbvL9kzy/XiWaaxNnKvlP56gn4wCP6opscStyH3pTNIJq48M2SAeR10/B
/8e+uGUgcYvhB6ATm0+M/K9/pBj9+hUxkif7TIc8G5+EmhTs+mJ2q6fCzxhqzLYNiBwkcycqvbWB
5AzjjmKsQTGAeDAAww3m5k7AR6ULK7nvMOpxIpB1uwXSzyyttALqdYiTsWLajIyIxJ+emSLcEvyw
sMDbU6DXrWpiwdfXTu1DWGGHbTcyvML90A+j1dhlz3Mw0LBMrzM25z4cnItlb6c6LsxQk8wy/4ig
5BuEGYz2DRiAUJf8cV8L5D4Arsp2xUme5pKsUeeZ9BGjOvI4Pes7YwylNRAqLtjew0tIuj1AeALY
0Kxeqj2W8HorcB+xZosMbMSPzAjmcZvS+LMa6W6OiZDBBPaXzJemHl8ypES3KA7HAalv8MhakHoM
/1TVjaWRlBBX+XoWydT2ZyGVJiTtNEf2o4GkxzXMGp9ak271slgBQQ19EmnyCvdgF51a12IdiZnt
epk53XKX856eF+GGw+LFuC2K9M7G8YsRwqL7dzCxENK8loZgqw1J14+hcY0F+GE7Ez/8POCY3uRo
2OegI7+Qfj/1Sqvq/F2CmBQSHo9Bf54J+e4VQEdXJ9wxkxb6aIu14WZRJkjFKK70v7OboxxT5SoL
6PlsUDeVx8lQFK/I+ImkVotZbQ9hVkaxqYms1+aspDAE0rsMAq83jNRS8LygAcv8hoHw7hkv4TdQ
N/RM+pjAf6J3lWl2wE4WtixuSmFpLECpox+d03x1OxY5XxFWrpMYix5Sgpf7jh2FQy9ayI2HTwlG
t4wMyrz16ysZ5aZF9jt9o+IVNrYfNE5wOo9ELUjICk050h9oYdSo5+TMvzp1LuajCHFIwoVs0rdN
6x5b68rnuAFY/Pifzlt+h8utEkLe+q9bnARAzE7L3LZcynQm2mBvT9JLK2XlqYcTd3ji84HTLW/t
BbCQYMgzuI+4TKG8HtHAtssi0wxuvMPgMPx2XQkjiQEkD+2kJLOcyVmyba90g2n1VYU8+TmKzf9y
+vI9SlALl5faKFOMnU5aNcQGO2BxeIOtk8a+URmR0yTI042Tdx8ecGagOkTcRSwGQmEdqAq6+2o1
KyPLm2JJWxfhV/9e/fl3jxFZyzUzwRMlN9IHim0SlgJjXFPh2DAZGTpVuq8xumm5dkJKEkK09Jak
t+bQEAbGnwXkgdnZPkN0v6PF6IUc4VyAvWvq5DWIlut2BjQV8mixPmRFGIAZfHL5PdHCAKLIVNz3
1q/N+jSGip6i80e3B7881SURnbzq1fYUbTcTPCvN68fSNckjHd3LCaDv34iZdNh6RhyVGWVsP/22
JluPXENndVZsB8uKajbYk9yryFX2NcUUcrVZM2WBytvL/4qN5mk5s3lyQgsSeiFyXQC6gVwhMLq4
GVhjpSGboGNT5tgX+3xtxZk1iYTYXDrBnr65acmEsh1t6v7Gr/QWTV5zUTHzvUYJhIiNTyoCYK1t
bkHQlqc8xLZHVx7Vs5L7glR4oN/ACneWeRm+pJyAGPWW99z8OXSkElqGW9Re2ttprfYCqFzsan4k
wcf9vpdp4mVzRTbU2OEtl+kYYGcCpB3RgPEwMb0kCbetacs9zvOcvchHJZwiWdvbSBCzQnBZ2yrw
lbIlVJyXzWSzNGK5mo7RapD47+JaisvjDK219lQUSuripstHMmoXaCxwTbr0J4quErK5NWIWQw8k
ZjAyQWVDNRSQHXUrGO66YEqW5L56zkP6cGUqckKmfo3fPBM6rNHqdpnoNz4UV+BIHbtZ4WtfQnEL
1nATJcPNYr+8iQOebQEVST6pqTHbcq82teHAfxOKb2KiBZlzvwuAoMk8Yr4DnSguA1vCHCNFDjRz
s04mKgiUDDy8708vGcT4qUM8vT3VIPPrGZUU2DBAUv+2NEhwQAa2v6/sODgPXOq6acaMxpqtcE8T
Gypa+vXcnxYuhL/Jj7Novak8e5LcYzsNIuWEV2G70QVUKqLOuF73a/p98BEoPOJgdqQ23NLKNxrP
W1r83Qe25K0uyyVuLwxjL2Lw7AWJXaDXaeAKNdNs4D172lTTBUOTNOfi3Vbz5B5d6Sv33L3IC5t8
JUUm/ZJ+bet24WLFeSTjVk/8gBcHYXF3SO7JUYWDhe32tGLqcWiHnNFJAsn5KBWZiXYBFa2XQzL5
xdi8952zp+C5Kzg9F8A+yXDpuGJX2GebJasgcXQlmFkzBtBxkz4fQzhM+mJFUU4gb/c6MnAQ0h06
dkq8PDxVk2byrW0QtcAinX71CRejBGFLkoYYnQ7Ony4gGyRB6qhcAtTNxdFs016nuG8pJsgoq76d
0VCqH6yGCK1vMYnFXJuUoWIPfYSQE7uRv+qgdzNbOORbSTp13Ckbeh4ohl4e4mfGgk6gRKnvHW0/
kIWOy/2nC9XRfP8+21xaLNBs2hnENpNs9xJ4hv8+TOjyj/H0cYRbVUKkiBBN7LGT8ffsyLQFjqxd
KU5j2pHClXdtDUW8msro068wRrOk1aVIvWE3S5E020lfJfV/rxHnlY4Oiq+PInQeM/iUy4xG+dhP
BGNqQrVnnFzZBPXLtmUPKkdg7hGHS76b61ZeWjBVQAc7TxJhM3G9Mha6TLPjMAguXxBxymWK6Y3L
qLwQmwtZWI6JQb35Bodui0owLlPM7MPSYPZKwYVKD4zlCRJtv2sp399O/72fWb+ZFhc7QXbhC3h/
MbtLX7g97nTvBi5uvqPKrAUbl7UtmFUmNcMXXH8P9tIlVaERRdstXLS7wu6LYLMOOJMxCXtvTUdV
OO8EtBujUX61UaGNanMYMvFJKih06G4NFHjtMMXNP9jcAMcKOCCcJ9dNG7uYeHnurb9ZEfxl0XJx
oOoXoJB40o+KDsIjb9KOLlgpPEBajppMbEBfeOlt4VyZ6Z8lvDCYmq+oetQGzto3FRNlLZM1SFLv
/XQnccaqLzT9NFr0IFDLf1rqV6izhCSLDjNPvz6GYgPbTbkDB3CmS4qVxAts9S+j3KdLEvbEoX4G
ivhcFItfrG1D5HKfD9r8FBAf5RW4naVEomStVEn2VQDRXPO9GiNmLyqOsYizLrG/bd7rhea206Zv
QN1CCLMs/cd2SIKQkEtDMOIizT2RjdqcAdrO3H2S6LXZSZ04Xs1RuaBvjLdMtaGFyp9Xft6FLBSc
pggK9CJB4aMOEjyitzGZ6Z47/LoajgVDK7aXKo+huFUgySX23TnQspHIOeX0MVFTKDT9ZI2oGm55
mGxIkMNGQWGm5OYCrvQS+6VI0D6pm22oCCzolsfHjt3B+qBRyES+F0sqHXm+MWyhOOcIRCENhH+l
vRsH7ZQ+2LeTNKVhCW5OYpVqiUg6MAiQpKP7tyOGw2GadcxK2fX8bJL8qqLnrZGs+T0T7RRwSFC/
2mrT62EZg3Jytc9ib/Ma40PowTVdSqAZSuM5fHGkiGBsYzOxyQPVLTryYg/u4EZpsyIG5PPKlHjk
K64HzjaPUxl8DtxbUAlgMGkzrBGdDRVRU8ZXkHKdhUj2W8XzElkLfhkOkcBglxo9kI5/A7OPOHpx
3Tnq1NxKL6eovZ5ha31Rke7LBUXIWWG6rPpubLuVLRzMv6EXxEmmjoog5ESd4ym8//yWRfi5mo5r
6ORko87AIIQV/YNPWpXQfRSzmQPtCKy9gvx/Xpz/wdgyYNalWATMyZ7IS2+046IBMc+DdO6zHhJk
miW4rOooRAMMAoTmv5c8lE7QK6T4TNVRpkWTO2hXtKocApe+JkAciAI7eMfTh5bH+tfuHdFOTbe7
pyx3YU0whvcSdFKxmwv+rvkpzLMKig3Eez12NVwI7Hqv6aUM+n2J7Pr1hG/m3w5zNVgQdyDAjrzg
Pr223pSV76IE/9i1QGFd5ZEipfvs4tZEbfn1UB1YHoa5RDLU029UdWsJo1P7eOBeem6KJAnXMwek
QwHfC8GokjjVZfOiuzCZhOfoByj2l7xk/OpPuPVi7IpIYnBRF6+jee6G9Egr2N0CsvpXSnsd67WI
QDUz2dLkwZ92rQs+BI02epATHyrWTSjslCkz8L6P1ZhPn2DM5qNEBW7SmP8Bck1SZEVVkpgkMAwg
0pV2rXaNV3UAfopgraPpdypx3RRcOF5cAAp2gMJ1DL08TAr6AyfDkhQE6eAEKNnoDiK5ipPYwcd8
9Pjy7UTF/rSqS3/PrAUWGk6nnBxXkt1wvKo1NwD0Q0OjXyw7ccZ7LFyNoHgWzRNNuIbiFiOAlwvP
CdKVhQVEdCLUIYE6Q9zIBye8ryqGzRxRJXE/sS/+pK1qiDnA8trMk74AfkoXCODBuw2Lyjb2wIn1
kr/sNXivhgojE7o3LuSovDuOC5UA94IZjZVRN+z3SkBQn32lkaKhr+8WkhU3e3EOF1FJr2EJwyvh
1b58LGEgi1o1zvhwmnx092LocUMI27e52yl1WTRrYOpPPaKNhLJZDJuN4mwSWrzo2R+EZ2rfa9Kj
t6OElijGke1KOIoDgZzute0uAIDfaCMtu0HApnTSvTFzX3g+J6dex/awFVMt/od6Lajrcu4nuIss
/a2OpcBclNheVdkv7Os87VJGjzyT8TQcpmYqTjPjtnMACGGZCpqumpuBx/QoNSKmAckjJR4LMKRW
P4PnpHmbggxeb7M3B8sJfy6V0+bJjmvlWqW+PjEUIuah5Rrc9kbCbksypst9wlXOu24zLFrZOq1z
AptlrLuYCJh22dWxlW2UuuHilcHDW7ToO2fvvGSUZbVPkytkwYOVY9YV/oormwkj5TWTwEbBOBhD
EqNjvw0uwLqAqaSsHJQOyrAOArqYLvcjBnFvfBq2qtyatr4jo6Wg8jiSaSoqluS9K+IDNtRFbqAg
5bZqwoZgs8+HVzDSzImjW16bjtZyNDKdMKnMP5D3MjEx4R2bBrRauz5vy2eEzmahLNJFdOGieHyZ
PgutsZd4tMbRdsZ9+IQXHrZ6xRviWG1buydTtC5pm6XWHwwXBQc3ZhLx5P6uLclnW4AWVNgXjfJM
/vGDQlCqeFxBwNmx3Eux96//1yc/4QjnNj2NtJU0djx5AP3O21OlPMtNhWgx3dKkNxAuytd9tXI+
I3KRkcZtbhdZFlYS1OYnjNmNhINjnddb/wfiAkP8D9Z2vYBsRiZOdbEl/y/rN1XHUmwUKcPRSJA6
JflKYULGgv1VQo6Q/qOShPrIZsaufyhFiezA9wfnaECP7D3Xw8BNiVIy5XXyXgQoRRaCW/SyE+gH
D180epmGvXLgtubqYSGaZBX23hzm3MXh2fxLwhf6rlhFE0hX+7PEt/EFc1Qa415LJ7IGSpAaxLX+
Z1gFvGfKVg6Y73AOdAYXVAmEOEnXgJXJCz2hpDjXhNhJTszQrC+6vtPdvtWnZ/cBXE3XLTMCrZsh
NJFljmF7ldfRM81w4GNJ8mPNsUcqUa4mjTlQ1Ymnybq1oYLde55puR20sLl77QRN5CZqb83zZPp5
9KqAfb5iRkApjthndAK7wSfhb8w67IHqx6GP59stFGvlhzu7MPRxFppjTBOaPEUjmaEelSjQPxwG
ZR/9QXKgHFMMdZBop+Yo2pie7XCoCaatoIwqZDDQCnIc5OnKnOaxBn2ZUFKy/ASrn3U6xn5HYRhc
ClUoQqELHSGqs4QX1X/DG9E3QVLPbjlZk3Gtyc0uilI7jxtl0g0r7n3Gk2djc8uKx1mtuoSvNqqb
xhs+eRUElsK05LgXrE0fd2V233Dl2sfjwjRXyKQJRk39F+xHlxX2DK5LnbVh0GwrgNK9Ymt6W3z4
QRDg4dNHQgR58e0VF7Jvcri8F1umMR+NmD5pnMe4Dj7IHrFfsifXzPSfm30waFAOVp9/zdpaN4Rs
N67WrzZiIpHJsMlyrw7FnQzQP3VdBUZlvDpV7ZLUmzC+vF4wg95XoYkBJESQMeH6BrEwiA7TPOcA
OZNBgWbSbHHWFVMyX2V2XIvIK6+eE2i5xSJ0kXEeTuEnOR8Gf9nblHxtszcxOUy4xWKYLBESTH06
huiD8jblqpFt58NvINiCrVemH1iXlfBu4SK17r+BkSTk0Iy2yF5PKjlfZ6JF7u0/fI4s1ssmE172
sxtwqsuHnGjbJstrT3Ku82sjVJ+CPrdvGyeb55yuRKWmMX0GPxThwCqlVP/0vPsrGCg/vF15xwJY
LyMtVUoeYr9XnIVJXQi9HNHaiZxR0z21idrhE3rZ24dj7os3FEKRIRy/9ieQ2JoYIZ4WmN+jikcp
uewPcmTmv8FB2JtyXpWWZRyqtE9uU8qeASUpI9p9/y7SAqDFpjfNmivHQqFwVbUy7Q8FPllGEhDW
2NE5ZcStEZQ5gVpzhTJ5/I1ry9blFYHmDj2wsNG4eaezHYLeUY7tauF0khB3w34GEgzX32Yv7Vur
Xk9f6lfNePhVsNroa+KZ5SMmJOB3ko0C5dRRHUw1k/y01IyPMQ7uBLbMydffwlU/lpCOIvwuu2Vg
rXKaqhTxa2KFSxfIrraBiG5nQkun2dOt/NwQp6DFQ4jzW6gAAobD79218MLNAK+45RPL/PWrpw1Z
sXOW2LyPAXq30zRp1RV0vcFQpqcoaFcIO8P9AVRPVQRnFKK8RBB/9PhaAushH3YzGOwdd2vmyKcM
Wkk5Z0FcvjbwTVoOt31YSUkmLaVO0ZVRttZi5veaLCbmQw7/urZPrBIr/N9WT21dUgrlIk5cV4Iv
YtgfKZptAz7pipxDdeCL7y2o5QZMle7c8zFmzRUKH37RJtujrTj31A07tyUbCid7P0LB5S45QsG6
wkvVz7xTwDIdoVCKkDSmO6VSraw1QshRoAYVvFiDj3a1nuNQaVMYWa8bA2ZpZjui5AGvTMjnP6hS
wCMIk/BlHgFqTWFVp+ZhhKnH32CHAmJNYPaDoC+FVMsdQRPhxuvhV8ikc1LyvZp7UZjtNy2abhtP
CBWg6+53eqrIJMTbvUkP0T5v6du9OoUFgg7vKGMsH64yhqByWVWjcSwRnPXlzk1Fj1g//yVFfY/5
v8kHqtHBs/uYpyebuMHToMxAQ/RsPITyIsIZMC7eIK9bWtPEbwjGiT21iHSCHmKUte9nxnTvbBJ8
XOaJJdygmDm7Mwy31Sqbv3H/qI1S5VYEPoulPe0zKayyRfL4QcYnvXBXy/swqDkL1KL00pQLMOPY
ui1q1eFa5+ndaZocbRTIDvtAniyGPQuQsT4AXpsGS0pCFoOKT984c37sBkvINhTvZNowALkM6zyr
sNzuJy7Yq3W3fiHOas3AS6gxrDTnRnFG9ip3IThcYZeT3ZhwLALMlDPyLkcSHjuJvhuG3FRFyYSF
OS7T5PKiFQOO8LWXeXlxNzRlIcVi6042ulfzl4vgkUwVLXVLzWPb5DGv/HNcqbh4G0jIevvQijv4
ExgQ2IucuZP/mEKGnVUDJLOKGbsQ8jScytsQqfcoslUBxs8QFm9sIniWjQsJ9HREh84WK4GR+bh3
lv+UU41h1KQ0Q0BzuQdi0DB9NLDZbmDKRu4FDKeRkfdQ9hGPf3OS7YxsZjd8mgMHEWrbwJxhs3Ld
wZz5PipI3Nld5umm8H6t3YX8LkBj5T2rHdhI+3X/I5C4MNM/UEjeVP+ti7Tl8SEqWMmx3UQui4rb
7L495xWq+YjPYMU88XhMzOFjEs0T4glKb8GVxYaN2PmOM33UkrDnj1XlnWI6eCUY+RlOsUxohh93
U8YmXN9v/hjOBVqCw6azpdQDQGQTq9j+NJM21hlE3fwttMaxfyPf27lTJuPxluRmFRVeThosKhmX
aOv7bl6YXe8euRmSh/wUzeCkIg+8gt6acy/l+XC4sMQJ2UGfIVj24reBmd/13UTwDH0ILxZ/ZYYS
cEtBl2agBK8rKOwWHvbGtDQXhtX8jWkhOhwJOl4xoGEzYrerGrhlGXbKhSXYrCLgaAycsamPKxhR
rY2VRjmUDI1qWMhY/wj3DOycnyWM6SzJo5x8CzCBcpKGkaZC3wm7NA4anGgR+mPt+/OfE8z6DUYq
ZMK6toFc7SMRsjGGqOIuujC9byt0+Ck7PuSK+WnsTPRUs8lugALiB/NhWy7UFcV0Gjlg3gUZQim3
v35rVH2lqkj78Op/p36F/ENnk85CJv4mr9ijHjncnnl4ty2k/TbgraZfadgMNwvjQ79sszmr/TPK
rBEUdBWeT+H5Kn+r55E6jdR1GPcuSkN+78x8hZKaebPWi3gGrl2n6U+FwPqYttum46Y8t4ps6sfZ
+PqHejmj/hpeTfqZK2erFzt2xrTso3q6VG4O25tp1QPQNQgLz1K0Mk2NHXwWfxy9Dvr9pwGXadQO
CZp3tBHGVGPRJdk48L+1cPKQS36VrTSjuo+Zp3/+Ymt68Ux+4ZZ3e1KbHhVYOVBtnLAJj4g0+LBr
RYxYI1kvMRJn68OVW3IcY81aiC+a+oZx41lP1UPixLXREgKqfsxQmNW5go8/lGaXM/9maUphqszu
Zja0/Pws3BEVun7aJy67xaU3q7xxtKkKfcZcuITCFBS4yKpV05RhlYqQm84GWe9wNNFVWhZ3nnwV
8zPrQ3iQYvKRvnbUHGg96ayUu+KU/YpDP1HdOVbzyQYJbLBsDYobyO96+VARpagvx8IxzrQbnXPd
d6xBDAiZKyxXG/2sU9yVAfldUmzB+JbnLTOHO8o+0xodR0AgEVM9xqRZPzVE/g/JHrRg3TOSBjez
8TiW5+LZVd+M7RVwhJ8lvHzLtdgEeex6A/CKwq3L2ols5cgwNIEOi6KBTX6MdA007Nl8JnAMRPkK
4v7jLNMm15PvT/eATyK3rTYCEsQXCfxu1bWFOhY8L4YLPRFGWYvva+28m5eN4K4NrOUmgNnYr7o+
XoZNgFOeP7Eaqq0yRseCFz/I/3jLLgU6iRT9ViDOi1vwYiUrSYjx0hUv8m4yNpZ/t5TAo65zyIHX
fBdo6SdAdxisAxvs6QbYcNKZPYfzPVxOsYM1VlIJdBN+IJ1glaOrqBL55JJKQCiIclKzEFIbcmQk
3p6M7DbZYVOrTM8yw1XYazrMC5c3qvUxT22WbblNUzPbAseQyU7O0xcPUcxkwmHnVLsrqXVsxdP8
4ENr+OmUYIrJIrTrtiMxPgEbnJxw8GIXpMQxeVqolGYoNmT76KCxE5qTiWfrAVkvoJ5yW4J84JHD
2DKBOK9uW/sedy0SLRg5x2KJ7JVG1AIxj9RnqQXkq4Ytob6H9HWum9IQkrNkGugB2W/aQK0Dut4q
Nlzm6Kz+oq7oiL8U9TOuDTD6WK61K2z4Rj+0xqZ8bWIC5TAfBnIpHBrxVe2/I/B40wQsRh3taxt3
Cs14np9pZud/DqyBb/b5V+gBMMOvAU4H/tuSR5+tYVSjsMGcCBRRHpaLYiu0kHfVEV7iy3WERTDt
9H/m+zL6+OIpkCgv3hyhlouT+EQyoBVqY78nseX+sT8bfoiuRbrXcgnmUp8uBfzA3yeweNgvs09O
xbEB/pKF8KbbrgucPtdGXnUB5pQ2BEvYJebJZ+UdNrU2drQAftc5J2j/Bsk0PB2knXcWYE8h9l/2
PCfSLP5fXS3U1/BXBg206i0p6Mtb5O4A6bKccHp5y1UvoCG9BqskDskxPAmieEQlVl++sKsZ6o2E
UDgy2L5ubiebfuuQokGb3OYLhEq7am95bctnTdX0wlHKLC2ijeYVkO8XAIgp3O7s497EzwJl5s0q
MNgiXIC4ZCA8mdN2J6qQ2kFsx5yhQCX3npqfiP1h8K32NIGKWJ6SeuaLB1Q4fYRpyo8VEswI0GSJ
4oWz4FItEFrxLh2hNe4on/P0yApgkPOMldGckji6LDvHpEbM9Eekn0Whuua2WLQD0zWz/byGCufc
Nbc5bwO2iRFiphfTVR+HSbt7qH5rAnZKKTYGGRnHAK6ekGwnZ5vbsXGPcj9bRE9ASRdijfLkJpCR
5vIpx+Wytv8kmGW/IIrFz1dzEj+ML/i56rhjsxauvztcihxMKe7lkC5VtBIzdwpWOiTluNB30QLH
sgcWwC6DLqS8TC8lazzZ4T8nViCOAxCEYdkWHWzGhRyU/uvGVYqyZ1m5YLUGJfREyu+nKaOu00Dm
GrWmI+Z4BBupyU6lsmApIZNzpmSi9RuCvRCl6eZb7cRJaWomB36rnkiCqk9QavqhgsTKAEwHh0nj
Tta2qb1qOGbVtitKnewHDf3B3Er3Hfe9lTXFCok27BTVvI8Q8o10r3/vmGqJ0ILIXMkR21DtP3rB
xd7TxkwNqDh2bGBQzYaQEIbxDe5t+oM/Aijy02Y80AcUtUvAABCmPQAcP8WVc5bynDjFBy9N73PA
i3zerHPNU/m5pbBNM+dU6aP9U23DiEs0mBglqPJQ554Gh0kWWWePFUk8J9k2MoCs8uEZq1oOeVTl
3JzkBsRqfsaFipxbllWb4LYT52nFKKDWjV4zcVYmm+Nvq9hB4pQLUmnXS0ewvt24xOZ/ltR/xSN+
1ZiFIY/RmxrWMG+E4zoEDdS9B1eMDEpuhPn2UZUqvv4W2W5zV3U2pjxMfm01YXcFy5IVod4zVcfy
vrXMeivllDb5pIjKXJN4Xs2V47wzcEP/ncwGokgBU0YxH+B49TUSQ+hCU5f48eFmGnd8RvTmXNOS
gsAhZwFlf1MeU0YY1CuHG5i8GnzWF1mEfezAKkI6CSjddjKf0eWGvNQrVDeUhrDsSjmOeOWcFJ05
LpY4F2nVaMTRn3IsTwEeYRPGn83vlIQ4ry1Jk9kw4OiqGeDMAO5T12mh0L66LdaV1p3bRs8d6oXG
Y3lxICv4eOFUeLZf7oe5hBaKpSbGkOfF4RNaPzqzgDlatThImiv/iprtFVym2EFzG2+dP/ksrJhp
kSjXUNX7mV38KyKOgJyfBa1zloHVLu0sYJhaCmlN4xx5Upt/UBcvzT0mjtemDkYupGuC2QpJeqJw
5OD4bYxt8uvrAeyrZajUX+RIj3xURkvVnL5pQnxGUisTzgNKIka7S99+dO3KreQ1JUHdx3glVFOv
Km7cuIIs849l8lIOCNPa711y3ArEwMu8T56iSwzIyYSA+dFu6rJHVpS+5WsPHBkfOZt0Obqpahk6
jTXZWzWgGS7ecgETKMQNY9f52l9GzM8GH+xq+vLQWh2CKNdQ+Ayv2SebyaojMgT1oxSARklTjXZG
z5VrxC9ELa82ZZW8/9/buyW8JJHJ/BRvVJAxhab3zR9/2Yd0iS7+6puJAXMWRgY77AhXAfIOjmWq
sP83a0gDqbnhwrTAS21nDrUODvCgLnCPdlNlCpJBXeD3cgV+/V2jMiv8+nHdh94liaEflj6KxUnw
L6m+dG9Et8H/I1Q9R1IS1VI/dt8phKhOR9J9a5QOhmGzPZbNDnfWCciqFcqVq3uopGciZ2GCqhqY
vNmkB8rABVEKVO3uVMVFSuZBDOr7T/3NqqhAL+qcVCWt734zqwlSBzfZdbBtRLGRr0exom697Fd+
FjCV7AmvM32UFOFC9njjMFawpbmVaPgEQMZsvi2E+udgcikqfAq/VuA+A1AeXsDKR79Yiwn5u8Go
j8rdyVCg3Vs5M968+9f50JcfZQ4nBOCQ0CbTT1v4+R3Mqkj8A2aSU4hBUAunOLUe2tRPPruwHEQk
SFFCJL+OGGhv/GDLuMkR+w/zyJ0JF3JemutoOSmfaJrs8UwAQ08FiXYjUBGAAVatTXbOOXz/JNy5
fhrvBTvnSU8Pfk9nwujWeMh/EYO1AAkfUQG0JrBt6RpuIPUeaEcGrx0TQScxIfVvxVspJT6XBOK3
UP23IOTSubkqs0p6eJemX7W3m6tinv9vBaMfcVnbPlS3Nxw6rXmgWk4ZS77fsEZYKwAMaf4VP9CJ
/kKu10XoOea2wDR4E3Cy3YKxVovWfy1rSlJVuMhMPxVEHXsVXnVDxjpR4QnI7GhpM9P+07yfo0AD
pTVk+FIV9aBIigkPIdwd9GqOEGdciJlhzhkmJt/YVHXOTceYg4sX2JyWJH4FDuiM2nq2V6TxCAou
UW0Bwqd5HNnibpxm1sR4GyFmJHLlsX4sJwnnTZ7xYqcwDXuc4fHcRC5asXrv34MMbplEsiQzcJ/p
yYuyJx2sl5v4IBoRFCV8FKCviHPRP+e2W2wE4vrUZHD8wU1XqBbycrwW5jj5KjYRNHLLYE94VWz5
nmZlU0cLYDVUuVxdRs3hy2eHWPB+mnTMppKcmJ/5c/zQsRhlc7qXm5Yh1t3gigfZRju7VtNDmSdy
YWEVol0UMKKkV88Fj1BE6jYHawVW2OEwDZL1/yAm0jfWV4AB3xc9GpP8V3DPKEOeFjf0/hntlnKI
8cXhx2nxRoUBw8WB4BoXGTAU/8BYttRp2B9DsE2WFXvOUV71BsnnMU5g7IcU3bAz9G1tbhWwGOxf
qa3U0Vhxyh9rFqvrXQpHcsBPcOQuZ3J5QXeVApWz+1Q7ltaegKr3ule1XkhskuvF20QAqLMUrbZA
lUy2jsmsmRElz2oGgXJxIdv69TB9rolphgzhpUm7ZHgPZ7wCi+B+hLHHwwp0ggioLGVsljE3vhLy
CHIQsD4S3NcUWUrfGqcmBxOeNrUfQvmCBrEFyGX5/JikIEhp826oBWBaED+ixJCcjSAO03UCP5Jc
836sAEBM3/haMUxlreppjNYju+aGJEvN6VdEnc72CuEJg/1i2Z+dxzqrAO9NBoDbEp2XBAehZdqX
tCt7eSE539I3+xnUgMLeFOwveMo178Apf/wr7b+olD7xmnero/1KrwDmCF/5QaExoQAjamp/yA5B
y0xKdLNUvd5q6f4sZsQN028gyKly2SG8rExJDHboi8dV378NEGbK7VXA0D8aP7QDcXJdCyCZgegS
vzrqBlazKHGHmdXsuxEL5ra4tfdTIfjWlEZvmSpMIDtW90u9nIhWBDT9XuEkVA/XvI5ThkY4+2br
8v/J+7dcCas6ihFd5W4TShb+96F4JqagNKplJXuUzlE4HyVCfw7DQbGB9bXF+3CRjTJbyUXRfUPa
EVJX18oz/qMTFA7PWmFZX+D1zqFeqPhcNinnwwzPOkZgcpvwRRGcPqh3a9bZ3dHRlOtt/QD++Zv6
NT2uKexcoQnYTbWoWGpM754gO4YwEh3n/W42GALe/Ns44R6qqX/+odmClWJl4YMs7DfvrXuM9pIn
CDHa4O28EKapMBMN1/Lnt0jD+xQbJMBbbKT3E3kxVSO4i4pVVSjFRa3n+109QIo3EnkIFjgznfPV
q/EeaWrOqmfXq+TOvc/QZ5wPF9Pq+2wRwNdAV/ThZivqttUHmEB7jfLK2oE7Jz8iZe5l4+wO45n0
Fozsim6JwByaQ/NZiMPsn4Q6MlkgVRwL2D67xRHutiTuyX90bhnBtVTFQjXPwjJb5M1AZEfCbNu/
7desaWLlRAdlsHlRcZHPfN+LGMpsT5hj43oCUgk+9hAdst35WUnsjUZ+IDxnbcqKm8bD/zgBPBBI
QJd4CEvlUhs4yvM7iko0xk9U34fR0fb5UpT5KpfzqBBmLe92TBbBEwTJtmAGVrTflct02S3B0uTI
tOjLZR5y5orrjafMxxTyXZrPInKjZ+6JoBleVdE6rKUZEi5rhnJZNbpzGKCuINoW5/lUF2/P+lnZ
5WtFbZjcn9a4SyTOT2BgDF6MPwr5j0VhiLLrMYZNhUeMe0mYNFy4vrx/lgGObL2h80uC/CYM5ABf
ZDa6Zl8bY9bxjrBeQquYVh2d9Op1i3fZYm+pCo/n4g+T3Rm4auNK7FNmZjSPZTvtshR05dw+gqKg
eB4ajV99QfeYeuYUAGnc4yfY13t2B0oflLD3VSmStwpdr208Tv63iHwlBBgSTiLx2nP3sTc8Dpbk
AvOe5KIMND9yKEzK7Caf3mm5vntRb3cxV2x6kYekncvwIk0/ZLSb7Px9hmp6zYghsZTdBdMdrhsx
5Of1HLJVsxBDSTRWDOiVF0V4d347aB/6GeyFiOVKnkK1pkrc6GdS+m5bR2yQfyQDOyNLtMzvrf7A
KIQNnQf9667gxmrME8XE4L7GluHTOShEmwsBQfAcag/KId89hyi6Jw6J16NzkKyxykAOL2jI9OpD
W1gErxwdgmUfBgw2gFUXvucAKqm2sBdIbnq5HYVrzcXHtcO3CgPHOxBiOEnNoqIIWQogakZxmeSW
h+SDM28tMin7KW+IfWJRrcsKTCouU+tmYcaA5ZucqMxxhgFzjUFFp5QM0SxEYC8UGGUTOy17QUIX
/ls2llRDWGLCezhkoj6JLKGz6mOhN0JMm/KT31pEmNN9JGHLy2uyM7Z3veXImMaTDzci10iSSdFP
eYBbe1WBCXCNwB6qiJMLHi5bnn7zpoUB77nWMhjzUhyhytGCHVHJvN6itHTA/7GQJrndm/qJAbXc
ziVxnTt7eE57YqOr+gpiJ9JgGvX2RVH6PU61u9z1/luwelts38squmDMeKzDe+8xJkbRXT8Z8bdU
4HDbQWxPNBQhhHmoFnIlPrSwbiDLZlyhGA+51YcbW2JZfNU8ey2iaWHdn4kwmq2x9OQBU8j8WujL
CLXFAJEibOpE3zOsT2py+vfcBJgbTwVlPcgTkw++fPmCZb1nJa38pX2Zsl1+Q+Cjz5vC8QbAWgum
80r6yMstIOyWiRIzvoxfQRG6OZtY9u7FuKeQ+glei2dBUx3/mu5HQoy4hH7OLsbyoMYksElPfzga
VA3dPljiyV1UFve6jZf8bB2BbMb5jfO2kVrIcrQ+l1dZebs2+MlPoshQxl7CTetYa4+B5yg6j2V4
jeawbrXlhpyuWWOeWAFFUxS4Gw7JN7RCzcXgwhexOpA88kjv/gvAzoPfTBYuZEKEb2Ia7b127Ktx
e5VaH85Ftu8BZZU45+lSSEiCqeWEHtl+C97372pqjz/L4/0fD02jr5XxTwGgzbM2xLC3nlxPGUHI
O9gokVznr9LvBVZPhCAJGUr5LmoadWY4j7iYPZip8nGDV0rKYVQn0xuWKEL0tN5jPPwhoaqAB89B
HKmc9w+7Hob5eQkioKmG8S96kRfuBDWcUR6vu7RkhxxzNzy0rQdB50P7bgGzYsSYUglPIFOU0TdP
/RbusI1ld6VKfmlZYoRWlifLRk45BT9pUzyuuRG1uH4R7timwKC596TnOjdrfGqwCHLGR6WVqRKT
dFu+SkqvyFNmJOwKWdWRmLxeV5JqaHjit9C5Wk0cFCX65tpSRNClcdanMTO/lksKUuLxDp8mDsfq
5WQz71JiJ5mLAofpx3OTMBdiIlZ4ed1Kd2FE+Skj38lPFvt8Ct+zolch4mSAqRrXRM6RdRJ6LTj0
zEeU7DyjlRuoR3qu0YDo2zhhIoojisWIAdZyA/qW/z5Cuo4Lnqpd1wzcYQaB+ya9l9ftmkUb2twb
3LlYkfXGsDszxJJ7oYUASfmVvet9hhrSX4hHPLrp03MUz1PN6pSph42sd4rLrpPDB60Xumw68viw
wkDJEuwXlTDYTbC8Xo8p8OSY06yRyX3Ff/6MowODwBsuq7vxs/aYOimubqqD4noNyuBrxzZdCyBF
QoKK3FObZTdZR30ZcwbnZloeoGzLAiXrmY+T0R/Oc3wpUHThYXOIz1urjlDWQSqBKPX8GTN4wn4d
Nd+aXyF2ROHh0AbaN8eacAg5wM11zOqp0M0ZGTK4L6Or+QsSyULwXUk4Z+X8Y7syx8MLkbYSzl6Z
HSjeFZF0/fJimNxtC2SnrXipHwSS+RFFwshsSVY9W0bsy2PWKO4jyIip39NZ5nxBTsP/VDPAOX7P
TK2xa7GsdV26FjdxapbYBF+PvuB4bQOG24LyAekawufF6mmffxqIzOyt58y7iyoWD8gajqQjMHyY
inqdE0mV35TZ4hZWcMPf89JkdAN54u8/gyPd+lWkAJtHq8WXUgf4RhoAaNMrUAc3b2KHa6KkGKz7
UP5dEZOuVSBtG9t3f9KEhDRDW+pRL057n667prsr2tbGD+HEiLnmKpxyk1MOEFN8XaTb1h0VorGe
BQa6ZXrtXLmIRYu6/PqI8ehLxyi9DjttQbvLiLwtdTCeBcjHYHwFCBOujFlExvvfAGqN8v12DOvs
7HHM/mqz1R3vMmvN4Lu2QWS1KFack4LXFjauF5DQs8H5rBLzRPKIAtHBxrNH7KS/MatJ3CxgpIbb
keHCgAbpMTeTXkehEGdFkbnUWtwQ/NBFE0m+7RpAtPQr8Rykd/iGyJGtByRQZgsyPBoiMhCVqUix
WSwhTQeGVYA13GxlgDe2ALPnBQ3cvzImJk0wzXxKWVpveUXDY0c+sjcv+ScyyyMe/y7AD2wnbXBH
jrh+0p1Ec1w7tyli7HevcZqacGsbuCTRLGtyRhccMLeZfnH8A9inP7KGKCZs+r8HZ1DBWOO2TGEW
CUDGY8QzcUFheoCh3lpael3N7qwwupxtEFWZK8mTorL0lVDvQcvUpbV7OP5VE1YK5t4vClIo0JAf
7qYojOQUaTfH6AEgkKh4ulGJGEF+t0Ka6HTlVB0lyes3hlpFNIKpP1bIZj7brPOD7ENX0EUqTpxe
EgBV+qfHSdlc5DJj+iS6bNsvkyISuvGa+NXns6Tf+pzSHD7Fgfq5B7pXLMSi/70TmXKUYf8e2SnW
LDBcEEg6XKzz4wU8vUJZfnt2/jpvKycOPLhzUyofRQ3AnNcUSHkjQloySqgRDeOpnAljmBlrIlay
e5DKHyZF+8mehl3cYR58KM0wNeiKBLk5RrBIrkpKu//VpO4agn8zQXYY+1qnI2barKsKh911iDEz
RuA7Y/unsHCz8aj5JbObezn9TGzlDS/SLKCxpB6W2HOCFkjApguZV5LAC59dBzHoMtbvmnY/7V22
sQBzBfRxBEVspMJjH8trCPors6d+nVsqHSK0vu617kIq8ZvflSr5IF6R8UKoDuRSuMB30wh97Sm9
mpcQY4T8JrYneXiTz9lBgi+XDKA4BWbSRgJG+l9dY3OVg07n77eV/5zlZzp23h37GoPuBIrQz+6M
7kNDtiqRJmkEWxdVgVd1KJdE+fEjI/WT21senMyWHyJRZZOhHZecyyozW2kSywR/aOV+Vj1CGXzC
8ncSLXl5Bt/PV4jdc18LmgWvUZ+J0BI+0GF8EBREhTiYW7RXCt2ATE7KdGeO/HwGh27ukn0kQnuN
qkuByfMoL4ZFhCM49ZgiZS016i4ELRFOt75SFdpI+aUaLU8ivZwA9r1Lj7rgzl3Z2OFnNd7BsHV5
GbzGewAK2EEBdJ3CkmoehuEwBf3c5m4nbQAJZva3il3Pp0CT5M8qSO599VjdI+fy45OHN7WOrAtz
qY6vzceBd2yJYPqTL5AUQjkIj/VJq7ycs1Fh3VerQQpCy24DJCZuB7ksyJdIqr9VNjaDsvj3pSmo
Hl+10cSSSd69SEyepfBhmkMAUMkzUeMBhxxEjMfUJR695+Ji1T+kYJiCgXyJr1acekVLpb/3uZqU
mSeUiGoZtpNECg9f23U4HYFbdIgLcOUYOGOOaa/StHrvfqBTfWjFTwnEsyfnc0AkuQ0fqabpKesZ
H9oGhRA4jju9lodt4qFiiJWo1f+2szw8vnWQZNd1ml9JMs2vihvtgyqe08bFHllqwD2n/aA6wxl+
hSd+uRU0L+KIukQMgRTsf+BBezELsIFVrrMGUdwpy/up00syXQjMd6isadNPlC9yK0Mfoj7nhNTa
Cmag+IiZZw8wqV3RKDmzTW8QtQFtVuq6Sz9fVKHFCmRlqr0R8optAZ2qhqQaZb3Z0RnwCbi5wLBl
Sr4dQz2rnkYfWMiLEDig+K1got9Qjf7Nr4lYqtFhV0gA4Ldil06QGwwdcVHGhRJbUBGu5msDe9Wl
r9MkS1kyljDuVfrYG+nzn5JpEOMdIBL/OBKQ6D41jcn3PhJKQlp9Cpmhe4JTqdmwOS/Ga/Y5W5Mh
vZpama1Y4AO9OWH26SpNy3naHcqStqAgX6EuQ1KLrPxQ+X69MDVxPml6swc6A5ngyHLBW2vL6kup
dpkyuEmdWc9iSE1wBVsB/k5kVplZN/kym6npZC1keEqrbQdJp+68KnYMmh7yDp+rmqqm77VK+0dt
OKpX33JOWRQ4WEaFyYOCh+9sE/c1LxFqU1krjOaUPST+qQY4owvviegsSCWmlk8aLUM3gMIrPNn8
vDiO0wpTkLLCBaRXie5rAS6nx2dircIAYYCcGE03xT4fvO2oI7UqrYzBXLPFr1A25TvgxCHOnI3x
EjxcJnS4QR+SAMSCajTJYrx+Xj2TrYI3V7CcDZeK8lQ9rRXY6CGjRTMJBGXW4lOUMx1eoVdqpXX1
4a3zKXW9SIqu4CT/gcAlSz3QdYMzRBmoh9pBvyGuhWvXN4uwfO4DntQioSLvbt7dtAtjoPylL778
2g0f36R0QN08lr900hcaBHvrWVdyvevgfTm4NdowdBCf7sgZiI0YbzDn1jGwiJY+fc6zOU6/ydVy
eb0yJ1hjdDCdT0Zsp2lf/ZwiClXwJ2BGXP4U6S2Uom2Kr9NNxbTp+AfIgqX81Xl/LXs0CRXp/UQc
ZbHft+qnRzIMJYx7SjMmEmUAsUHHhUtjDMKcVICugOmoiG3HYUNV4h+IwSkPD3i39cRlkgsHfeuM
vhP8baGk5C47p6SAmKWnVexRTFeImWbH/jBeMvS7xobwY6AInbMk2H9NIjZminbYmQEv4xuUzoOl
/gHsgFBtHu7z67dXCll9h1DGvXfnxjOdvmuJZpyyf20vOKw7AZnGzZwN01G/OZiKe+Xk7L59xIq+
g09jHTn0nXZ6gtQeeXq9R8x8X01MZfuxe++HkgPCKQ7un9uNOo+t7TOenRYnrDzqRaQHY5y2UhhZ
lMaxs+CIDAtfItyqTFqVTjfKCHDa1C5oFgOu9ZozpxMvtNIsbEtmOYHBezH+o4HlM+qPIQGGIAb9
cFgY9IU7zAf2pfkfLFuGxhBU5PxLptn/7ntYnsVMDEZbnkWGQgIPBaqK84sknIOjvbDAq4gL3tnd
7BP38jj0SCUNKTkuZEd6QWMCKlhBFmTc+fN5XQUIaK42VSDaQlfhrehH905fV866NkiOgYKPC+5D
aGcKGtPXILt0wvPU0zorpAxi+cOCd0C7gWRC4zioSbgGjVckWqbNiw7PFXsoisa+5WVHkP/xz9hv
MfE/GPDSYRAgJVLuwyziKjdz+b4PxeW8TbwNSepJ9VarcqrCuSuTfxjuN/YFvn+HwrTUfftGKnEA
KnlYxEjtsKeWBmkpcQAZPTtbOeQUvR/559dmkCczZ/xcZkhOK2GbSTihjKWZA28iOJY+oisIIH0V
QZkB5RuY1CQL5Ajhbkm7PKOMbJLFDIssyy4sCziEh9eyflyi3PZtV49vJktIHQ6YKlL/J1yQ/r+9
0sWjrzM8Mrrt2BeEqeVNx4EueNxxOB86HHBu/OP+GQmQDJ+GGu75S86ygH0PKIEmOGhkL4Z2OOTh
947Qa0yfu/AjKzsDHWunaE2EMkWQA8pNEqqs8DiYxFdlWQ05qXa5yz14GgQJ6nrfYttUxOT8Cslm
s32js7sf81vDpFPCOOiNaZXPiRnYErxiQXbSVfKD98QI1KRmlH42YaaocNPIUYtTDaLVHjDk/QKv
GKihjs/Qvb34K04cGoeSUGin3IaS3u5+AdXsCVHCoAZQrQa0rqclXBbssuMkq+weziEnskvLwCL6
pOtCvBbyXLdrH07S44hX77T4o6e4vM4BsvymUWgictLQmxgIHgosqI7F0WjTCMl1IIlM2LY+J20a
iM3KBQOsOp2iB1YdJDfs3IHArqgm93ySXmcQctVSrMO9tkIYnpYkeEI/UDpq8pRvGxnyp5zOnfl8
SV7G1trwVhcz+P3n76sHGtl02/hxKsiwAWjAZQA87BHNJ/O2+DIe4tgUUu/fH8dFhgjQQaMKhgHm
b23sE/3gDR3VniYDcTFstSVNS3+pQ+IwDescqcAoOBUD7UrJmZtmlSbmChXeS6PeIMEWdDNh7Uxa
67oQnI2OC7ZixxzEZqAq1pGQ/MBeSJIkiki7eETmXDej7d0wVhsQyOVvuvldF7s+OElReyxu14YR
GJcKC39uI9iXkBOr5Rba/23viSZ8djMPSyBIXNHEV0u+OZs6LLVEKw3biKJfbT15EjyHWRwj3yuD
TOZHXt95Rt7mVkZWG8gr2GTnen4KJXBgEB7ir3+uyUcE7ANioK4yJYIIglQW9UYIxWnF2l8/8X8W
cDjwxxJaVH/jZHCkO6kK2lx8Hee36N8uCneoLa1mOVpxAR6QXFDFhHqm3WTLEBGWS+6dnodpF63z
8vcPvuMqN49N3Br0gEmrk3mGzEuMhC06GO6uWJXvJKikRTT/0u4M0CIf4a4XeVVLYuy2fddBdGRx
SwsqWJjETTgm5vcxlrP5QpGw2WBwjAFhhsZGReE23OlTu9a4BQ9JpTc9c1lBFwJZDw1+/HRblIst
HaeqraQEP5LqdeDBWC5NmlFKqfTqkwRn/6O1aq3hnIoyCK24cIBpYKhQ961KJSK6SyqIgTgoWx4c
7V7BiRjBq9L4qRQxuyuTqC2wc18wuroQMYXisYMxUso1IkmRd3nZ09pBgFqNc8ldwLLIAVHmTlW1
9QVN4T86rn5svjhspxB2J3yoDi77w3spoVotpRx0EfEGZpdT4RpkfAHV3F07/S4YC9AFmPQOBwYj
HXcrf4X5GYxNm3hL7MxJizyCOlPLQbGAR4i26jFdXMCZvJccZQPt3FKhAwdczXndPzWxXaBUhsxs
Y8ETpkQkt26VTPNbjWiyWqDW8WpvzKRF0cVYVitJODwUwx0XTcZuYToVFI/7Tr2hfYNQdYrhIeXT
odpUIx3Yb7tyC+qtFBcgI8SUr4iaerHlIHTBLTXsNfPOUm339NjkQzO1FI66kQJ/2ZGfgtq+hqSx
3h4wd22IXbXwmKhJuXNWT7DT2WnJ/RB1XuHUkoWlBNnFhtclhhdG9bF9fdMMzbj8jxQCzn4ZWPld
G1bDl5Xep1QDObNBbVg/r4XLur+L8m75cftMcQBZqAfIeMtG0JbtGpvTINCsuaxZF54lP9xWPTzK
8ehuxRO+6Uu77TPxIc8/XjgQMGs+WtH/2WeARLoV8C/mVbRrE0e5qcYpY8dwM4DDbmHkucukbiuW
P4Jrh/ZSfstE5ZRv635aPSXNf++UkGvStt8Wwmv8Xh+Qkhqyg1Lx/eBggWamn/Y7T1CW+GONeFzj
aUPBAXzIoCKsN0EKXkv4qEb+SClEeA4c/4j0BD5wfOuMvkfY37wgr3wvzXr8WBJkicWAEcEE9qfR
FHcppLULUFM6ltkZ8E9xujTZT5AdPdSM5PEXB6AKbjx9lodW5e8gqgQt736IaMrthEE+DmJ+P99B
m35PhBQrJRwWW+4F93ZssaKG304e2WrbhPN15VylCWToDgBEtaqjA1pHgdfkOcmpkvnnxUyMr/NR
2MZRfVWbaar5Yaho7FoX1ILA6mQU8jJdtp9HlkMIFd4mwLsN+kL6ySAKgGFxuFYb9iDreR9lyTVP
z9GxR1yMb7SDkExAd4o+vRo7I4SLQTgnZNDI4cM5IWSUZyu8Vp1KV9jbQe9FsUKo27uxmfVD9kO/
bIcq3zqvTr3GKahXhwHjK8DTW3Tc/E8h9+y2m3UzVBtaaarv3AJOZwWLUr0nfzNIgDHkxGQj9Jan
JzVR3dvbQ1sEsdmdhsK0IBp//EGdYovj1RGTB559PTDET2OhP4FiKjE8ldE3NqTvab8533Ah83sq
eKP9AZzhAjrfOctwhNnEIf0pS4PFGbiPYU1BYbrTSLp+o3grilEG2UAhesNDl9d/ruwqibmo2lny
RV3OjOD84Vg37szyrx5cX8pCDV/c67y0m1xs9tKLNA0I5bq/r6KuivMhgkhokJmEMGY2v7vMHDgs
T1MiAjZzsVET8hkbzNhU4jzDbBAJdetuG8NgroD30lnbmGsN26/DcbQ1v+18lDOBl6W0B2x+LRPu
01eTfxXsrrsLdtJtOgn/71bVrK5yL5NpephprPeGJ/9PCTF4wPLzGCms/zFalBMvOYu6pcMvRVaP
Gn46oZEx9vD21fFwrl+xOcN/WylcequuSa2X9IIScri7kayikiLfxenx0KaKTjD5+5rRubYHo0pk
mqDOH5LDI5pm15oY1NR1TZqz9VKGnuSclwzrlkzUUrld0srrhTU3jBV/xrgwMN0iOsCahWIsbfMS
/YInFliJnwgg560QHz2c65pDB18VMgHWypQ8OweCcq72fDiXPKCtzcMyvmQHk6zbYRQhiGQzc+ZA
sIkEOuzDu5wp0BGeslr3Q2Ufhfo2OVo4JxfWe11jGam9X0lVfHmfabjeZvnLwm+W+zuPy3tc6Sgs
qpvjCycrL/pa7C6C2RN7awqU5+MIKSisW1frsWmSXhY+wcNdoFBKsagq2Igz/a1wYfQ5VNxfNtDD
dZ6O4aTjY0zJyecNCcQlwyZQ30LCW6AbWjendwA3OPLVL5T1kk3e4Yypg1L4ZBA79t3gKNsC6lCy
grEd3AelcFd8CF+F03TU1NBJ8Ji328kKDuaXplBU3uRDQJYSnay+0bDuDnFROxjij+J3NNgBaxvY
/RSxdFyDt4wN3Acp/lPM2B7oH8Xj8288KYSHTtk8arcc5jQegDvh5l+JpfjAdXgJwQjRjPXgyC4a
iNHumpkJ/pGKqJerLyrUKSGIRRwDPgTT2GYU4ZTlQOvwS/T0+3qdJ+0SJSkYc3otpPTGznn046UT
11wPYOpLDlJ7Y7+pacyFsbHnbllT6eW5ucodZxlvlLdBzBW48jXjLMqhJ5y2MuxY0Mft1q9V8ttC
HLfIedN0X51DB+LkqcpUupt9183k9MdEmEO33JzBsczXFvHruFi2yJPH6JE3r+r3CvgXE1p8/MN8
xAy0Gh8TbVID8bvtPku3o7kfZ+w2AhOFAy2TYeiIOq/6wUk2aAg5/o1+gIKyuoAQ1/Of2qfRTaJx
ErJlnPz9i39c/Ib1CTjEedq32mgFxO5Et0Gjz7tiIKEZM/Iy4llGIasHD4wR7IA+/iKu0yjAZiQ3
YKRtFbn2gzW6/mRTNB5fCbNjaecDdWSGEVHCGoPcYOHvuLhhEBeQ0bQnfCRYULDP1cwRJihg3khu
MRsn2YbkZ2GXUCDneZD3b5PHedHnY3veUW1vJ3/8NWOHAlLaAb4gLQLw53O7d+qiR5h19mXc3y/O
PdtQSahWlnRyIgKgwJaFF7gtXgcG/gx25RWBxkYpkJfZdJ78WoaOr9o840tYWs63Gji5C8l70H56
CyxHpGS8UJ9KGio4zCuKrsvzqUZudzrwWm7zajX8bDBq1un4yo/OarKG/ZROJWh8pt5a7NBqKnp1
fcy2fVmiwhqyyjJBHBUN8s7p2KVj09my0xhcb1CIH254VYkurBO9e9ipDkrrhSuq2W8rlYQoDOAi
StuHgxTJ6hPgfMLp/su3ExOiBBKDthg2uzaDKpJEMCF+tpMJm0RZ0T0ETNUz6L00huStpeiGsUAb
DkPVjHdnferlw8Bn8rjCSQfF2bLs6iXT4Fh7idCyr6ahFlwhQcKn+7B19hRB6qW6Neo6KvOUj3xH
aQ7Nq0zQTXP16HIjzj522mJl0SyghKsvkK1ZdE4DSUW/F8/EsJ/ketCbTsbS0k6osb0V7S5EZUNQ
rJdUxVndajbN3LpDEar6sDrbOdHOdacHC7Eccs5QHhF3viSAprTEYDNeyQgijVm3NQ7MSoZytHSl
v8UcCgGtOJBbzyTDXW0gSddKE5AIl6ydI7dNAXdeXVbAMAF6OfhLvP8OIogGBPk6+Yji8XKSHL04
Y5Jj9fJ0bf2BgP/lr1IdVrxB+0db+skHsaHPEU/4ZprVyfQLzAYgRzlxJLr4RzR1OWEgFNKPrjs0
2OP8QxEnjdkqhshI0FO+Gzjx2Y8xxnHgcpcJxuGwCJnkjn87Gl0ThjF7omXVjTsRWl8FtzCzS2uG
SVxJtxYylZ37x5lh7iZu3KEjIlqqkmHZ94sxkhPSdvOp4OszcczjTl8JYxk6m1SKH/nTDJWw6Wt1
4KnrgMUtBuXRpy5R2PhtUjxQsvweD3dQFf/Z561+Oq3DL+2IG350NOX8oVNwovIhbcwUnKFIpg6l
FC7cYQHCIwSzZbLz3cLPZZOasSRBWBQ/TACjyIAswuBCDtUHQsmoQsGXXuabwTG/r+WTt/qLL6Y3
xTwbed4lLUXM4Fxj8KRygS6Nb4Smyqu3BZFTaEMTh/juYrg1C3yVoYlWQqd652XT7FuU7kgVELx/
1PkNzidcUI0doNY0c8IEnasWAn3/v7nvRScsvn1jWPAojRLmiHKAEeYQKGo/9d3uK6xytRrsddyB
jcQvm5mQay++Iz97ViEiSlXecAifxp3VEHx03ofCf65ZNyk904jiTp6XDBNLeaaXipayQ4PU1hM5
reQ7oe3eEbgTR61BAIyQmQjuh56Dt1ChQaxZMLjHKljGhhgZSanndxLS/0T4VkdeCr38AfwDBQ/4
6t3NoMlcy1fwMUnSOgQ41FUeG6jbUhomEPEFHgY2OfGIDfrFAC5nBfS9vvzLYpkyT2TlTbovDfoS
QCGCWK3E7ryHryIJRVv865Z2GTmBwtQ8DtVLbZd3yx3nBoQox1wwaeAxUwkxycbSSaEGtfY0Uniw
RfFU8ytccwhDqkZxKAq1Ix6zeK1PzRf4PyXuZxBZNWaIWJZfLTUeIyP0GpInGzIk3eCYGlofZHCL
oxi/zLnu03xaPE7mDgxNg48Nns9hRtsbTJUIVHyrpJjMEPZ4E10NFJ9AAgqCCkP5N2ka+blEwq8b
uF9FJsFqEUGAmoDqtnNkzrIHscz9atZjgDsMMTQHpa6TrVNVS9h/AkFLIOxdAnZpW/s0zitAs6Mq
cnugSvQQmMhJMAk2Q+5GiBVv1H/KlC7y12jTnKUndfN9yDFJ+3aY81ul0u690opNcFJyvBUT4e73
IrPZviBtmpUBQMzw7fksmbW3ej4HVlUi7bk0iTNvN1LbL1mFl55RWBNZyvzp/Uxg5eDLm6R1DF2t
3LJaLARI7sAQwAZWJvBmA4Ff0aFZPsbWI35+H9wNju/GxXrwaUH4IyyQiN4kvYeQFWYexZztto09
1MGN120VovSmgBTP79VeMRsL2pm91QLh79ZDs+AKdnAWyUbVa1gn2QUGqFXiKCSHUdgaOhpJUsca
2AOUMv3Sqfx7B5UQikWHHDtCuoRIpoEPt6rF6iQdaYoFvEgkKPx4qKWP6A+4aTbJn67T0o5SHK6M
rFQMkvciWR3SF9kFM9Ouf0tkbzd94r30VV8iU+HU52St7323omZtcPLOei5pzkPonj8aU0OvPlr5
aMi7uh8fDFc3uk9v37T8INz53HXRy7WvyVj8PVjRpFovCZvCnv28ZjfSaeEWgwCANImJWzhtDbpD
RAzG/ckekJIw6+3XojxnpfM0/mDVmUhM8y1GFiGU4wojTHSBhwIAHfwxCv1m9i0BnS1XXYhXAyd1
YGjqWw2ZRNPG9m198On7qAFLsQD0coBq1DEl6AdXTG+HB6uFRbyGXR6RWVGBy2Y3CTukivcYht1F
ozZmyZRQpk0I57pNw71Tx3myqngs3NHGreMK3YTuG9/IrdRmjDqYODYjFRgTULKovp8eFo8sxHPP
H9qX+2uxVNemRnu6USirppbOf4SiHVs31TaaVKDyNt3XcgtzGshxz4pQ8HRLJOkdnHKmfGDHCd9M
bKdCzV+fZiHSIqFVaW+D4FfzjHjcQ6wQkK4Y1rScsqyIvD5lR/3u4/AGB0CGy5lTHefquXQxRWnP
pJomY1WBHV2hmf2/jT6UgGe/VpKHiJBM4KrZKsLNquXZTI3JWLMqESlvZoiGXgZm/4WmZ1sZIYPK
26RihwHURzgp6nLl1/IuWanOzbDb0kgX9IYlAmwP+xq+FqjKi7b1NeTEATMVQgVmNaPSWyCI+v4O
awG3L48/xDtkSnnxrfA9phQ9aGTUCpKsrD1FYJEFK7M/cpjp3F63XMjVPI+GoEgQNUx9V1W7V1HO
VXLjmz4t/wjTCyo9cE3UtTae1fKFxHiJKWwpY/k4Nwx2ttxO+AfonRnPZr+GJmVjTq/bJBIN0N+9
Tv/2M4QKLgCqvQ3pqARtcuP+WESVV7UbZVk+HjGfZyf9dtSz4q9NfXxSvBoVxmOnb7unpdx0nyBw
vu8LE7TYye74LJXXK8BAcjYXACdj7MlHC3eKAKBbu7z8BH6n2pwtx9DMez1OGZkJVN3g7NrSgnAb
UCqXmYyuCy+FTWFywTp4mcdWM+W3zArFdZDW+b1lX1w8NhhVdd922DQAiTj041YpXMpr0I4xvr/8
NA228hy9etahql5XC2gbpZVVz6GoXLLlFHz1LgkQ2e+DUrL9Ez4/EJ2gZ7mFa00hhlKjmop9rE1W
k/yrgQ+QJMK0alfddt3SMyQj7P452RYURgV3brfpOnHMkB6LcLU6aXA14KNUCgZkWLX8tzG9CD4V
E2AyLjjWha5chswcTsOTQvnV4aGvY6sFv9ct05mGB2CyuTgdKzgt/bglTa/Ssp7Evn6COhX303J9
PMn9sILw7sLb2GglRHntSZpfq+FXccKdt2XT1Z9XpZD5TK8cR4WDqpYU/rV/U4jT6WTxWkZbMmoL
u8VFg6srACCOUx2nya39f0uZKZuhBgYKniHmcHdvsvqLz3njM431gF2/St9GsCU5t26QCOufo6FS
VBsedqk+slMHVGsUWK2dXoRbmYyjRDuULR6irlZony75Q4WcrTjvFKC7tY92b3jz5QUeNcROvVXe
F5S/WQgP7IOPMJeYrPiQiIleda9Ugy54yNlTLCNd34L/wwDNQ3c/f6oIn1xx9W9YHdz+sbe3nORJ
goz8Y8lv8+B4abjMCKDuFur63I4fQlobYcHB2DBUH0Q6/2WepZsEpwVMr3et5B8DAWb69r92bYgk
EA+3WJf33ezukTtA+QdmsFZmJfdQNuDZYbWdta7PfBWSoPDmhiFzyB6k/SDAZPsUPnneRgR7AgvD
ZIV1iEKjvjMF/b4sPe7CeNmjkTZvc71uKvZFsrTPMfPtnkZp4/ou6pxT32RsBnqQdhtZ6rq/TaXz
OJLqkMDJlYZY+0Qce+GY4Z2NdIoBErPyjKAQnphBw6MRAj8W7FHNJ6DHBZivZGmEHMeAt+wJmaWc
MSuyIZPijYKRme2f38PQSab6lQH4vDrOCxMwR8HtToeTpXHgXLOhcuxUzc+vHnAm5sBe1c4CtHaw
X/zGd44UQMQiJR8VxCWAU3XThs5XhFFqnXnKMOc8XwgZ9XOWH7ag6YMfp3FjDhF+FvIFrxGJ16M2
4EHtx+1QLTqQBwPHKgs6Acj8ayLPytWW6c3dGp/5aM2h3S0r2eIBdTMYEwOXjXG9VwGcUtU+gSUf
wCXY/FrPwsyZ4fV1mjF7syHTSms/yQ+RKXyPKIhPTWAegWvlVM8g9fh5aaon8+zF6WuEetipxWFh
KFw+zklT3xlPzLnRJi/wnvGmKHJy1qxgky9L8LOYJqwM7UA4pmytBLa70OU4dAdJqosnVhWe8k8R
jzpBx8R7Ao/HRuwHZk4LCynmAhMkC/Wwdn64ScCtqaYUSVKWw6QeI06piNNVF4GwsxTNwJWJbhxP
jRhsf7CQdifVriLmVj1uO2rWzmVcedNZOPAPAf+8FdrFIE415Gv874/pqIEgqT215XRt+YKG9BEm
ED7frrY52xyO6Na09fpSs2M+dYlgHnn4lnhRlWVZn3E9Dd0Jd/QXrDXdiSq7oQCTsC8HmI6paSeD
GjUu+TorHHanniobw79IyySzhXMaJzQNEkxTFxcLRaKZlAfXhzpHMNywF5YcZ3RbhFNTWlDBnJtW
K85qubG6Ozig0tG50vvY4zCTyZTQQN7aKaaOnoB26yDTQMOLry5aZZQbFctjYl2Rmen4iT3SMA7i
CbFI6RS6doU8jBVXFkdaqOB8Rk/sacC3IcxgCW+QWVr8oPr1VyIdFpoHpEdr0lwXypCmgJngmqOf
YhxfKYXtyWakUsjNZQXMe6G4K30MfPLBbGc0vRC4RuWYSpN4zwCo4olaxq8DlSNOnvNYPyskFSDU
WbZKaccHtoCHS0DVTJi9+XZgH5rxqDLDRMn66Z87l06YZfSmeEkx0BIOapURNeFpA/4qIPX12jo1
x90ldY6Z3Duu70PO8czeOQdHO2c9H73iLcVbdAzNPF2RvXR+wXRpR1WE1/Du/WMNLB5c3HfYJcV3
EYSjujuYPEUjEF58Jbs3i1E8j9VWvjSbK6JT1L9Sj4UlcJFF1BKnq4NZq5ke3s7Ce+Bi0cHwZ1m5
2djfFtW4ZdydYLznaKBKTBfmHyuikBxmLkZFQpoxyYeOuHtZijBSYevH9rfLjbQyrCQ9947QuV9f
ckoUOEG/flZivqadF1DwkJzRYxZJPHsR4xqppBuzxh53Q8qVY4MMmD55lS3UHixad3aiD+2+q6jl
wcdijyv/FIiF44LOqIADdFZyJsTGSURunzucVSxvGyzg2mzBctHC41AaTtTEVrDNNJQfe5qcv39+
byUQigPdJmUv7M3FsyewXZHj765AqIjgbFROkmvtAbF+qmbYrkR8yzMTJUCPlGO3Zc+DvS9CRHBE
4P/4ZdXVMD4MrA5JmR9ZTONRClHHtAB1c5KiuBvWtoXdTCR2fjDjjTakicaPjTjfpfZ6YJpZdaua
OXNvyG7Y7TfzaPmNa21Lcos/ISB5WONkmk7cpUStE9kvQAoDCipyMtA1XYu9v+BRVfQ3m2/IZ2pp
/+SFxU8XpvjjnDX61fXrTc3UXt1lBtZDf6EB1yxXk1sX9EuQPJaw1IvsPg1hNVhoikTDe30gjT1x
P6OMw5x+ot0lH/Xnofv7/JlU6lotzBBMVSUSFLWqEbqtwJw8Xk+rhhOr3kyVlFnHnMlKGC7wrw04
1SOVlIoTaJ8q1rvSXH7cBrWiULiFYBqaWaYeg4VsC/jCzhXaHkpbwDTLCrsibU2XAgphgd2K7tLd
RiPB17PonCAt2oY5SPExRBdtaBQqzIGS/ukJRgaB+UaTtwTdvevR9KM9g+GMVf0+qESO2TkG5NZ9
cvtPrLJ8Dj2lDH7PQnJouxZ63ivcaKE0BWDGpUvbrF/pTsLMQZzuArlilX+J2WeYKi8NOQ4aNCVC
aMmXK8+4ZNQjc9LgZZX4Mr0wsb5WpA08O2n3Nwyw0XaDCnOnIx78KXF40CvrryfgEXgYo66++e6X
SScdzp+88WYIzPDM4iwd+9CoJ2k+6JyjLJ9hMIDzVlRSjA1cQExKSi/FPFtY6TJ/ZUUA1dOdWwWX
NVYAMl70PKVFflR7dSD05pSN4s2f/ebWXpsypNPPKg4vUjtgeunfQb0+dRYs1+as4ggirlqsvH5H
OAt753noXpzHYAXEXNHGvH+WrESFz9z+uV0+ISbtQAeN//X9lSxSnlnXu0oeSwOqWzuMmK5ng4bA
gRxhFvHI4FqoEsooJBreksc/Bs3vY74QK/qQKeY10XPfZ8PMbxltJS7TkF2dYL0fZvtyZi+clZ+Z
X/B6gwAZrmBKLaotvyWMFoFpAO2YgcRtWyONvEZLEdByWpfJxm58jmPV/9XOYmJvGtE+harZi6pC
SIzzCmta1UIDwJRP+TPDsPg6uHIjtCKT4qqX47zLnBCt8ZjWK5Rcw7Oy/Y6H0vEchy1o8fs1o4E/
vI4LThSPZ/xs8UupncANoli45j3njGo/0JZb4YgKbQaYjRyClb3AwqoW9A0GQ/XIDoD4sSUUg2MF
FXHYxlZcjP6sG7V5jpXwZTmOhWATzHOwBcm+9I8rSoWGuUtHib5FYhrq7wqWSsRJKlKUwZY1tmC8
bl1h5SK88k+sUI2MtZYPeyGph9cQu9Ur3p2ziO1mAHT7apoZj+bmo8rT7vpOSjemrzwqoLcIUSmv
eJ5NefYQGZCBBMwJWgq3gBuNgPlC0Jd/L31eTFiPDOOs++poKGJLJIZNh3H7aHvK2utFXJihLEuD
oAk3PrxOI0XT3zvvtHF81RyikVDHO7q+MGube5DSKado8EHh7jceF4j00Ygqm1F4Z3UsUF1wGTs6
IF0k7SQQmmp5AUrL/HKdGDmLXVt2ryh3JcNHgXlRBLaSvQ5dcJxiZkW/8NTdUiY/BbpGxoNcIO4R
G8O88rd+EwREYb4+YSNf/iGqHKbD6ATXJH8P0qbONOzXzRHiDhHlXpRzVBQgQ22eSpgmqS8NXYVf
gabk1osFQDmdpSH2uaCwRfDTPxMEah02mZAM3ZpE0WeJLZQvmh8VBVwzbNFniuMaZsXuKDtjlVwC
Iun+3ClctVlWlrhxBbs5fTRWfbLjIBdN6mxy/q/kTDaXzoAcr9dE5o2tU9eOC6GDgp+4ET1RSXA6
qBq8E8SD/5jwXMHEYQWPjgfyzZAn39UxmyVv+Pcsryde+S5YX/eLxLyssONxLbGSO+CATNCMDn3B
/eucEQovAjz5T1S947DkHBjTalwQySRp9Buhz2CKpIrHHBk3rZ7RBsTdQ5VSVSeHjcNuxxpFEwaA
mxI20pKkkxnqTCEk/qKZr6ulquStokJQtDm3e45iU/mUcoiycnjTbFrpiwHkY3bzKtb/LnHH+4sS
hQOJxNG5SN4sJh05iyk0wNdOC3geAlHfaNujfUAD4YMQfcuPERJAL7YuJyQ/hpRIvfoRlCvsvLb6
EXymNoxX77+9u37vKE1TN6ZA54g6VofuzF/3lE2+fQWncHlOT1hpez46ZjpfRcZ8nhvez1Ul34MU
0/St8StO4V8LLS2YkxzZfpDuitYistsNzOHGpANWD4imFHKbVTVjghJslj5jnXR7w4tYBFj3BVYq
cGdyO8Rc5G3U/JLgpywJFKTFS6W8SKhTMOkNJSRsLAt50NCDRPkjwXfbIj2dF3Ey1tlV4/1iwqlr
KjR6PWpd2tdSyMwAc4AGZSWdeoZbmeQjGrfEB1K9dxYoYAo0nb3gbDU/ixJSoBuQPPKp7eyNXJBH
UtXg8Gw4p9jBJiAQ8B7efNRmYnvDc9qOJBRv02/i31hW9Tn+rhnuoXQ/wJOftpfhr11QArqFjMMw
GB5AOoYUczizpGxGT2EuY2BqgJWjO3qAt+pq2DCNvqXJ04ZgBdWfBe2YY1LVrgb1Au/Cgd/6jjtZ
JOkM5C75ixJuoKL8XGp5gzyQBPYdGGXC+k0BuNMmrJ/pTRqDjNhWSqNb3JAV3diX/nSTThQL0sDl
jttUSePVwTlXfjs+8mfDED/f9frLDX+3YYvVroka2VvFK9EG/bDfHBnHEJ19PHWWUVnyq05t+75y
Y+lCj0JNS/jslVXwOOMz+HerYvoHnJy584JpRmgY/Lrc0bbuEniLT3lTrIVA5Mc1TQ1s79D91E7y
WChqBoN7+BYwRya3Z79JWHJbDB7CKh6Ez0ZodZNPxVrrzJ0upCf6W6DRrhsPijP9i9/tr7+c3BBi
pjpdR/da4m+jZs34jfSiFD722e9tb83j4uMhkORBocWHYDx8OQ/DzbeomRsjUrijqR2gK2gCuiaw
JoQ3tvz1uFy6Wa9L9jDer3bo2cQvkyB0c8762StYLn55LO35KZNBJQ2haXnt7HIDL815hNnqwfAi
VEuJuS+JatucyfZRISOvltOayKB81lWs+SNCngd8Yq1sb2OyiJSaJ/JMsgdYmLeKFqzxdBYaDC01
rLsLGRv0mPCBsTuRg2afT4CrGF90h6GxlsspHwivenNCIqFJ+nihL2VqixlFsbCoDIqoGVLCaFna
ck08Xi5advffjIf0S3eiH4R66sW79OdvUDCfXU8X7MTvjCNJlx3p1Kl2p2uc0mnzpd0jyW4iIO0Z
QSMyGCti7LS335TuqVLIxuE12TgDxMo7FPm/iFZaeWPwwhRR9HEsGmBq6+fG0m72+0Km71+B6CKy
WfUVhhLMEtTixMFps6HN9buq7U21uuL+od56mi9IFW8McCVRF7Tc1rhWwWWJY+OKrjYD+HLHBWDo
da50feQxY/aQym22YlnMq9AfIuo236hWzqm2vsDSSNSbMNtpUSGFSqKc6XeMaMmW1t0GwfSvFgIV
rqadrFABEOT3gRguz005076/Zyk5bxOC9r9ExUMoUek7LTHgZEremmPZYFVJ5gk8POn/d9aiQrBq
+bIQRehL9MtSZFRY2CPVcRAJn5HeOLifFkK33jBulWQ03O5d3IV5CHWouea76QlE496s8uA4H3H+
2Ju5u8ItH2NW0cXicdto9XFzb1wecUNnUWsAiCAulgFT2XlHq2Ohk+S/IpyXeFUGBjUa065TMwLj
k/+sbKqxyF/9G9kjgvuk7HMc7TJdPCVtD0jytO2HjrviGsiAjVn7cMl9A56zj7QmEnnloWD5npy+
OCTQ4HbOxSGeM88TdGvLfZwBu3J4MMBkiK744AQW1vwkhN5KfDNY09HjYZQzqUxJE5x0DROdEZPu
iS0ocaqNxiVU0JC4arKW4mbZlJyzgqJm+4dCR54Y8Fsijdj9ocpOSIeUzuyRhMDcDq3KCQmIWyPb
QXNIwHC6XGtjXo0PHp5BPlnXkBT3dxHrxvU4IydPUAf0CB2qFilDcUVro83wXaShN+euTkwWyM4u
yuNV9C/EUQrEwchvRLGiezzKGPaYrDitZSRh0qJj9JH4M1/LzV/a3LX2I7YYVcYowdr67PfudrQx
0X+Yqtc741t6vWSLmN815AFYuXZtJtMKAFuxVq4nu89016YS2DcYaspuiNnfxGDvNuORURPrh26B
+FPG+vXlR5quaWBa5wFK7sGMPMcRZp/1jI5PXCYafX47lRJfZr0Z6szvM5bwHEcnnzJRV2TOwyAl
dlNiBF6vBhHRbx956BGfL9YIBWORDnRUcGOUQnHyBUH5I0blkc+GZg3orpWMKBVhIlUv8dwX4/Vs
AGIkTN2/q8rejB3nVZ1jTF3yYNPCBLvqJVVPh9kEMsZwC07FBuTEp2UeEc3cHsxnjoWZ0r7QfnVu
ZEOMzPlbxnor1FVbpYHOlGGG8uei3NSyPmYH9P+fyE/6xYvu37SC5NurQuFMfHxRI26VcIfF2x4p
kCXm3jGXW1VzOeuXUilQVBFrQYzra6mjlN9cbbtalYXHuMUEJJUotI0b/UQyqCM6iGqrHoQzmUYj
Rj3DlnZsErSPkvlRS4xcJuDwuWsWKPGnVAQQduUbPhyoUdkcFSmJHMPfriYM52k9DLQH3SRAbF0A
E5LiyrLeAfBCAD2kaRHR70fktsy6m/nAqGzOueSyCgNGrx7w+3lMi/NES5kMXSEISOp4HtMXlW6s
MuinOA3LBakJWbZcXLsXM5IrDI8AMSxwR2DCQsNGhw9jTsgeH6WWtn4aBavO8qE7HsHCXISGZ0cj
GBm+C4qU8qBQf808zPqWiBgr79Kxn6rKCI7YPqv6mkfZDXvm6hI8rlq3Bf/q9l4tE/XNE585zHtv
k5oPnPgv+gqf+5VvSp2xdcws21CDR/s2vkch+uo6/xvkCQSxKwxtO2JbMLrcd0WgOsNj22rbJqDP
a1yQs5VLQ1QAbXB67AAN3yEN4M+SeY3VCWf7VRiHLydXu6LpCUKJCUyV98MQF7SKXgDWK18iTEgr
zZdVZXK4v3BeCzbJspihT+0DhSX/PoQ/kmewTisFxg9mB/tkGJ2i+SkkImDLiYmc75DrXpunAky+
zipCVvQR0dUww0Z4vwweOZFtVyZpV4gTZD4fQhvzfyi7okf+iQ4eisNfnugiC1jHtpMDgd6Z8qmT
ostgkoAeuykM0TXc1Ti/WyqlRSnTQbZeo6T3CFb7Oiy2Aaj8v1iXnmkZnP86EpTS0UgoBmdZ2jhO
DjDqbxbNt/P0nV1R7Rfuyik8Kesc/ZvT1zUylVXe9VoAcBJkfUgN+q+VZxThXE9OBZQX0RNnBQXu
PMdWyVIZOKCTpOyGJCG9wsKCFvLMtoHkyTHXQSg45pO/CUgpyEVIO+J/Qh7SCMtyIg07e5aHhW8G
m51SEUBcovKtSIt0xjShkFVkomAhIOqLTvB1zoeQDdd52qvv389PNg88k9o6kurZyfm674+yeAsN
v5auddWi3LcZ1THuF2meymtVogf6BzSatdxVv2TZF9zJXpjxeU/viQnpQjSbe02aAojW6JgQ1vnj
eaArAyYEdFY4eA1OzA/7x8gRbZrfBF6UbT3rud236lIfuBJlS7QHX3oAtelOzlwvZQe0H8AVLuUh
gwW/W5l4Oz/WghdDK3mnaDktfWouB906S87mSDE4uBKRmMf56BoTpakgk3MNmO5MNbBtWhbagl4d
uWF4SCRdzjUUJmz1hsV4H64PJZtOZjvqj4MWrD3f+sDnWr6fyCRYg3se7DsbudYcTr7swcvboj+3
DgFvQ8QBmO9wfQsiQbovFlup/klLyUIeYhAvR5zi/uKBdBswIhMdY6rmoJEi20apzJalAPHsAAdI
F6Hfx5TwMB7Wjm7U8ZmRJPFJQ5C5Uoqxj26ugMP2YoeoQQZzG4Q+UK+QVNBUadB2SU2FrE1d/iY1
QCYRAlzT1sO0jpb4gAZ5ODfXvBQqKyQd8Us/cpclPQ36Z1YTtOS9hxHfuzdezNAajeDsWxCIIBid
M79vl926KNvBUBt2JWrd6GcAA5e19JB/WQ6KXWwhEBOPlwugB2wL2PwnWDiSDiQeECZ3vEg15NXM
1PRbbNy/EhZxp8uwDCyVDUFH5Hkfy6kGGHdL5S1p7V+6IjD6RI/KC+3pjrTLh4ifOTeMzWC5xapM
7s0yIvPt4aDzEJQUxOMEYV6MMr8tVNPppDUrbML5MDL+577C2IIc9Kq2vdCFaPmfnO1wE39Vv63k
N2mF4a6D8qGNmwkBnAx+vRUIZKSbLnn/lGQh1CtzIVsgRuudESwJs3gOCjuFaRLDBpQYDkYNcpOF
MiaiGZZI6ZKgFv/7niYghnbrvXnVr0+qKItp2pgAr2UQgW/P9F1wkqxNXfwE+iajM47ko6aVKcVd
hs4uaVekQ31V0iqwRVbqKjk9XzlDZd19loQj893vNPmwbU2owSsZsS02YuitLF2bqcQYcHY2fpOp
GoyzYPykUTPATfUaMwMH8MUwl7h58EwZmkolA2c/WlyhTgOqqJLGLd+TNjHDmfMTKgfzbZHfa3UY
iWAmK3Ykgh/dQgzidI9ehZ/fVv9VPpnxStVCcMnCtMVHFZ4ArYJWJ5DP3bepygd9Qj8uVXFD5sfJ
Asa4s6wyMpHCQP5o6vviyNjGtY8SKwTgypLWmsHrr+yGv9LS+ChbkFQhVfDn0DmmZsWoJV0v+F+H
kOlu1kA8QcsXgKN5zvN8G9D+FAPm10JW7mk2vEv3ZauuVV4bgeOhHlrYPgyxKFqbAv2NOU4B+s5u
lrLILprE2mC7I4AMAFzpxqXsjq5Xx4aSeEMV3ta8ndDjFabSpfKPhyA+eNQ4B1JUoIO+/i9yaYqQ
8PqKWDYPtikd14ZWow8m8FUOqzbZJseRfnA0c4FtIZbyylbjl40liQSDYf5qG46jBSgHm62DpOA8
89AdXgtL/HiTYz5M+j7tiDsPj3XU+FbV7MlnB6ceRLVv2PFdYIPNqNm4URs/O/4zmI7IY71I+B94
3tCft6uIsqLqb+XwRvjtgAZqhwhgbl5U5UVW0oZUN2QjXxQ0uTK/O25MmdS6raOrehfTCl0P+c5s
laq9xTKOep/uKombIJspzUjT+e3c5ZBy316AUlD4ggjBBayT6T6L3+NGh1dMD1S7ed6AfGisq7jF
fzkBRYfHGsR0i7xBZ9QlHunS2xMwKrl5n49M2cv+GwgnzP1X7fu9UJRuMWPxOEw6ZpwN6+Nu6/d1
aKgaIWrTgAYi4xXemw34BJzp0HdWKZS27h+N+d4ahQ3nzhyNRp3yxe7Q/nZoGeAk8FNQj7WxXTuQ
qv5ObD1XBK9u7ctUNDDCQQkJlTU0vGceW92M4Y8OesJl1fgk1vTRKp6F/IKxOprJuh/z8TBi8+bG
lngRlT8fTzbaRT5km3PxA7rUqYwT8ucETmnGBJdM3JxCoy7f6zuhAm/1JsabEv7nIezrWu+nNJgk
vALmolOpIARdJVAcN4SgSlsw9IP+W6PZ4RRXCvWAlBWuiKXq+s+bmSggjxGMCBgM1RPUKwamcGZj
TPCl07RPnVsba45X1mu6nY2zbjV7+JldBxP9RyEvcf8jI0LW11coB12RJeGDpI9OZHSsyrlBNpaf
9qR//rOdaJdDcoOu7fBm5cLhHoJcu+SSD9AM1g12w40lgE5HZJvFGAFp7d7dhwG34lRUAODiFCVb
H68VNsG4gouVMxeVefqWXPajKqzs1QPv2r9NA3elhTHpYC2pVug/yY8ekiP1k1bEgXPlT36yZJUn
z1HkB9Eic4jVumJ3a8rlOtX7zL3urbkCaHB4icB5dzrj8l6178q2NtRQarn4+qvobP2N4dznarn2
5clE60O//khPr87IvkgmQWxKdViL7FZdcheX95w8HUxuz3NRTtoYMFcqxUh3O1DUELwwmmgp6LhD
fAaOFUmGtxVZr1wEq5poQErrkOg+FngswFpJFAulj/s2q21Wr9KDEPB9lLqS6oeZFwCkoZv6wZlf
S1ad719YHoInSs8d794XieZ86u3tRIQ2L1igAnngAgPXCpq/XSus4i1BXp83/1QAh6rOADvR08R8
vQTAsx0K5leyhgKUrxw11VOHVjHkvn+0ykL2TBOGKMGxcrVNXzxImyJyrlRBujQpMWlIJgj+rsJD
k5LzD8ZJgYENJsCXNhXppYcl66UV7nNfdo1OvEQhnuT/V9b9jlO1JAuaIzYl10aWW7Bv+R9kkc4f
Iha8t0NACFrYwhPzR/U0R1IrxV499Z+k00VF/dWVX2nKDYw6C4z+4hWGrTfrANo0XV+hWkIl51UO
SFV5HhBM2N2DWtKyHJ5T+XJHdRevqWjTJBNShiUy2dpwcNkhuAXfzYI1TBF2ipUNUN6EcAHqv8Uf
dhnvXSDh2nSMSWETIdvsXN2BSDU0d+nX8794zABE6IrqRNIj8okDIztMezU0+JJ/gDLPMYPxhidT
c+NbMB6B3XPzxT6cihTUiuffRYUHjqQ8MEr9cAFd/wvQL82pYDJy8uAN5/N1JsgDMsDejLQuEP8D
tadxzQ8iQdDPnF7g08nVK6a188h3QHbhIafLO7i2gj41MKcgy6jLodOdlUpzdGLcGdgAEDEM8L9R
oPPsc9KaqME1gydSi7clI51twZpS0UjRGZcmFxLZhlqPSFiksYJ+zZ2pPMDHkb3Mvh5N61O6RtaB
IfVCfsckI8G6SUt+pWvKmZlKoKpdsqV0FG0vmoslRSxCjw+7wd5n5b1EaEumLGh03+v8f15I8SqE
ljH4dfJWRQ6nG5TEePFDFZuyRybACS7Y25C1oIOKwdFdERdDr+8n+QigWLFUGqgszCLwL36eEWSG
NLIGcLh3p5xWyEy8ygy+88kBs7AierguyYRgcay1zn5uizi8xCq5xKP3E1nFy/oNXSM4In1HxVBp
7mhQE5JfnO1IpTcuGJdDHwcXFFLtz0AhE/5lVeyrjN4+EfRsvePmGQFZPveAZvQEtbAQsPVgxkke
/QbQu0mGvcMMLBBKwMM9ZBeCI+rXSPmDdc9o76aST9Jor0yQIgWbYess9zWiqavHIS2VgUVqGzt5
qIGKapS9MpMr/Xpc2SGHTBii8EJquRTsZxegN0mGffLiL3glzIKaz9USApwhME5o2KqQelZTmCGL
p5EnG2oQRgAVAJjZ1Dj33v9tBNJLuANlQ2WePEF+x0bmssdJ2AV8XSQr6bMsACs5riaEaCAf4t/6
t53cXSRXyZQ0WWd1OXoaZvMJFgAFHUdhHOL1C3J5z3fs0Qyb+KS6hRTuFYMxHeItRfgh/CuqAX8N
MSL5zGaO6DfPQqNU9YK7c+3wH2U4VS8kUmFamTdQn2ahtqrK44o1yraY6dtSD9PH6s7AXoQ85nHK
doxiWwslORUK7Wc2ASXi/4QyE5wVWqUjScMJAkevBD+iGtOFeN7Hh416PXPDyVA4bg2MYRofxLEM
uXVNdvMiF30iI3uWDilofLFYNvFlYoM5WixuJzacsazi4aHcm/P07hD/0TjpN6mmOPNQZT6qwwFA
+3e/yifC073bFEtTLf1CHOR2ORBRP0CizEhRZP3ZJZloi+AdjocjEMNg6xG7bPkjgXKr23co2q7L
Vhsjd1qB8YNmi4wM0xe+ZKxgD4hjNyqBV7D0Pwivi6MjXHofO8bDKUGnKjyxYK6mXCW/2DjTsOPM
srz8YWp1HEJJ7GeaBXH/jDTf1k3Cw6IKOWuGagmImwLt3kJ2S/jE6a0v1deu8tIEDu/9xIK9ifY/
PVVwhE/hWuV9eQF6iVm3YWwbYwzftY5FR7Jc1K5vM34se8Be0YhwLTCLdnee2JL44LYAl1WBrJN2
0L1nGfeVd4VzdozhjdPYhzCdf4TtUjycqqY+c62Jo/lMGdtWXoXjDja+UzlnFNalqQs7Jpd2hBNF
+1h5yAvmyv0eroNNZ56kYqvBq69Z/Y0g/qIRM8M6mVLrOZ6RxK/kONd9lN+X89ajsfBWwVZ++Tnu
CSVFRLtH01sFSvlf+B9dCiksPJL+JH4e5WOIZK0ZZeZns9TV5i8bUha0TGO5Akexb/vLJUzg5KY7
qUGQ1NDg0V7QNmHYrIIieC9pNp9vVk+y4ykT/3eP6Izt+UYn6xWAuGfjQud44NbRIoMFT8HdemzF
+u4b+PN3ksBsppyy7saCzvWkbEsnhNkIrQ3pbYtdeOXpbYzjaGLAO2pn0BWVhctMSZtGDPC//g1M
dEZyj8TJikr/CptjDeAgdaA7sVk9LmJnXtBKYPxcJ4psLJVaR+jrEOusmkXr770eNCcJPSvrQVHg
Pgcf2NzE+uU4JIAEcc9nJ7Emzd9zG/nPJYbl+ANIoe7lt1DGUzUXEDjthkdP9ivAA2Coemou4R/B
A9IMTm5OB1oF7WfHAeOdSaKf/XblvkqiAHGd94Mboi9jZ5wV7KeKZRyS8c7vJG4LhLhHaeODp6UY
Ua3E8NrwBLuRazKWq7TxYfZwqPOCRirm96jgbVIxQA0ByIkmFfv6eWWNSMONWVDwlokN6SxfAhg+
c7+Dbn3nxZWGGkwQXt4/c7tfgSw02xA7I5R1vJTPklVF2QQDfO7GGcH1hA90WXcG6d8Zs59GgrgS
kGwJHU0+ixeaHb8VBGIyaXk2SWdf2Eo9W0f6SxMfSXk+lsO9+ns0Me/B5ZvAXiZX8cjhP25Gsy0p
BYFyhVlywaGtOSMtej1xwQQl4KEHaXUKA81XEctLzfAJWoftnGB0JRZkh/ymMPR7VprULNhSg9nV
/AT9yzeUA4SXCRmAhNGh23psoaJ4kUqa7sfjHRQxDMW8+sBKwcjMZ6+kHyRMpkrTHAOq3kQKmSIG
tVTHBQTz8R5Gp1Ujpyt2cKy8o9M66vm7DvGEVqLSHg5tYVmr9zkx/LIiBadBqTR/z/zjQNZAy+GK
AlUxWpBH6Hw1xcHZnDK0wP0/Wna1e5c/83MikYDS5yhMUYuZclDly+/tBVPnGE9Wg7Qd3soRNApr
r0bCLhsspwWZmBc2SirOwHupI6Nwn+U6uCnkXIUQjCB1LX4X41e6ait2f3Toe5Se1rrk6lN7fEva
rIEemSWD1/2yTVLHo9e9PMEY6dPUp9F8qBw4suMaAJmVAQunM7woB9aD641fTPsftKUu2KXuNIXg
NzxVe8DkbV4QS/gkO15vn1R6kqr5Nv6vboXPO7fTjzkKLfQm9+vKVqXm//8WxnrttBgRLeCGw3Pr
L+NNjVohieLrSiM2HsOgMy4h5VxEvYFpUTA0hoviaYzh+Bkld72cy22WHuL2zuKHoyTdBGs9toyx
u02uYx8TBTZUs+kTwAn7cTjpBzKc12PZO7aupli9cJF9Ze6+QI1SDRQ/b4AbtvNkPbU8mj1+bS8d
qyAv11V6pteYIOU+qr+gvh1XVYpD0LdzMdn8v4+coPZFVWDTFUQY/hP73PrfPaDoTq5Z8efs72YS
/TR+LvdYL16XtPzi2bgZVUssKWnkCWRtGC1spi/p0CB7aYsWq+3c5LVoma4QC4hNj/nohlvrbX0j
xaI+/brZq1F/LKV25coHNUxyevFReEOaZqr1FRj5/2B4zEZTahbYt2zeggahLG7IhFhGlE7y0fhn
wcfjqbqL5Ewn3FXq+Q8GMeGQQ8HDxMQ2UvDVfDMyF0TJBSF+OTkIsM8gd9Vtxwdkuk/RH5TBmM3d
0rUAaJIbCgHo7XfnIxgLet9VAos5LsKbpKHE3U0ypCGjMHcktNGlLl74JXQLDnluPeFE7e/3ReRB
5TBKok4F2Q727NIZGet3C/9SnzMqKJiOZn73mzHM808EV0WgbuaO9gHYU39cmSlp6thE7kMB2ine
JI8Com7AExBZUIhay6u1U/D/VvyNZDCd5JhGIlTzmRKcQ9mk5/G0gvdX7vh2HrMhGd+eeEtA16e6
ds40z+i7tilK5KkZ0Lwi6cPF/fuvvBVxyVfAi8IR9J/1b5m94bBKr/Z8imLoyjMkEHIlWP7Czbsy
f6auHeV+Lpv+MGNJoS4h/v+a7fNARkgSs80/SRBNt0mdpBbEPq39aBiqg9hYQXbPJPYrq5WGs4/r
tKAMOTFyHRXwuKYphDwd7sOb6ylvLv0twpxI9RX6DS6/9gUAO0Ge62cBA9miyL3yu6TbswIujcfi
BVP/HDvgX8lGdHCM12M1b90/INgWuHUnNRVCHE3ee0zimZUND3IpA53PENozAW/rkCPYNv2ftkF1
kdXvXO/2b4AdHXe1QiAxIPtScpv9CkcSOTd4t3gqslq31AyZzIFGl+FikqOSHBZbsIegfCyzY2T1
8TJG0Dk3M0zGTAZaHHHG2lBvIYUr2Ii+/NI1UzHg5bfEdvBnymiBn71vGNicdva/WbjF5IKCSvCc
rX7riVNZEm08Qtxk7tftskNACIxVcOQwldEOE8+KOUJzmddkbRdhg4VAjq9iKyje2GWmUHfa6UhD
QIdNu4Q7fgQNNkThUzHS7c4EdIf3jh1Xv1SknrlSuqhHV36BB7XvqGbMkwIIqnT0YVaPrBarFyq6
xDzmOGnSuf4QMa2Zu41euk0S1rLiV3SJimMi9298X93/NuSpSviEduD0LgNme/nUkWdxlfFuSPhu
OtmxvSUW9amfnHAY8ew7BQMC5H7fyxvr4aSJMS08k5pXrIZwWYrEsjmjAl4QsV2oS+GoOFcY2Kv7
ZtyTbv6Hn60LzvD5Urk9c+3krMFOd/5mLKQ01/6GQd6124ufjw32RpkcWaiRGyasnYMHm13QnQb1
75QeCQZ4565tnaRI/sM0tU3qCtAo++f/QnZD9K/3i9eSHsekY+30svDx1pYqwj1VD8soBZXqj3C3
/P6dDAqeWKfyN70AkC/xO4QNxeXTDO0IqiQs6C2KfUNMaqYYRd9poJS7KNpecm6tluQQ076g4iP+
lc1KsYsJ1InOu5j/+uiZRO5VfNpY0jQw3EoEiN1kik1tQ6wYQI/JWRzi40B5xlGW0I+/DidX6HMX
H9iZXTHg12xqpKXfuy8uk+noLbkn4jbS8fEjsEquJKOpmuOZ8EoYnjkcong1TfyO42r78PhgPuJi
lFn4rgGGVcrWyT+NfvohY/WC5oJ6V4bg4aSZkcGlOSKZZ9sZy+ceqXl7Drzsz669LTxwsuCg9TTg
jL8GBk4b6Tp1SkXcwwj+GjlevBuDyTc67hAKUrSluGwQsmRPmlvHl81j0GoFQbB2+nvhe96XzU4m
EqBBJz4Qwwfytju+1g90hGfBz51Fki6OVf7MV7igXy377pyQ0QPbUCXMlkXxQjKsMzToyqndaaXo
4UoB26zk1zmSP/cDBKMxCIdUOCQD6vxN/CWpdpOxPNUtev4MjYyFHsUDQ6LjitCNda7RlCtj8U5W
NlW3xKOqFPzrfSa2zvjROvoYdpzoeDBFz1/nPb15pChBHSAoSuCTyI46X4eXqj6gLfa3LqSLU7SO
NezQa5B0cWkNrClekD4tbGKjSjcuc9ncAzI/+0bgCDZNl/XK4u6aV3Dymij369cEogVXbKlAwhLP
rhv8O5MRrGqGQBiGCDrlFTCN7Rxmef9WZYo8ZGa8y8TAxPIa2A1SqMbXF7phAnKLarfbWL00MESN
jpaofno582v06wH4X06ktHV9IT2jvcjVBrT8Xw7DwjitKeUOk14ufPwx5U6UHROacLtptZfN/atL
jvMl0qazFjm7UoigE5nr7gIlvxwcAhbRVs8M/Rd4Qz0BX2u0C0UzOMnbI+MU98X76KqpFBwaTXn6
9QjPOCyFnWxI/CwYXYIcV5U6IHQQdlZThPCQk+VDSB1PKdOBghX37afdxZwfFSM8az5F5g4a1lWs
O54WaFo+OBkJwqkygFlwyTG/GNmaUiAFHlL1e3d2fjtBQtWJaZjKrv7ElvNPskh3asmfdCVxw8ly
vT6Z4OPm/5MLh6smo51z2KVFQ8ZAJvyLq/T6/u0ZWBzb5G8vGW8OAD/8cMXqV92+CGrsaNwJSVCS
MW2aCoVc1mcTL8pCg26dYsbBYwZkAQzjzt0r0VwDiZjcdG5FfSfZD1xHoCIKd41dPpPuZYw2grtx
V+RlFm6V1gqdKwJmq9yS1oCY+5l45MUrRWBb+XM8iFLsUT/PyTM7u/FW9ZnVMrjhnCti3Yx6imxD
S1hRpNCTYNTWGg9YwajVLu4XF3qSaM/h6xPOxtVz4iB8XkmZ0cdYM2fJLmCHDfpYISDYa//AmtV9
YdUF1GeozVd0SCo2KOX0PHKhrBI0oLRugUalFNeIvwrVempufaJQ6gN0d6d+u+m3J5iIftSTpYWe
Zgso1rGD9wOOyXEvmV4zqRmhAOvdHpYWQ0gmxZwlNyP8eQ7ytyGPTRMZl2ir8yLhAyjnjI2AkLkI
/GMAtEE3MC+XSaKJsxgPtwBjXdDm9d0LKI7DY3lC//P+JMNqIKaiD8aEuHlCAt5vly49AXqgAPRq
yLgsEan6JJiK/LQsL15BFaahOe1EdOmRxM5kyhI2sK7EquIXts5GiMB0hE0VJ+gtHwGBtKCTMh7N
vlUeFFbMyp5kIBg7wb1hGqW9CEq/Td+zPgqxNquWMZ9VZeDT74Sebtsu2RZCrZhNN6SFRe/e89WF
1RWdtjIdp2kCWws5wV22qh5+r2CZ/FFSoOkkfI9KLQNPIU8cqnyJsDpl2J5MboCkX7La5NwDFGJV
O0MV9JW7p/zloAOu5VL+p9sBrB9fIcInbiaVJwdOtbN5BlU87aGUBTu40d03z50N7X7V0Oly3S2m
Zh6guAlf+lp8sUmlu2rY7IEZZV4/79h45dfj1zJ9vSHkOlvNZ/sqoW+5lBmhs3Pc//qqgMQl3k1z
Qndk0bDD949euAvxB45ARezDwGYy4ZX/eCDmQgflAo3TwjEkOjnTMBGdnJDHMGlV9riYKqmLdcdl
deSx9nwVEt+Fg5hi8WV4Q7DGaZ0uofWH5p6mNkIdAyjDWw13F1zxkYYHzX3X3QTpggJ29dDhtfRH
O5tJvFe0xzVn2Z0Hh2JQhEQgLA3uWP407iwoOy3o/xVfPnDFVIOBk+YZkcUSqL8R6SdVx/V7CsMb
20xrrMUs7BbIjWdUG2F2YKBQX+T2Ls3YlnKkPp0CXkmUTz+U5w/Ghs7nGr++f9yZi6vvefo15y5O
cSpieLWATZqAnIQSPk/epOX3o8WUgwiNImQ+yHPCCwJtsI2+Kf8dHpI21pQf8hCTLG2q2nm1f/QC
F1cjWzFK7WB4UZq8I1/10za0iEIa7fvPy7H10fFYo/cxE3Mp4jeZ4bCX65acdqLZvbTuC0o9Ph2X
7Fhmqkv/r0fkwWeWMs80dc7Rm5uR0zFiikqB+XKa5ph0v3+UC2IduykJbEa6v+ENM0qUSyD2td5r
WV3hx+eNdo8X3YIt0lyn33rVQQ+r9OrSwDWp3290Zbe8L3DcI462Ym16eq9VWNt0BNqveiB9+yer
w6+9SQnq2kxjdVyIM+ruSDxS9y4KCHDvSd78STJf+aNVfJLS/4w4rAfDnbUf6pBEkyBcRsUa5sXS
PFLG5OU+zR0W5hvXeym5yspvZJ87lNQApNOTAALDn4qAor09EeCOLuaJd/Qtq+uosyGwfru3zRmk
vNkSXw3CSEA43T4y2h61SkF19MYhqDGC497ynucMTfzmr3vlOoU3fELwuLTyWKQafK6uM7j/wxM2
aCU8aYtYXpz7nBZLhOBgqmIofpVJcAbeyHWgiCaRCcbqNgBOGnepeL628LtffbV8c193gvDSPZHh
iJOjeEo57bYPYJGtazLOIyS9KilVorYojWX7QfKA6SpUgsK4v1i8vofCbykywrDMHiIuNqF7sfbx
3mteITeagk/HG+SeqhRhzDZZOfsBn/S1OdFop/svMmMULypHkX2GuFiJ1Buh0hqN1srrjjceZsn9
tiwv7pzEtC/sPTtFfgJouXEe0Yi7/xi3dJylBpjXW+mYGc10uOhlthMcSh0SqxZ21oKacWq2BZsj
3dnjbnoo4RCivsHdxdcfgiyxpoZ33WHgkwswKIG0Krr6TlBmjfpQpr4x2KkCHagvmbQzL8Cw7Vew
Cv2a4N8piThhgLfP11PqCNeLQLKTPHq3EXUMF+LjJVYTNhHFegyti0nM8woseOGOmBVSoepLyrH7
rKqIfGWJEhYGSIUpZZZPqE+v6ULpOLlGzXqxSPZjqJzqFj7+PPiZziZXVLdpg0V8LiWw5OyH8R9t
64eJfg9DSoExX+YX6BK/xM2O6sO3W7KYpDtniZIZwusPJ7NScppdhgDpFK3J8SB78ieiDF/X42TR
BiPmamGVs3mGInqAnX4j8iv+fik4L9oyjKl/oO7CGA/eU8Vna+nBTh/DQgqjXWUIYQYBjac3F1SV
PkrgIisNNwWf4VoAaaC1kYHojJOmi9ZFqjXhDZGyAqbn9eJQXydFUw1I0bwnOpwEm2hOqotEk8ke
Zwb52rMW9xk6lL+hMv2QmE5Whc9alh9ZX45D6BJAD9DkEGR4AYY7sQLSOaiqXwEpBEc/z3YjgxGU
uUc6hlwMsJEQp+UmbWDi9asPSSzNyumHhoFhRE7D9SI6+S4PxtNOeb2IvUqbEAGeMTUflk7Kqljf
bYymqcnAIwwaUDZJt9FoBvVmRCzcczoVjuHtIRlHSjW86Y0CZuq9KPoksfUQ04T7AZRvfA3M98aT
iXVSxDcdWwav9a3it2AneTxmPjD4os3K9v4VLjp1pBRL5Jre9/R4zMKtxTPG3NKgFu7NynodmirW
Lr8b2Ijqu5sG8r2+rZpUG2cO6hZ+uG0j5t2EXHCmbRD/EQAJ1xjJoW3lRU7ZjxMhRdxTkZsIUq0h
IxodlA3nvoz4QdKmbM7N5vvvejrVieVEaksYzSMGJP57sPuqxOoKVzgtTsr3rW4Ljdfc0bcW2LVc
EwVr4JLF+EuAFXWmoktf6elNmd0WW3Ex3SQUUxvete6Hqau3AkVy10WFlK0gPp9Lxo1WKSBD7Zcl
1C65vlPRiaoxCxgfzwO+JSXhAcWOu0t/c+VNOhUBzBxY0b7qscMltK7j6s12p+yC5UwajAx/vXwS
lwToP2Z/i89NY5Wg8xT5syA2oDXQ2NV33qP4bz5m2aPkJ+CUfjracPJ/GJvUk67qUMgarop7XuSU
GWHoMdXxZoh0qgYkhJyegv9ncC3pu1JNUGnwd2YgLR0Ym+4Imu8jeNGlxHnJUNUSoPewactRmh1C
Fnc7IuoewmlplyTFFlYWquwNynncDbka1Zmncd+3oqKHzO+fmYAtQR8j9DGGI24GEs+SNtIGye01
lqB4jS5s/oOEOERxnGn+2G2o3E4EpVqvCH3Cziun+wBB0nuvIDKpFRfNj/em95CjbJs9fxDHDJ2B
FbS+SBWyBi1+aXfrruoz0cBamB5qFAlDrPeYK6mAC7IdD+lWMynFortOsbpl5Sl38eTpHMedSrxO
kRsnoNEEQD7W0r3RgYZFo/X+KUpvvQYe8jFMhCLVM6XLqL4m/+LYRlu/Herd3aF0QGKPPw/zpocu
qy5vA1pxnawnAA17yp+LsWPVdujtvhjKklQgaA3QUXlrdXF9BSELl7ZW72SyakUY2Crsp64xlAiO
Y+z1DmbHxsPIiTP97cuTtXryWRXviBq7Tr8njz8UBD0CgpOK/Rfb1dkUk9VLLtKnh8/8coB8kFQK
LJCgOVzjxRPs9SFU0xbFr2lfp8nZ07mBFu0wLW+LewDnXStVwR0bKCM5uaSCO/jaWZ30l0cdcZM7
dwMMVP9Te/MHtHhvBBvqppCAyu15vlPRbXd36k81Y1EEFwbwy2w+hkQ6JOrBNpLx4i0n1wMc1xYc
VphLOHIePjVuc3LwwiK1e8xTVVsNw+qm04B+szGoiJxumCSd/vARX05EPOqXcrlodnkiDjuQpYjV
lnWIDj2iVwq3RtO4U8VAul/xnWEiIBR4tRMyDqBSIDnAZib7HJj2rmzyUIbbwF7vRj+U7bsJJrzO
UlLZB3u3vJW4GW5ytdJiUM9BEapF9VWGxJbklag2umqHx8Cm/YtYaDIZtpFTQbMfUfQHhZvrj2NT
WeAXlFSjlUY0mHr4e3tYh/y118v185UGgx91To+8vAyFBQI0BufYtkFto/e4hTMX5yZf5cHAUn+X
hqJx9WlL+l1GmgHwR68S753ooY8LoumGjjXaqZ5jIiVrUZAsHc3e1hqgPy9KCeR73wUvWGzcXT/s
LXTk0gCyF7HgvpMtHpjeZdoNPl6bsnBv3F6fnYqnHp24yE+iEXR2fIJWK/Su6UDW03ZkQ3pCUWFT
SNw8LSWXsoZfpown0hxol8tJunOk9JuoidxGN98O0kgNbBVIfmh823zWi3MMi4kQCWdNEvFaumDr
rQVr8hXb1c7rlBGNjtovVQ+d9twVBsKEXREVPHkMqsdH13ywY4fkyOHZX2ZgI45JRpz7QIHpVtLc
8T0Nt28DNM4MLT+YFxzHIK5+chWEPZowrg1QAmT4bglukHjUSUePYRdvURbOuDLEyrvgHEv2H7Es
UBm+wVevnafFzJ+cWag1XBBFs7RCe/CPt6fpd3wO13tGwBRLLCoKVJoYmLa5aTl6nYCXMsnidnZI
GMIpKVfz+WmGmFJXzfYByYuHeyPlViOtOEHCQ2p3p1bYKoi6GDMlw4M8IqIazk77KLdJOF6monbW
uo/Xd7XysQCgWo7brzcUDKqDPyQwSgnOi0XbRfOWb7tQJyLxtBvR/8WkkeHJDlA7x7piTwQOjka4
PknGC5BpBaD5+jsaX0Is1kXRkzZPBUVK6sEK+9RVyjZHhHpmLjqrOP0XfWLwcKXFqgiwVVAkUNUJ
rCVO6rYf5zmvGle1riKq84SlR7ZAn3vsNe4rDuwrGSrCKDd5SB0OC1KpKR9mca3LcD8v/6rvKX7E
RuAdRzPhWUcYeKyJTBVbRAY0sXqDn7vj8v10Rlsom34fzrwmJVhYLuP0QPS9ABRICL8d61j5a5qn
ddGrkSULE7qQH580A9Lz5mkYZ9ZyGFf42qY8JtOrN/PcuMnxe5koxlqv7AF6wTWLV4c7NpRA0pop
Zhb+ueNUfT13hK+PDtNON324duRpkxEyrePCUemLrnvoMQU7yOORPVYq5MTPV7uMV99ZySPGD3Nw
Q9x00wY81nBLk89KE/MZ7JcAbWL1O8+WPZRJNz9crLl4xnkPjrpyO4Jwd94u1AF4tmMcCOn7so4J
gPB8YagUAOGVYvoVMtniyeURs0NIYdH1jMi0ATEuFVunCyrnW1xv1T20/8LsDRpNtaF8CFfip8LH
MYW1eVpiyTF8L6EoP2xagSU8ustniMY9MsSHI/3cyHQNLeGBBYt02zqIARVllCFZOrQYuLZLfSeo
ASjVmm+8viFqIFfNzY5fjv3JpeAED+NqpgGBPuHs8lonq/WX2wCq7GF7yxGC3jim3ULzZA8Xs80w
ik/VEQN9mq973lwq+EX5QolxTQLsXKuO/3MpeBJCa68HUxfxqCz2R6mapspH5FFKf58PUAnmjMlp
uj+t3JPbOhu/C3o3KFHCDDREHkbdZgaHXk7Y0O57LyjJpSmoveY7In4htPfXrkR0mc8hmkri+WXp
i9HI44JjCKL+Fh99AoEAXjGx/J7MJpwO9kNPllZibld0khFxB0+cHyw+RmF0NrOfQ5qSl1+yWrzw
gpRsa77+j4Yvbll91Np/Kq1791vvazz6cCzYovtfgOg76J1JJQnlOi2uzSNeK5TJ0G+KkW8cEYxB
BNC3Ji+LzJgjeNOLwyYIJ+YgQk34zLoNxZp3YubBKYPn6wYLekPUsPcn3eVGJStSGEsq7V2rEDf4
EsaVxy4IQSqY7vEpApAaXFZJMjm6YL2luUq5Fk/uJ3IPZy2Cu+Gz1zF+I5l/R3uPbrHG4+iVKs5K
NtAXVVp80Tw/nXMFJ75e5k3juFVle50t0GueltVX2jTio1sPiz09OfRbA2XlvTiiUtVC+sUnI4qh
CxlrD36WFHqJ9Jqof3Ttu7iGO0CLp/qZ7ZDbzxyfusF7vc9KYmwbfn4PnolP9ScNEV1cXSvJe6+q
bqTyD7ZlqrYsa93t+bWdhA5VKygMEC8BCP91+busKWa7LGa16Xv5u3KwDIzVz2DAqsCu2SykhcPg
AxpZl2aYbg1cVYG/ac7GXmwU/qPRZpC/AAteAcxetjdiun5ne/FHW87qm8WXBDei7W2r1OR/5N9d
wc4vBzRyNeeQbgOjZFp2ib32kMxWddofl3TSpDJtp84YTVWKprn4dFVf8hT00zhf25TuOlgAfpn2
Gc5YewoVxPqiyb47jrXoC/3RQtayieDhFsgkb64ecFWsOF5dHHDMBHSSvAGSNu8fRl/QWxQaoe0v
EGpZ+zwYWrcB5p/nSvi9W4+MUDu8+hNoJMIlVkx+g1uXzEXQi/sWNAfMj0NIFWQkERyGkoozMWrd
aGe5HyxT1moEdnUcSgaFgya0PK6/hyCtdYkAKc1GwMCiW6eW63crE2q71uXWkwkXljiF+T1uAwLk
tKRG0XSrRD267u0fE+mMeDYg69R7Fzw/06adKP75sVw/EgpxuptjGTkomN2cqy9o+hccSfBsxoZu
vZutwl4agigRF8ewCyrK/BtQYy/jlpl/crPud212vqncGZzyVH8rdRUGvLkFXBlc+/4D2lvBUR0m
p8HCb1K1APmJJRhcTMtxM/jGgIVsvPmv1APN+L1PIOyum97hSIjdtSPHI9OUz7FOg9kTkCa5/Eyn
WodSPuSTlj4twRVfIEnwJj/nqfsmQ2q7nBR/02om1fkke6ecpEEptjmsNTqoDTX52ILLBfrqnpCt
wiyCfRamPpfTm1w6ALKVVNrvpsh/KI6SIFbuoR2nTX37jiFliXq6XBqgMOC7HV1bRrsJE6g6vol/
wdvYJvlrdmUjhlLsOq2EylnN/qeNhV1oP5bRpmlKcMpVXgOKugf0LoU0PHpeqADZ7m1x+P6P+XmH
1VPU4f37nWXIDxLXcwbKLFYNUYDL6jVTQQEEDFBUEDrFMi484+XwZvPV/MbpxlPP8B/Crr4FMAl7
OnlPTYXSAJjjvvMn6b4p9HtNteN+CrwVkP16hXk4cJtojXSLy8akhB4oUPE4JWAbeTV/grBx6yyT
nNHD8s/ZVgL7vXFBCSctgdYIRmnFtjgMuBhcqvc8im8n1Kv2TyypsLcJQftfS3MslzfgNFz9MHDJ
6tSco1rwUdckSQl4Lvx+9hnAEbiynLq5jDFn5XgSMWYItU+pvzSQOzgcBuMfDgyhlA+XkQzQqlFN
r1mnGVZqws6JpBErEbHnLaoZRasj9dO7r9+YAB7QUPdtzFgotpX0e+7ExgCCdRE8rKkltYud/STR
3HiXMQ/1ugiPQ4jrfL23LQ0BRdBD3xRgVZGGEStwdz73FhbTW/QSficuw8vMli1J4kwAVe8wyJA5
4EGRlX0LSm1eE6SMmDeePsZfjuFS/GG3/9yB6vnaN0mr/Hxhb4koGXWE6AjjgtYekxWsQFrAoYul
qFT0XMnUk+0pv+yQRGkiyvOyentKXcyuh1wq6kt8dfsMFC5Z8Zvl/CQKn+xGcwEx0dA4zlfcufa1
hH7wDxw0J2EUYB+YLKOlEgNH9GFh4PXQ+o3rCk1aiLC+WvsLQr7xnclSqjyZwuenMaILZqlC9XUd
uda2E+xR0nJQOZLDNbn63bKWy0jkS6/qDXlVzGmQV/XzKY6GDkG1jBDNngF3qcQd0yjttjNOUXsQ
v2qCPcw2vmO+C9lPHl35gm02dvICgc990tXLCtVkALQuThCuQf0gaoF4tSnmH0h5oKnJkS9q8OhA
wnQN8jrHiQUhEtxj1MXfEDZzGS08ztqvfK4LUCs373fgBOrIMuO79iXAfojnr9rAnCSb3s+3ksmF
TKzOlRs/QA+TJ6fMMGFUuLv13XjON604xSdTGYyxKsOhg+jBt7pGXetwVgJe3UYZLVnDutNxDOCR
MNf2Zig1zY5YvpJhR2zYnIdPUTYsihM5gvooi8TSIag1eB8OJDpQcUTWifqeXwaT6RTZhjtmZ1wN
VVH8LHEfgc+PUscC4Cgdif03a7GOtY9xqoQQXApPC/HgU2+iXGJZQ31+zt2irUl30UoNiKePGKIw
A3hZNfSfETYJaN82X37Rgcr4tqwJS3MzuW20xlFPgzUoISIAPlbCem61laUV9XLv/V/d3hJnAfBa
pDxerZ2ig3Yq+shcWDlDcL+MvRc+pU08WklxpeGJFPCy5wCSkxL9FPyW99OpiIgzS3K8EHHm+u/O
sE2532a6Z5dCosG1Lw1gtC5UeeQgWcYJ3W7QHvPDQKIVtzBhJts03F/trl+78/dbKbMAAz1aI+IR
VcPlNJBLMxAfcE7hwWmhOIpyfnkpmHeQkV7rJmYjnz9TVml6m9PppBQ9bNCsgGA/xZOtFVSA88XL
T8gIDJPf61XCXggQRNWs3jc9OGZF0XKcPa+20GLXnjGX4i7ztlEbi4y+I5XMdeNVSmy7Muuca0cz
0X83Hz8TFUuvj30LWTr2WpGbompqVwiz2999Rhl2pKLxHuY+dEHAye5140XFRy9+xKUJF3lsZTZ8
bBUAJuf+PFR+yOa0zsptDmVQ27/LK7Qr9v6F/JWBuT2o8UDKfuBn7/qQj8iCbFkIiqDeg1tS/AJX
YfNX5fRX5oEun2FOzisdZ4qYEfF4qJNQqF1E29s1UI6QuO6my2dUMc2/2ZmM9kawgQ0GT9doJFdd
4Y7V9zCnOsu+V7YlY2M8liOzhhAA//CJ8lvjkoEQ436N+E4Q/QndOtqwRUjvmHt5tS3S1DliXx0s
snFm4ORRkvJerHxMxXaf6nnOU3Mcewkft8W311nNU/eDXUvLS90AL4bXlJmNUgVqit1wJascfwBC
Cbvj1eij9N+ZxJhe7QNtTHsI6SJzedc/oBBvCbluHlrx5XgSDO3otDflA9qn3w28N8Ntc5GsRcHN
Py/nPSh+2rm6LlpxNATC/1hQj4hcthnC/EH3ECF9ncqfyO5YBof0DJfc2IS1YKPZtFX9lNcgwon9
T2qAvbnfGwZA5GO4uf/QX+WkSnpQ7r/nqs6iKeXTL8e8Js1gTzyh7CFup47ge6Do3vqGs8NVlGM4
cZOwGcqGUGmaNTvARdrnYrMZ10z5PeCplMggz+AdVxhkXld3OaO/YXaA2jPjRIdLTZ7JQ1zuAzmN
I6/Y7itU2jcyPPBzpXNbV+8ig0uuPe8WyAJRdHu+m66AmRt8GkPcZabOOEW7k55oHYs0WXt/LT3C
eZUx+3EHfRC5FLzFApdqJhuabCExAfevUbuKyjLFj3wCl0hlpWptVvnvNjnfJ1TkYEcHNvs4RlGX
x1ZA80IJXUeErq6/bI/DmGTjJbDBrmJHP9m46Q1ceVMJqpxKSamBrY/TjbYXfDM8z57c/b1ZOGEk
/n5epdbOzDGbQvb3Z5jteVe08nARBNBMM+NBqYjCwsIuCZfOCargn14bIfE7Sz6Ara7LY261elz5
YfXOLj++KdyV9UAGddyH7Ij2/UCmCAOvh75S0feHXS5M61FhWUnVia+H0yYNvEmnePJ5ACbWXlWM
60RLaB0gztbC4G71mQul0ay+wtspWxhusob0RAXgspXO+ILYVynRcotKMNezWk8IVbw7TGtS3ZKR
EvSMX7Ow4S2cSxCbahNOCwfvUGAkupk8mCwROU6k786c2arOJhxpMzoVGdcxKQLYNyEdbGgX9boJ
cuqszD/dlUbqQjgZCgjlvhfneejSX1dyqKceBLHfbh5tuXWeOmBChjA+RGRbEuqBLYBbYGXNJMYh
9RpmcpGki0R4TkORBezs8m3cfT64YyveluS1T+4MRTFBzPOX5Hd0P7Qof3A5XEpqhtu9rSLTvOsG
eEgVVd4akBrWUuctMtvUsGuBUpgH6rf0ta1spyW+X5KiLDQPQHncigk4DQldHbfknChgrF57iFaG
trxyOve2B2px4WV36ySSoZQ0MBjJXiShI8e6RBE1OHZoU1nowug5iqW9kxmx5iWRa80zMWkB98kW
VWH0KqHFWGHUBDg5WGB5F86KhqhKFNtHjnMAS3/wDDUgcMbaeKf0MN3OtnuT+AxPpnvcqJ+fNUhf
VG92qqJT3vi1Iv0XpfKR3tehEnHE8SMWnQJAP3fPyoR2QafdWwaTONBi5Id5w6toDje3kmYECrOq
u8oTnKwvxXy4QVrp7aJG89TSAU85JXxZzMtF58VNLo91TIIIr1Uprm74aVkzdME4cUxE4lwuZeKf
uLdoEEzDtVoDXg4nSPy2IgbzJyYnEyOcou0uDx9xNxXBCT1QRVO14sFTCA0dobVdDwto7tGitNfs
SGxgW5t5Jb68+7G8tMOFclLfNolGzpvxYdmJdk/6C4xoy75ACuK52H6+i1mmJBbMsVgiUPke8Vne
lemfauJVt/4P2/nH9fvjVEHJQJghr3UEzntYau/VO1OkmPQmQCwa/HnzMqyjzA4AUBefdTBXZkt4
0qbZYB8t4jxHdAPJvCbJivtt4tCxNDjYdD7e04dNVGGMSeXdAPcpeUf86xxNDTUeMJN2MZg5vLOT
dwJHGg429rXNRIhdaExNx0e9/FBokYoVhowSoOLBUtI0ZDvhz0y2m9iT9o6nlpuu6AsgYxl6wj43
EP1bAJjnaxC2V9L63aO3UfV06i1f/O9rN1aYuc2dZOeqyUVjUNTOoxNuSqWDCK+wOPnKp3H0Z7Rg
2brydLoAe/Vx+ULxQy1BlQ3gikO2yv1lPfMPsNjbbZuic0obPZYkvAPzQB/ElPQsL1aRDC2glnpY
RUL5m2RvE1RBBsdgH/DeS1ik9c7l3+ac7gjZcc4O8S6jE/zWFG1s8r66YPLGR99i5F+UviZKivKu
U/Od1CHEBJBtBCdo55UztExL7JcCebXbrwDfDUnUihQz5mqPjwJ3cM+woPwfFip4cyEabuMxSIX6
BUWUd0eK1/IxZr9v711PweCPZpc/Yd3k25x0T+TK4O1CF0apbG36TYhsf3Zy1zCf+4TQzQ1295TW
5HH8P+XnNQFc0RAXWaJwyyxuM+ccsDFCvroWuxa/nnDq91V0GdO44yFGPLtIE5q7VSCSfVphFpnv
1S+CAdsOIC0GgQaI4VQ+0kCkay2RbG4CpqLLnW9td2xvGeHqDi6gRFdarm0rLMoc6ua+LRNqGj2a
OE6zEgNaYnlWDgggqcM5Ddf4c6yxzJpFm7oLsb885VXlmaf7GjZkX0jSXjjTtCUkzfkkDLj2+H2J
pp4MKheTEB/YoQMjkUJxhM2thfGtdXaYgEtDZoIXsKHuorRdbKYJYKrniCMg19PXidS/aaCqbvSV
yNbginiewopZiUE92hrX/wX3FLXrVPsZ/8supCGtCoBpXLHYvAT68Qx3JxacfYomk/seHuZrmyWa
ls+PnUYhxT9jPWjAP2+3qHtrgxDHMU6mAYUBJXdHgLFQjixGPu4LtTpWlESG8j96iA0nAf8nvq76
IryttTiUTdl27YsfVkNfCDVR2FWKnRw3FUKG+DaQEygP6I/KHV2LcEGSqhlvOs163u5L9cnHe5za
BoTjSah5MgVCniAJLI8VYweIGojDstix7WmIhF+U9MLzCJzx7Eihx4sARWgkrRxyYPEWTD7JbRaX
sSP7un+LiufMKSj2P8ILlr9Kf7V01p97Uxsyofx/N7Cy3KTiFoGQeRwN3qIL/Eqqh9nNk2uj1FpB
eiMKdFJFDNeckEKBIlSOXdCP6eHMlkizBBhkfBhDlZf5+Uat4TAB2+lA6SOWzTCpoca13Z7Nv5s2
MAo3cYwKIqO7WuygTmzahsGMBVIODTPKZ3IJGwnr6k/I+txzIQqz8NWfmj+4xod2bKWMKPGvWLcW
jOfquyKEX36pOtScQ6BIbv83JTZiXtlE56pD9Te3v1TjpwLNfTk4Tnj8S16SthiaZ7Tb9FykRc1G
1UNTll6hcTxVzZcj6m42pRtJVGxAKLSS4LpfUo73FZ2faDhQGFvGCHYgbbU+EEi2DwhmnG5RQW2t
dPfT8cfe/uKq125C0kHx/1LVvg5VBu8ydol8oUaYwDmp4JXXhV1mEBGp3Vh3aM0SGz97WYHOq9Lh
blxLfMI1XiXWXABCXJmFEKYxLZ0vwNGyTCUqK6vILTz2sYc7r8ayvO4911PYbaK/GS8oSRkdrqG4
g3OAq3Ifz0opmHl6GJWrb78FN4Wl3Ck6WXSnlsZMqVARUxlVBa5tZGQFBkaqkuvi6en0JIrRBdt/
6A7mLt/HZD+35M6hObaeZGff91D9GyuHIGOmmoCKKHW2AR8qgUWwcHMd4UkMTLaeAVx1tJScvhCd
hec7Jp14k3o0FE97LaThLhHCFBVz7bzWqKYlMZY9MAaBK/cvRrZyUlUz9+eLcPVVhH9WV8hw73KE
LbFDPkxU2eN2gzof48PSxOIC8msMEyXJW1Qq4kmmTAZtZAXXQGgCCW3eN/t+pYIytQB9gn5T+YJ6
HF3G5iFfadIKxC3BbUIm8tyM9q+dZZmvyJDjVnNYaLJGUicWm9irP4o04StRmkLPCmN7Ihy/jqIE
IPaij2RjvoXKSheFe9UlBpUX0Rk+vrS7ksJeBf+7uHieDobS/F8WG+P8qNMxss5loU0sHun8pErB
S18RTcLqv98pXZNz43IebkVjCxcTOW3W6LK6Msvz+Xs+jHwxLxnj5DW353hiYzvD9f17T0VEBfdj
/K7ovwS+CCbpeyDsWt8V3BNHoKgEP9SGR92zXCsinzSMf9kiWqB1jOn6lhORJQendxbEA3OW3FZG
E+uf4OcAdKqqdbp+9TuEdwPp9c4LCtsQqFVhY2M+rnMw2F7ptUT32jy0+d8RNsaz9+jrhxulGwh+
ztYC+rDFO9yuooxvWjtoKqIXoY9YKK61YbyDkY8X+67wS6v2BB6bqRPXDnRhRLFZxit/WR8X7ILl
6iCHVeaYJdBGDGzPiYkOeOmU2z0vIvoERLLf7qkQWPRCx29FzfDkrdUYfPN6hid2sOuJbHVji84G
CEAjjTwb6igsfYbjqxJRW5fteKN9byE86/+Z4Y11MqJUhJBOnlyY/fY15UbOQbaXT2I6B+/TuSjn
3Vola0pcYoBkjWlrUVG29g4SMpn63fhMGlUfzYgbzb3r/GSgJqbUp6Uvu2m9druqonT9WvQOkPIc
c47hrq6Wcsl63zrNJzNc86Lco8uDcwEimnIkcLKKD+ZZw0XUF/GJ8iu6kTNZ2jlX18hRTc7vgSYa
4MJy4JhHdmsZWxcLT7KsJC62DXLoTaRHqkN9fdNVcdEYBtNGrgy+9RCada/EmBREMsLxrtZAr6Lk
EZ9x+h665Ubbwr4o6r2Htw5dhwAVx94lxPsEQJQfUVRWzNt07AzsOulAIvfPyPqYoQmEQMAQFN9c
7ALKIWWSnMWLr5kDkayHI3V6j+binU9+TwoSlGuRmza2nQxcro8GVXz09/xFigy/Ko2Oq+z+BxOB
H3xkIMv6MtB+5d5mAGV7qaZQHs2I4dfdUILjgQMjoVxij2Kb4ecuy4JJa/jaUGWl3YWKDmSQ/mXm
Vz+BQ6ADqtivVjAUDvht2MdRNSdBdKGOOSZnKeGeSm8h3MLklDQSBSgXaPcNzH2Vvl1UO3Q+YUAV
ghPYekl9BT7OOE7FShkMeRk8OLlS13ilWvOgoi3d4P4J+Qj8rWHm+dMAoOUPx/pHn3Mwt9rQl//c
GcOrVOLe4A4OR+24n2Bs2UqoetHIw0HWajIOeKO5+y7R6oktFlri/QWlZIKpH1j1b5yEEHxvOWMl
7Ty2vre/t4EeVEzD7/aCfXflX7ZqD3SvfX+jJ8zf19r0SRb7gJP4tEoQUFxj2ZNMpSK407x73o//
TxIEEy2Ere9yV6gupDLPY2TxNY10irCrXl+RaNqGzLbhqKM8F3Yre4Y998/9cxqdZjVhGrmm5nxs
DyDOpKpLamQmhGagYLvZj+6C6WcBAaZqETKHZnBTBmeLbNqPhTUcCSSCCwFC8cyRQ9u3m4KJ6IVc
58FbS8WJTemQ+OwOYA31N76J9CHJGlfUdP4k07nGR8ceCn82VNdviXJN5ZLbzsfJJLoPMOTWaSYE
jni+T/epSOAgMT/vvVkN/XbpCJoBL2X/RFXcDQmWYg9trwb+M9gx0gR+d/ogMY5KkWV2DcEaohiO
cthJz341ixdV/m5lbmRUWpF5n793e6+gGRTFqelVYVVJ854y3j3NJ77nc9wVxyj8mDwFCVNogy0w
1wSGCsEOvKm96BEyJ5dkhRoOqCLzcoDEApHoOASppszs0A0sJCC20eYfaDLNddevvUkszREnnLo7
9zUTn9xLB67bAFfcFvRV7gVp+DrKe375ciqZUsyBef4c9T41uDowUFEXwTwqixXqwzAFqbHECg2v
XufpkdQkpY7PAIgbRxopjKHVHXcrYk8JbzNBlr0ib7R57qXmXlulVN0jO4ggshmxcGS/2yettQ/b
MDkRU+Z1IqXO42CX9ZJm1E4SM3ickrB4WWDQ+b0Y7gfBcVZuZCjhH5Tu4qDrXwOjWdXV+9eK5sc0
l42dhZ3SwbQAomWAUd9j7ExTmcbQjozNPbzzpuw+yLiD+ZIOjOr2/nx2myznZSN6Xl26sUMQmTcu
nSL7AQpERFb/d6KQKRnnYd/Nr8M4NAE3TK5Jy2eqN3Rm8uopFE8KHStv0yvCyt3YoSNMhbyHdqp1
hsXgjEKV7/imUwk2EDHgUY5NBYjE0deIa5j1ODjuyAX2nkcBBKiITxePAAUbT/rvgwL2D2BTM3vi
GvGgDy2Ys7lPbORKZy8hcKyPmWYq4h/RoE/U9drEbCssGKz9b5TkZ7QCIztq2R3qY7rz9dRjQZtC
2WmcL1U/xRgQKW+Q/O6zv48ARrSFcGKBZvKfbKugawkBsAW+lujfgSdb9cRBSJs4LB+7vpLwACVl
DUHF6JR71DyCqmFIPCu+EL3mm8YaeZSAuWNgcbkxVADjiPWAA9ZH0hG2LsrYRIqanqTBanrUSTB5
Mland9jvYQ2pWu8zsB4TKXT74mV/5jeNmVhS8ARuvleceBEHCbCtZifxYiSW5kJbZnmb6/6aExvS
vTzTSQVcnrXwH4lvul+IfMm1rFMN8tHclYGWX/v8EEBOat7GbpwGUQ2aFm/y9ANrwlNCvRXr2WCt
qdypfrNeGBMS10Juus/DZXl8PBczRRtW4CkYrjCLPxl/GKX3apwa8PJ77ZDI1kl+sYZBZ9TBS1et
gzC1CEonRuz6eLaGB8l8xk4fBlUEA6YRRf2nNKDo7UpDymlm0Su0li4LeA0gCkUYieOtKGgnmvbd
7+KsTt0c7zrXw5K5KN69bCVc6SeE7dfmRyAd+Is908ucJ4LFDPiJE89X7E9rBZcB9GWkEoCjq0pF
alxRqHIPykkD8v0QoVzr9iL4ELuGCa1UG+KbgHiDWMP3FXY3KoVUOXIQ4P/PS5hEsi0VQ6+UGC5t
by6OtZYanEFgaBD9hjiEmXeQiBBUVeQe7N1D107YqwJfk0wNZhiVOY5JKEW3iDU2y6EWDmpYcxsz
CGDfBnnLL9ZrYzNIaGwU0YB4dWxGzhqF2NzwwDlith7XJmCFK5KMNJaCugf1jtj1JsjJbBhvxasn
VCp5jA1UaJMaLxHJtFnf1ekEx07x8JkbQdbEKEj4kh0R4xF3dheNNKhgy/+EcBqeJZcPSShDcX2V
/X6vIDCPloiE40FvIsgOh/Vlw4vittVkJcMND+D2Zy+A1hW0gn5IdTeNf70Ojms233euWBWKynF2
0UUNqnMB9nTqnPfTbe2rS9qKj8lxe++hc7yBPQh7R+MDUfXfTJ1owZvrrHZE68nszrTTX9qqLX4Z
2s0M788Btoxod1Evx1xIlUID/yaxPHEEuvt3B4KUX98IoYKV2jCjVEPyNa9KgIQbFkS2/RvB5JYc
IVu2gPEMZrJBAaNqtMfiLu2l1qEZa+3Q3E+frm4Di1C7yLgJvgDzxWRa5b8iCrfRqx1RdQ+1keX1
gnXVFtY92q2cgDdjnN3vG7y4bH2i4rFMyVxqqxJZJHVA0Qh9fDNmyoCw/IfezQx9qb+N044bNA4Z
AybRgF9ULbvqeBkKhX6YblIv3x6lrHNyEbJk/mFi/zlN48pxqUIz9HmBqOX+G51MBwwxjOaoinjx
FVgq30bNz+zazPn99X+pm8LlxFCbUrTQb73c3M9TwVeJ6vulawVraNHbkInM4PQMxsW/gh0qoWxH
WtRUVPB973I1sSdkg8kzM9t7S7HU6WEGll2KAcF/asZRpLlqEl63wBvX9Qm6dxbzGfENvjmuZrvQ
LuhJ/5xyqijvOC6HRDwhDUnx0bAUPsA0OwA3y+2k8noqwwdu/Ov1nPBrIipBlAVBsgpOk0tUzOio
wwRXGj5Zddi/Kt7JZ1gzaJN41+3ndMvaj2GEQRAkazFZ0LYWVxeZVcdpb8f3Z1tKESY/N8DecwFv
NefDZWoanta/OumSBKEYUYIEzZzts7kz+eyatlAf9Go1Nquu468jDpiqqkK4iMCx/SlDmWdve3vP
nn1alWodqDW1w2uRJLwVFHmZyA/oQf1nA6lYJCp/mFr0CO4FHsNEqtyJpCGuBECUJBoOBhgURCK/
tcRQ0ErE1RoQELy9PtkdnEL/muJIt1S0bReqEkKlKqrc5FaNYgDS/1YUVjOGLRtLvq5dZioyBxPU
nxg1Bn3AsMANEkLl+2OnhVyt0k4vFhZSyys1JDBha3a8CReKhUGTekK3DGCOXk/D0nnPr3PEaXH1
Y9JrD8NSMfBAOxwibhceTn0219eCOcvshxrOMaQUpMefV3Qr3tYc+CFG88/LJ/LIhs38WGC8tLZY
zJ1ogsi1ExtXim96uJ96AA5OptymXG1zTGE5v6u09iOJsfM7VrgsYB4i9mtWm3K30zYjWHJ4Ip0t
xvS6cF9s3QBNPuBCcjxdE0irVrIDrKvPbR37n7hRXlaLleaMRVQqR+Kzsg/7j2OQ7zOWCBbS6xhB
3LhzBdc6Rpo39SkWcRyeUbFPvkWXj2z/2mRTHjV4OpXuIlpqVCvGKOO3Pm6vtkuqA8iTromMUQuN
undV9N9Mjev/QRJu/kZjxSzzz9FGsZrkHGr4qf10ada09ITYLwkeV3QkG0EEex8INrhBwVPQQq5o
IPabKbIipVJySvYbnoLEEJ/BpyKoLh+JNzj1NH9j7XGGh86AN4XBM8kFqjm1wxV58vi1hK58qp1e
xClHcfvRiEQKb/L1qFxRtBny4chEabBY1OKF6FlAFUT9qAw+LdEpOe5L2MfDJEdg4uP2Cb4le/gV
dxzpWDLsSyx6uojQ1hYYRnUhv4lnTSltIi9pTbJe7sXSJ+Rpqhc0rFqNNi8XAEyAzUO/dC+Gyq+h
F7Nevps/yyyJmjusCFYaot6OeSUWVIDSrC+ymoKxxAw27WKIHoci2NUvqNVV2jXl1Ugh9sAqDRj6
ZKxpeL6PikuvFw4SzcC6agmUKuXyLvjTUYfK76fpLh3yNxMq7Hr8+X0troS2licvxDVUUPuhT8Xz
rZuOOUwvBDdsYzJ4bnAvo6HXYL9zCdZxzJVMiKKboEOP2b+iATRWTDbLpv76RC6NlBvOHkZGUZ2f
U/hZOAK2lNTRxUMXwVBB5FgwrRQ33ZThom0bCZDL/Bkio+L+EAgsKLBphmPaV+10HUsH2A5ushV7
emufCJpBP9Qtu942PWJk8n/a0hiwqyIRFs02GBBQvymUj86Hhl18mjD0QP951z7+QsAvV0RPT0h5
+QKo1QTMJZtw2legsjOyu73RvQ6Z4C6GvSQBZ2/lwg4zOmig8jje5dcMZGbLsfjv30QtWCoXDxhe
PZtnr8Pr8AdxMdKwyUOucDhnK/qQWdkfXvXxB8J2r1w3Z5kNUcC64WVFptfH1oM2/nTlgJdfAeJC
ApKsCwhgNwlt1n5KbRD9UetOw+oXgdmvq7yx9YqU9Y7gtxt20rv/1hnHah26/9BicbHU6pHf/Js7
HtQvfVm5XLiF0KXQ5Wy4DFNqklHrs+cF4oAZ+oQEhv921dgvMUJOkovcw0KR6Zb7NaEMpFIlWl5b
rvxRvXkKI+xyt1yvqPD7+4AIsToYXWN3AjQ6AMH8aOJrprIbOqGukbDKX3qkxpOP60wEZzRha51o
Bmy4cRp5AbOr6W0t5Bkyp4DmhpPWMoz6faD+wvQBfUy+qtorA6GdBgtsQbiZrJWwdrAyXDk8+1By
kxjDmncqCz8ZnddRkvlzBnuJFfvG/ZJHAVwFwomt9m++VDImUu+HS54p1tNhaxblLLMPrfjfiKOw
5ptBxW+Uv+hM783KYxUT34XLFG/ARSW2e/MrbvM9sdrycyw2gBaGWZBbfJwdc3Yp7aFgGSZuOOHR
HxBZoZjsZQHoaRKbVd0Bbts6SASW4oGohohaM7TJvODjYeS9RAE158i8qlEDzOoGa9AcV6OqSRxx
pIRzS2+HhrIDkLxR/lldYmAqLZYC8hkNvBWj/aUr/Hzv6fumTIRfMarK74/j+QxI0cgRwFNLGuxA
Wti90T60DLuUjGa/FigIPB0Q76BnFrteXk54/ff8qkLDYR1iKcrUf23PeYzFj5E8nmQ2PshW4WQ9
jXoHRtmy8ptHKVJSU7ITcUl1qMedlmE7suFkKanlBJ65pFlyY0jShxaXRFMq6aHaitbb14ovfusJ
IwQjyERx5Smods0UQ2HKyNO++PYLjD8xlV9FqR19+p9TDm6T+z8xxOxD2eEfrlTXlNjBpFCFusQ8
WZz7JlIEDSOcPBzizRZ/9wNsATjV4Jb0Qq4J4LkWd2QvoVtiniilZoml6/fIl2IeUdzqxoc8k0nW
aR55QEEX28reX7NoMZTn/IF3E4q8KWswbeLV2RWuRsiSQklJgDNR+vUV2JcpaDq1izI0VwL3SiwR
9uJvZUTXou+1kPXTjtsU+BVwEIGqdrJ26kEnutmM/LAmAMkgcMd+BX6Wv4xnh+YVa0jOBpddhhZd
trvwTLa8+MOqTpyDeDMRwPIo1LsRiNO63wju6Jci4CA/HeRUNcMODkgPTWKKmaoq3BpV/OBWXsrn
B1SJuAXL4oYGyEuFtflV4ZJTfKcDH+dQFQ67/Fl5uU2y8mS7dUByvBQI1mUmnJaD5sAeavyvlnFo
ffEhUFortg16hcA7fSuXkLYxp3YqsymWHiLZzlGHOaZpj9YtLj5I7zRFw4mnke5gQDuw1JLAnS+W
orSLeKUBx+tUf8jCcnMwFrIZ8jD1qVRUxNvXNpzwb38zS5BmR5q5nFPZfMEFyRHkVoyTKv12neCd
nCdKuCO/GbFICFslcX2I4YciyDjGnY60x6HhE0mF2r+SiG5J0M+LQQzIHpnWf1R5dyPIe3GwfzO8
en5SDMIcoE9tLYTlOj4Z0Oyiw5/kOqbWxtAYzYnm9u/4Bq7w3lGaU0Kf3iGnv7Z/1LrX3gHrm2oV
3frAc2d+Zr5JK9XjaPbF5s6C6Zn/BbBgG3oyS5Um+be6ZGcyKTh1N/QcZAFPftxKPWVxFaXU+Bnn
vEVI+QJ9NQf9sudxdkEUhFmGXFuOr72RJAdcFTCM5rngyzZ1IiWu6DeFBeUVT2ukcXvh19KUD/OZ
sws1oCIfJbTrISO545FYGlCsjxOB2KCAWOzjtRMBKIt9RKb6LOEmxeOMR62gApDyLll+J1Oi37AB
6GVwQ3Eld7Go6bdDpDut9o6cI8+EGcDsKjd4Ye67JqkLjY0SsxHFgoJ8ZgMwC0uNmcWqaDl84LiO
njDP/0M/qdFfkBUra0ER+po/Z0cfRtmWtEXtdVvghcY0Zt4B4KQg5DmcmajuCk4cIw9Td4xZbWcr
8/dhryGJG0IYL2qEBw2meVKIyhx4COK0G7D3Ag9TNsAdRIuonSwbigX8ZLoCX9KeisI2Q+ZopjPU
loIRKMKtWX1+ExX2Ll6kktN2G9kOl4jFQOB5Hv+RFM2JiymNDU9kbFMpujwl1zsiM3cI8XAzUAIY
B5ZLe3a6mV3x1OSjqSe32ntdk0U5ilgaqY4qVNoTY0WZhTKgYmM4qKdfkhq9BxgdeEuohXGA7DWY
ILteHQBwj+R1YxAriHnOl1OjpcRInEqKqSD7wzYwGY4O+9mp4gnZmgIQCpUZ2vw3cEVm8e5lezry
bPl4PBlWl5S22rQ8T1C1yLN5/ICzENs32ApfoVaU7HYMDUS7dBqoUabwZ8bL+S8Mx+9jN9WluhsE
Xdx6cBbUzO6e6o9cbXIrFdT3CLabb1pMVNhh3ZPouqlwcAVyeiuydajwWPoY+Wwdy0DlfHUDj/L4
66bCgVDWXLILU0Xe4OXR6zexT0jGdvJZHMolaaTSeUO6UAgN4hipl6D6recspdM0PKhS05saLT4v
KJqtgQPV95zS07n6EkYCHBy4ZhH5inFoOGCCkPZQc6434a8u9FKwEEBwt2vCRXmdn58AiDxf0ey6
arvp0CVHif30BPdgtWHzkLYelaGjGbDSDq7/pRwElCpYtJUKsq2d08qJxV66MDTIEyacU+Aemsg/
VZ5baC0PoG8WwE8PQTo9t1kONfLA+p/+o17MteMbqOuTte9w5GoAJ8fiTLxj1YWQyE64t2oFyjzz
WGkL/ux9WkpjaBwswjd6UhbmAXnMgQHcN6VZZ7qvRVS33tJUHG091gR30s0h+bDqGiVUZDepvHxa
cSKRpJfyf/fExU3eDYySBtAeTTi4KmorJloYtg3MlZ5ljls5R4sXnXrweO6g9FOywTZYUtpL4byz
KpDaG1dd4x1dUUPUlt0iPnZnX8aoDiPotGwz1hUmIdg3ag7l1pDlvY/QGAZuA0r5PDrA4CJb/1P7
0+WQbm7TVaIt+wNNFWN+59KdY/PcAQcHwKQ0+EEy82RPt9XCxWitW+BoL1L4vVDSPSqkGLrXWDmq
s0roRynVb5gjszWE+fMb6eC9p7bEYE+bKSoLOWgCr6hvCtMjAxsw1o5oYPt+MEptnkOHQo5yUMJe
7X+5BTJtSO9OYEErLOctRwamv8dDLHg/tFb/SWRqO6dwQ1u+3frK85D4KVGVCDCot7M6hNw8yCjz
vBmZvQNAzniENWZEj+YqHGKySMh6W/0imPcA90w1f1kZ/KaVslb0ZLMUSc0JVPHyRK7UnQYuRfbh
5RqSe8CldQIjeY0Hgx698ysA9a1OvtRL1sXDGOSPqV9yOdPHG6mMse8eoueaCnjyv65H8x8kAkAA
XqYbRakrPxyEAL5+AgakmLUoxjgJUU6+hFGgev0sgBSWi96HoXXI+3DQ/eTpOfOaeSfdBefzZUv1
uEC8GV/yQoW1IfrdcRiGpD20rDQGooOknhTRiAe9sPxrKhh29Bb7PlgHBldGKKygDs7rMvhuaFf8
eXBLyniPXNgqxzDGx2d+2xOecJPOMK9kVE5DdtPu7+SsJmc77OboPCxwRqEVTjHwrfHmSHF5M/7t
uymSsEAsACEJR7lOs2O5peW1b8B582Njo3Zd5JbbRZkHPqhLhX4lJ++EecnhyfiveguST1GAxDbn
wuVOv84z32f1WBH9kf+MYHdPqQlJjCVN+GddMJG74NrvvUgrGF+mG8QH1dn6+eM9ZWcVGEj3U1As
nq3DeLXUFq0PNm1DmSSFazbD+hVYk3/djXH47DzN83oxagqvdOkL6CBmONl70sqioM2e4ho47vAc
Q0mHDSanbPmmQHQ0CIr0BUGj6GzMODL9Z0+NI2ZwTQ2+mGixFP3tB8VVuPuc4jwFt8uZD7tWh+E1
XFhbi86men8YNgdTDF1DIYvUYwBCkkWQAylYMiZOQMAT24H+ikb/xP+LmZiZ4LavfmqpkTwwxhFE
zX63LPAdG2NQl8NqZsvHQcZzpP0Dy0JOwPQSrn42GzpiIKAV9eRVNsdKAiYRAcb2BA8J68FdAlvw
AmVyue1YUrEkrcLY0RujiyNPfkmdMgTYOSWzgIPHK8upBpP+7IzxT7jX/68RE3nRYXi2tg5+/Knz
0YQq+3/hcvUGL59U1Kec+m8/qeUsMFjiNu+S7lch19tEPRdgeOwyMYmFuySTSxj4QY++udpo8umf
2acg8mQfMLSeAYYiEx9ZmEfNGwAdonKDpnQLNlxNaUjxFTHsp2kppouLGoI1D2TmFc3zj72b4vRj
+bn99tfwfs3GBwQ0fVw590vKxuvFboJrlsrguLxE8uXkQJfiEEdU5CZQzrU+Z/gkk/0mJQB9pC15
hPMLA65r/ZXmy3/rmxcKBq1hfwLf5JWk1VsxHNWiudIAW0MIddsoPOkXQ5ihiuCblI+V69M4g+OY
9WyaOX3idkJYWnGKou1NACEfs6sdaOSw2CNk3OfOiLmQ+dX8mdjoLE28jBr87PGKW4JsewUlCalS
HAV16jbdl0t+rtPfSr7OiJJwBUyWDegA0Z0QQKRUd1eHwG8bZ9MPGe9PWYPW+XMPIEDZtpVfhfWg
XV3eb7sKZaUnE+g3Tlnb5qJdVr0jSAUt0aRuqWG+1134IZ+JY67vsKRM3WBSumWcEql5nBraFmpf
WTLWj51wxnk9iHRAqbixBwvNH8qiVmbr5shT5A/YmyJvqC502UhcakfT9GAz86z4hT6u08gjlZO2
LPM7f/ow77yeiGykPRdF6Cn8XdXrzxZ5+lr5RlFEMMbGwDZaoeJCTBv5mFJ3CncxZdqbH34YNysI
UjkCF4wKA7pzy9rLaE7z4qzwgbFV67ZXiNM3P/xgnV/J+nM53c2bDgmNSxdoxwyRFOtHDMe0YkgJ
o3MLkFpNhduAq01bJVhKTU1TM+jo8E1CQDcXmwk2ZtlbGeh2WJ6ADIPDbyLQaTWzpqaXxS9r1xyb
QrArwG/9ulch8C95DCDLCBCsGen2xBfF+m0FQhdgJPFY4MNveQO3k+tH+WOHUY8ohq1LLg73hbo6
5GYVlgyDSXIh3yqGZHQw09bXp9XWfUh1Nc/HASnbl/KBOwM9lqLRyEgjRcoOg7Agyls8ZQGU6dti
lWBKhLRICXs/H9LQWb0Yub3SNTlcEl14dwbEYtTKElgIaPDmPUccGayC+6Vl5GgnR7ptpVLPqxm8
mgGKn93w31pMYXu0xN0ia8u4xr3tIkxkMDQ1qTl9IdgDvC2THLSJ3+ywkyFvrkw9R1npUmO06h/+
tWb9bIItSLbwnrHsx4bCogvpJVuNzopyIaHWJl5cqWtkybFrwXTODtmQaO/Xyz/XwJnY7jC2MR1d
ZL09K1jHHB/D/67LH+fe1flIiPFXfNgCmhwmPvhXhCPqCyophxpFJ26Rdk0Kijr/7nqhhHOF8+bV
X0clSia91W8T95oaBUEFmHTcvuxOAgBuv2s1U/Tnhl9aoK+swXsmblDeTi4Io7NnvDGrE887YgnL
rXdN2kNGwIhGqhw+jtDcUpe7ace45juQPAvATKZiXUqwFPRNIeD5SSf4PCuQhDx2bJSGty62aHFg
NW6pUeZYW+ErAARPlNh3rsZvx6onDbwTcp3Ssb6KKqzIZ5kyAZffE4HlhpQ12rTdsbyc/meaXOtO
reEfnxgcmhhxHQQ+huLIB1xcdTEIvk7pyU60QPTYQm+7UdoVD9JysuJNHd86NRFReKg8Vl3797lX
5P23A5RFZ5mqJv2F9ELebCURPgP/2krkQgZ+WDChFCPdXxF5s0TRMepKgToWeu83sxmSY9l+cQvH
SKc43isIkgK+3JS/OzFfVsMOqV2NvsgQ5Ty+O0TktoakQwjThzfrhuA4d0a/VqswXwKnhG1QttxE
lugJ6CRmprM5H3a4yX9QAKIOydh8ZemzWYyMd9Et4dqN1tZPYIw/bV3/Kml2JPWO4z1LBipd6Zvh
rrqKTb9gJVLTIyfZk46uQGNMiZYI+mB8ji806KlI6tNgqBx5GKNWlv0sAkS9gmywoXtT8GnWNenh
xh8HkEoviAZtrqeIBpXpIvAscPssICjc3yewa9SruQgtPkjM1L7bjKV01SPnyz3pXIuHYKzHVtCW
eaI8atZXwaM6GKgohD4Xjcqo6lPPHW2DHyBPWzMigJKRJ1PJQc8AccZffhAJccxnx7lQULEQZrlG
1L8hpEhxipnOyx22yg2s+LBFm21dDnvBSYRMG9518uFcUaoNFbxrVyO7Kx7aqalonOyaCHC2wvvg
e28eIh8f5RZkPTSDLgYehjnv5nTJnqrXo3pnqinWKnOxK5MJB6+ohkgLsHC220mt0gYYBB53lWu/
Zhqq6fKF/VzayTFlPcOYHmhH5q+mp+Jw4uMev95WxRyOT8HTJKrQYKr381eUBHMyZzNlhWM0uNqf
M8Ss+OOYotE8PsFcMfOlTjWLOxZABwj6pUAfSWL9qodANuwscZ1vUE5zJ/EwylP0BsbuH5ZY9CTm
5EA+O34zPMcSop0u3C8fkL+JTEsP7abJlw5WwuHPA3VJqHaC/oNIIsVoi+zmI/wyhKUEitpFurTL
HN9Iu5eqJ897au6+sMbdX44l+mkplxDGD/I6pJLd0buliSImZ6zf+gW44GMRrGP+4rLQfWC7+tXK
a+5cscmvuaLRKAWI1DyaFnaYDkqN274I2p108ynWNPLouyw+qFXqAlBD09Cc16gjmavB4w4tNs2H
FV5PeP3vu40h+Oaol+z1HEJD6/T+jqTWEUBN3O7YCqa0Q7wzhzUZ+YRA6RRmoJjgWSKL3vzJOZsL
uyz3u4IUNYKk12LSwAvQ94ydKYkMySjkkDhfANwwoomqBuQ8rV4CXrJrJ6v7k2roCYOpxaeD+V05
KdxTuJtql2cY2FtUBDcmrYa+c7I1A7fC8JweEOrIODl02NM+l6nBYbW69tGIBDdjGIR0SbAGTpmx
jcV6GP79cFnjB92+MJPwvQ5BaCwKVoHE6a+YkQnCFWu/6Z63W8c6LA4wZcP3Gc6nBIpMmveUjamx
h76xWupQwWJGQelKB9DmCp+JI7PsFqtWvnquhNVj90C459fXSubKLrWTFZvGqdVTtXUe6DkykmVE
qR5gkzrkhOdEZQ40RCAiE1pJVNBLhHQzWkhUDNdorVgoNChUxl5wXlXV5hfZDmEJZGCHLje5IXy+
FKprdsnqo3PrXi0c/0HHrAQ0FZIf58gn81nEptqNEUr53KnazEmkRJXvVjhEChp8/v8i+bQZnbqz
waz6eZ4oBeDdPRbxZeA5BL0U8dHTn38EVWde0IWVS6EoXnXA770o8mdhLJ7uGPayDqdE2FJjixn4
kOJUJyCniDOOUj5SM9FKktqYVvD10+qrrRBPnSrTOIVNgAzI988ZD2XOZ35vc0Pp/jJ/AuQoxiRK
qA+7m+SuQk1V3sEq8NFFye2N9SZoqjHPBDWGqLl2njZbayTtalD/jiXjl4eZD6sSIBB22NmHLSWP
fn/OGm37ozSE9NxuH+y0FutiJwfgiI0tmgrSDfb+DDrWPSTyPHRBXlni/JadnKjOsEt7k3pEaPFx
mwAkU10khEab1TCNawGQBR01ZmXfPO20pFaljHB3yH4o8Jon0UfN3WNfKJzBQLk9Yv6w8mZJ87eb
IOU9tI34WVd0sF5XShmAFX7/4s/6N7B655ZnN2KoP6SNVDEV7HnjzC16QGWxbuQ841ZcLttMtdN0
17Vl2xjWHEEicbaPReVPdOtrjVP0pi4I7soGjKXzjQHyk5jjSUvEwao8gTJPihrg7hiIECvwWqDl
+4wyabKfXLNYrZh6ZZoSgMaAgrV9o7dzLJmnrlGnvua6L4+vDVqWFIbXN6W/0zJhS1xj1+KBBt0u
X3OyACieqAARE+taWjbRAMvHMxeubmYHn6Bs5u1UiOOR5h66JMSKiLZoGXQ8bgPYZeZAA+P9j4DP
9jin1DY7pxtNCrtmzKnBVCa/CSy0HoCowmC+DzBla3N0zfDxDt5vswnjxRgZocdGKVQt7GvkPtbd
8obKSDBNzT2M6s8n7okpZYgbo/8UhVRPVBCytTswM7kctORldlBD8udpXUqlHi9vNUuZU4Z64xDG
sJVQWtt7zwTBv7sZdbhg9qIkpowhbFGk6VAaPYuInyATXE4eD+JHJHnP3Yhc55MbcCY84I6fmFh2
tx805ML1waqFn+yRBWUcQ5sBgHoeYhg8N65l5ND6BELwWDJv9vgPGjtRNnl2HamntVctz2HMjyfc
1v+xzwli7Sxto5BU5/1M0WrNYX7LWioBCJz/pz8qGMnJUsg1LpyQsZ+nmA+/Okgs2WPF8JjPGXdg
lpV+T1uBL/6eMKpQcywyqp+10+/Z9XE0ue5FpGB64SAjsvTtN7NLhZXD8BpQUcdgoLkuR437rVA4
7hO/GYUbf6GeW59RVH83BmgiXDJ8ldvHdoB2dqbNZfljReVLaPQ/iqMidE2yWGcTHiyq9jPvX1fT
DlL2IjH+MVDc4u+YxYtSfkz8EEqQo8TRVq63ifcAPkWXbEqYp7GS4yhs9Ap+UOe0j1Yg3tqJRFn8
CO9O49teoWXiAQVIrADnqGzLqH/IdWtQXcEo2oNulocuIbr8yUriQcuyu0rKLGPeizf5TRrG0anF
e2bn9NGIY6aJr8EmWaoDun5Y6ZDzRogPoyVk1Ge1jXBh5eTzvD5PdXKbbutUQvQm25eojNpQHHG+
Te4KzEuE/YUYiq0Tdwkm+iLgowmXEemSNsJ+ZtCx6XtXlPKtkXNHEId9Rcygh0QYk7zntGZyX6zJ
3/fDXvlxCvPRjCxHQZaRQK59fS0nNHpjbgPx6LTfUxUuGOQon5KOumvVgzfSM+jBhB5XBEitWVIn
ofCX82I6EHS+yXHHWi4gc+7PMqOD6Dy7MJVH0iflPXDu5Kx1k9vOYre4VU0J+GOiQUfRv3O7+HEK
BZQwkP916fo1mU1XOMiSOcilE/KEGj+F54L3qDEIdJq4N2fYweuhn2FERJzMjMJK+c5Wc3GWeALB
QVq4r1Pt1GLUCb5kuRCozcln6V+D9ib3Jjniv5obkS/zoXHJlOADkwl83YCpVCQ2e+lR4c0A0WzP
eOK6tcDpzlxvWkaLOXh2LKbCa+FMym/klTRUwbLqtmGQ0D4oj8x58A+JzDYZy1ymeiQtDwelWMHf
IVHmtRVzjst3p/eHRgjI/uRE4b8F3j9FRgnjMfuHrlRDx1OsM5mXkxEP8Q9KBIzbFRuMz2CpjwF1
IoCh1h+ITTHoi4BxBLXlJ5NblecDaFl3QMxm8j36amRpCdEI9e0ToiNZUbyxYB6s29ZBDna2u6Kx
O13kLd51+FL5wSUZJbRvwZg5aFdbXkvRAXn9DpdZA9ts1eMm/xL6k0KHeaPUOJDpxqGfV70a/1e+
BbfkSuzRtJ5h/GSXn6oh8M2pHi6AymPaOMpF0OThIgWih35MzxmxNiux1725KPMSgoNtOECqzlSr
Zg4Q9gZZD4C+oSq6G6E7+2RGs++PD+E5UU+INvPb5VANsul7E8u3OlGSRNku5ZW6p13QbTEmxptM
hNEStS5oEzn73YpABgWYd2/pedQq5yyWa59bv2OCOy0uPaoDWhNzgd+lPCeULbMUqQhYAPXAXxk+
C2TQEhmDeWOa/JqerQk/ElQh1h+EO+YoFDQurTmLYLBlYw5VnQJFRGg0f7lKMU6qudfZl3+tMYRG
9J6d5JADy5V9RKSi1eA0QEh6/Zq4susC/dnFZT7CxMyrPmRChpm9oeIepyAc0bCs2ZKVUpqqWa5O
YRwRkr510kFVCMbtll9p7gueSjOlB5E+GOUVJ6S16DuFYJW1nZI3kWX8rClazTu4ptwzpAuomVYH
N9DZungNcCBN1/cQIjrQ+PK1qkKxaVzBvTUz6/s7/as8qqtvovlhBsRemJ1/j1JXGItx+g/uEEtq
fuPRMZdUckdwKokqrH7GMFV0T1lEwQiedm+b9c8sGZgmUaxPWhSBKcPhIrJ3BScRB3GN+7NuQQGE
wLz5wT/rhhyGiJH+Tg5Pg3tV3liDJkGVcEgjXk6nyuELMlrNw3pOP7VCSINnGSSkiiq4IQ47uUCv
eCSeqsUHhFaqS7IGKs+Nvq0Wr6sHaCkgR6/xdmYXqEPa7+64LCRu+rnjbr2AilHARwIrwQHsY9dl
GLG8JJb4r9LIFcvZnD0943NbbdK2Nr8XdkIy+eXppDXnzgKqKBd505MazCTjWZm4eDLJNiSf8KZl
TzNbZLaC9fK8lhPv8QvPddtIZQFXFlxV08iRp2BsVdjODOerUMcw/bQ4tiYVEz7UASVDG0987Wnm
1ICxRc6NW+wGUkc2xDDPHw5UMFv4HEGypkcIRA+pBoc6W8ik+680xGomfF7iYL5pcDHMTP1yfi1G
k3D1sW86c6iaKWxqs5HLMnab8p93mLMbFtZm7qSUtyMiojvOjoKkb/qzMZkRNJAYhbWlrJtD7U8d
u328r6QEODoj56YRs/vLRXP8DDBe33kH+ZcBsRJqeLct3sdKMXHGL5nsI6olD37ZTU47vdO5vihD
cFd3euAOIG6flzQguR+XywemfM3bWgjgpOpVJFYD2cEPvY7RXM8zqSrNOuvXAziC2rVXNIdto6pj
e+ZgugB5mdOgLgE2gMGdjIHLLLFhJvYGxsJWmaMxo7ZdXMtcjwpooZta4/pqz/sjPs5P7t1NdEP9
tDQQkX2KMBbwk2B/FZRp7J7dR6Yj0IxiHCqf3EDAyluBjquEFtHGP6FOzfKSp/YKfJAKeWTgXxmj
O2tlOyLHHzpH3Xv3Sh5WvyHpDQMpNgG63lSQTInPZiBolHxl3pqHdBFzpsGE0aw5DXPu5Mm6Ix7u
wW5yruSHf+zEokp2+JeZHbYBBejemtsXy54FPLmY+4lGeexniBZ5aCQHKik5UzUwX4e/ItcmNqt+
ajTZroRlk7456Z3fPLmZn7zK188NbEIQgvdIxNVHSkqD3etQxUgIaZAfpGc9GwMO4Tp9t2/zPdGf
tpP9hxDCWdxE5tAZiw2RhAR7MCUSFt+UKJTiMdg4oepBjZaIbRivWNTl5jYDOr4meJcajnzBWBy8
cZpd/Pe4R7XY2Qxxdw1TNGL5cbWnmU/741nyrcjkBn79pTM0TLHJArFh1R8hXNEoYr4td3LUPJpZ
jRnN5D6+tZZA4dRWz5FLYWejGp4hc9vy188VTssqcC3RwMN3Mjtevr/ErOCiVmLetlWjaUdLHipf
DdejEc2eYsgA5e4ehdXmnvIG8Vi0l3DlkQcFyScrsE/7j6OINOo2JEq3Pw2326BhQDhnPF5BWJe7
ZK9EVZ+Df416cigZUKnhEZAurojm076iaKHGo+osYNNF4KTsTLSdXfW++ZuFIxzBLnQflDCKmeCq
gKiko4vUXPEJRxk3+jbBnmtuYe5ee84nwOgL1v4DXcNdYKA1uYiLN0SMkGTCP4Zb1d5Z3hLhf3Jy
79fg1PT3tkjLCU83eShDERcQhFhLnMH1UxjX5W4D8okkNYdmuZ2+xO9AUKc1J023csGOk93QWoCC
g6av5znTgIgXQ0x2hBqORN8DjIWuH9HUXyBnkZbID/IaMqcTXAWafQaDF1zh3WuuLOQ1XHDqxE4H
bRttDqzhApLfRr1Boi/+pIqDgNb712rAWZyTZ60mreTRZyuAhleMh3PjZbCmf0bjU3n7hAw2AWa3
n1Y1Jf7ZNlJl8FEgq59SqQ0Q7u5x6gYOlbhPax2gFLTaSYhFnFa4TAdyZ4qS3c3uQBx4VUUpl7A5
KBIIu+qkFhcRWdy2VHTTk+n7+2tfW85DxGJXnvCfjnleIsDeRfF7qvKHxAFkcgWTclSTvwFhGV1X
dLWb+EXshXupD9Yfwy1RF0f8moHUg26gX9zFzjTbVwSN1SIQsj+Gi62X0OY/vLJy7iFIAUt+1wZL
REZUF2kfG/38sjToV+AbAI+L0uM8gl7z2WzzSiB645Vt3fzwuaT4UunHbo6xrBFUh2SN8uD2YP+F
vSk+Gzqg/8/2k17evABFFOY52lfzIqMu6K8flUe4qnmmc7BQks/CQK7rQ+9wjkjDBdExyOInP6TW
KTfl1EkdA1nTb+3AsOKF1pqVYX28OSSmdCeFhNNKWNIsk9o9uiGHOaielLr16wIhQZ198CvWJhki
x+awy1TIoBiI2jXaUNrBuyPP0tflmEM0JaSwAvk+bmYzlC9Hj8mr0Hyc5lgtLhMtXedrHb0wlRFr
52KLGy+1nbjiY9FQoXJE/D27O5Z2IXrEjAeF19MjYd3HkYtKbfiR3wBQ3P30JTzDB/Bxnu/UhQYV
nhp0U/hyiX7eNuO9RssKPfkTvI71jDsreR/fqta1JriKe/PyMvHMN/858G3nHSvI6afOFnwVsJSa
bLAsAZTqUqso6l4lo8Wj4rUnduiLUpu/71lpmUI6bKzFX4RjVDsuO3/08aWgqyWZPq0mVEGtIagT
3q2Mi61yduWq3duiytVvcyys3+Y9wVtJsNi52udRqtX/xEZ64iZ3e4HcruPhEbAOVOy5+xwAL1mZ
rNEteK1AeZ0miR7CTR64o9QDPlH2Vm0CGBa2V37+NbpPHqmNqbluw/Ea+YMCI5+BrTGxgaph0Vj4
zS6VU5ycypydQpJqifGLwtrZ5NmbWRfG+oa0jQAKffL3uiz2HcV5+sUPteiTcCg/ffR+K4UCu4pK
nBH6S/IbLEl1fdS/a9u9wePlaa7LJ6ayBDPtoeKIlJOc+r+O7l3VVpMfXyQwCUsD8cF2gsSrTnLB
kxXB9koj4dHBB5TEm/8lQjuVTSoEyA2IFRfehgwlaEEsYohpcsUaiQiDef4qltYv/4sFERUGW4M7
N+JIau4RjGmRAoScRaD8pjNd8mlv52HLux3dGAFEvAcbxRGCzU6ZRr4lTtgaQ4UYE5iKMP/5JL2S
uh/ANAAtS6ZipKsQZEMFsra2lM946J2NjcCiFXSRnp4qNLJqWaIEqil8GLK/K9RXe/xKa2ITGsf5
pKrMDafG9PLOuIExxbom63JsJm9qa4o4aBG/d+Yrlcozc/w/VOl+au5GqXjV2Y39Kkdh6fzeZufl
PC0+4S55sYnNyTx+cGOi3faNd1qyqqQ8N1XA7+shxlCDvQaautG/32HRbIjIC0AJ8B4B4gGIQ/Fy
RbT9VrKx7tFP11DTlv7G2zcYPTsfbou4TOeGOTtSIf/ENZEulW+NeK5HcTFwuUqzpjeGDkkbwqEV
sJlTRBSkfyFcireYdr/Py99BNTdFBW/xLdVj2wUj6WI1ZDEw6wqzxmOoHOnrZ6clwLRGCRd+CpvD
adXlT26rinNdHyGNkR1HyDobVXEf8PzfW2V/oqJz9xI7MYR8nXNecYscE24D8SgASp5yEB27oIRH
NY72o0fOLZnDHckO/xXrqs2gaRKomNRdJqi/6+MkgGb0d/fYDyrhPIvQyZ4FBJsIzX/6/dpDyzse
0F7mITixxEY2D4QOU2I1uYnrSovehVkpgz8hduilDCz1GoKGzmUkpTb5dwJSXeMzVspvigdEV6iS
s01fbGyoKteg9snhdUrx7uRXVY27X6TrfhF4MZ9njsT5tgh6B9KXS0/1DRu48YqjaV06krJA5z47
LINoOePIRxjuz/TBMW4m/PFjLJa8YL3CLJX3zpeMIsJZ/XAkx0MSkZFo5ALVOYwYChryUtiM91xC
/6hHr+G/ExXdJ2SmWwbRPR+WItOh6UEFcx4P5nkAOEq8HpB5o68YVpGItMxr5KbUTW6DLkyS1cQD
u4RQYYo5dXSa615P3ux6CbSnRIrR5U5DQNwKS76lfWkpTDKskyvoyCbu4g4L7bC1osBecoSR5Mkw
YWCe6Np8g4JX/lGezz3MskZQ22DjhXvcOWiyR/bp8E+A2yNGUiI8ZO6Ul0IMWyt9Na/n0w7pb+NU
LGlUYPnfNOHhwQsHpAHosp15DAxh7ovKgwb+Eev9x8fD1WHkqOzxCE4Txp9VKCyL19DJA/iBYe7N
i13njdvNzznN80s6/g9LLjfwJRxV99IWllNxPibUS0CLvVirNMewrCk9ttp2K8TJEXOxrEAJXYtX
6BwmaHVAktKBztWsh/T1Ezwf9ygi5U7FprjYS1R/Vs/5pDSfP5UWw40yiW6SndnvvcuP1DumGv2X
fQVD9e4EWZLOQGfFxW6zAJiSpPQ+TGoB+NGERElqrpQWHRsw3aLvrEs0Z1zYzAJxGl85nAcB2Kzu
Ej8qZwRKDuMumCKfIy5fLwbw1fOHTbvf9oJe0ZqSqkvLAcMmQkpcLDcgdsWkp5ZhbOWob5CbXD3K
j8j0pjZ/okeC9L5q1IkmW/yHRHPZawkZe/EcNESNV/YCQFi22av4R+1wihWTRqOdWC04NIP8PUt/
iEZljipQAtBs8L8CnoImzYO07QV/ognpeDtH95Bj7eWi9RNXEnFsv5ye2PxFn6EQ7/U3CshB4xJE
FlYx73Mu5FcrLSRf7NEn3EUJmODZqqQqf1WSRsdYeGCLAi5Gc5N7mGOSBwvYJKUDDboFUswMyFJc
1J7L7jiJprXXB7NGcPV9tphTelF8fNIdzXFaVbUbXzU3uBQcXmLnRrIoxxTy/f9CY0Wn9Gjejo31
boc+km0GGjSY5C6piE1CgpLV+IrF9DFsQKH2LOhjFX4jIpl9v7v2Req/LNsUOJQ8fleMZpKE09Iz
iFou8pkGUgFY9GD25hV7F97StMS/fJvYIezIFXLrLJkj72xW5NwDoZazoY90mxxw9jK9E6vhCJ9x
0sLRCecDGKCCmatpAaSRIPSuSoJbwNqWV38QZRnjnb38g7X+baYJ/WfpFqHuraI2waKTNNiND0oo
QandZP/uZIPgYu+qYSjemZNP2PBrsQ8gFAVF1zYujsRNuoU0mKiHAp08SC3HSZp1OP/fXWi1E3i+
ZwphysFVBkSi9gFw8+GteQriPB6GV/Mn9xMe+l9lxobpWK3QavGzQ5JkorA+Sjp2hrIUDRNgusCG
j6SE4BSoyeX6mcrBNjVYRbz/Wgixgo3T/uF0gE3zIAddutmVoXQXl0a4Qe2GD9eUgjwDmJYA9lqF
RJWbXgDlR9Q8BSdL3+0zXA3EL3Eu2MHyYt1kuY0HM9fE3X4lyct6/ihN9u44Art1Obiy52Ku9XNK
79rBG0wwsRnYZ0BxG1F19R6Vl8HQiM7MWkCBfF/VHJiMQQxXZjDQV+89DsCjR++w5WNnwObEgT9V
ed4g2kh6h8Vkn09LXPunmWOZVWsVImytAdRFCADfGEswRdhXSKa6KjOofOjx5V6rqJx5Zyrm+Ylk
r0l1QwypBcwfON9Ylci1BMa4imoU887qBILz5AjtsSW+Dc4wtqzXu3oxW+EfkUSz+bw7Sr1mNtnw
R5NBwwAlp8sR2ALWgXDfBtUCh4SNZVdrmng84sKfB9HEzWSwKWY8IlzeKHMaeD0oqF3Y8vYptqEs
mhmaH9Az6Jvju6zLvSJExGzJjshhxHeU7mrqzM235bBoxVUwi1Ukqz6CS2gu2IAT3RDALTqMAQkW
TfjedHknVu2wcBZA5t6dJvR8tgCwBGDQLtY6Vt+jNKDU3cNoux3gU1h2ejxswWRmVE1fftAvoD9B
uGmkSgbJvak8dRcCIgJF9mgQw+VI2UgouKaktIeDqmbVwOw30cUCh0hJAV18KmGMpZzGVHaeHncH
loUfvEWcTF9DeUqWzB+BA0RQ1PwxB2HEwg8ZCBOmzp7yC2gbxnLHKhVtdufNZdoeQu3V+I7ljFsp
LPEbHuXrpKnZ5uxZqHpwgzYW9/JifdWn7fG7KrEVLzBqx3zi8X5Eo6zkgqxXBZEbLdoaT+KfIfc8
+w8oxFX3n9T0eqhwwMHMS289nm7fnxGQuOCp2NbgUAodMGrcdwPhCe/UnjiOOCztk6RXBjjvJi1t
N8zGs4DFeh9vOye/eLNaJGjR/jjFGIAlyUhEdIlnf3TkQix2JmrYhyFER4kLvPMfQeDSuD2h4kLO
5fCCmNV3AIbKlhBK2PIHNn9jZpkho3J0X+/bDGnkFKRyUF5qCTnI+cPcPbCYyJ8AeT42xzfY5J4I
BC47Sm3HqNZ72lumpHmnmRBBSlvh1WXxPGyF00EevxVkiyFZ6S8yXm7uPAvmS35YOrBTILtQTCo3
Lkdie8imVdQIpQ5uWszc8aKH0TIeG3/sOXtgjMYQtCYF0fdm9Gv1JsFMJjaNTjgsCCjK88AEPwsS
3cEmf7QR1NF5f6001pt0YqP+mnHq+bsbc77rDb9mGwuDmrWHZm5MprsN2kHp2jNCRox8VkD/CkAZ
Rmrt/0Bl2n/3PZUEmZvCT0AB+bTVF9oZHKmMBxj3/A4Sup0kKo20bGrrXmUIgF3hS/zf/t/n5so1
RMZx3KYuvld0B76ZGRrrqjMAdhIYQULPmDLoAv0ZbaJ6VO3kJEot5YnrXEiC8vNHVWkkgsiyNdNQ
U5ZEKb/Y0vUk7Bz3LFogdT/AHZi+2wuCVm7rfY+82msOxPepk3xIhxNt+C0ZAHtHGVZAOAdVnHri
2f/wUP9UIpZ1t3xVQ3gHvrRhTUOUSJLyllfD96JJwN8zaJ1EWxUtQdDEEw7BHmlR6v+Q9wwp0WmX
whM1TWnDMQ/KIU7BAipdAj+PmnJ00cQ91OCiTcufBma9SSDsXr1keHD5cNWXdCiSkd/MNyLYtk4k
ELQJbcKbWBDi+ygJ2iBrwEy0BLh9UW64aEjharGx+fcw+FUbmegrF4wh6gBMZNdmUTkXHLXSyq5H
xQRZJa4m46XZlO2b94iesy5g45n08/OwCGN5n7ZrqxgZr2ZCuANoZVu76nfCpw6RegI2Ch6b11VC
29XoJmL4gBObgZMiRLsWKBLSIZeqVuK9CSrldrwXsm1xSSPZlk5NpkD3Wk+jPfNt7YEZakzGq8qf
GWCGd0birwO+oNuZ1Zf13qwdKR3yLkJLh6t/XQTYWceNdGXWvhELZYo7k4a7higvhUjB6dzf5SSM
eFag0g7FSF7fsC43X+Hi90wiUaAaQU3kl8oXXAOqR0G9PHFrCu++CChtuNiCI1npMWUpnFiVq37o
lOSAX/Pl+Hnau3pAM/Va2/iIRsNPPEb7nf5vaZHKtAmoE2FBRCOTmparz1nQW/KAQrK+R/ZRtuCB
UzsGVp5jIeeRQtsuA7NC8sWMrFyksHCY2p6T/RIeVjk9L8l111pOyPoVa7h6vaJK6DKJzHUGyieR
lkRh7++OLJwHwGGZTFmTYctZN66hVjXIfjED8OOb3h5aojTAK+qUXVpVLNtYDfDHQ8DnDnNt3zo7
khrWuoNkAikxCTLIiDjZRME3bJ+MWhZZsE8k4ImdlgfzXkqLbBst9TOmfqkDrIeM9rmq6I/4Dta7
VMB+b2P3eNJvG28OxV3t7ZwcOlQ9DmlL/kQ3lI+YElC6xnG/AK1TIRE4amBsfM//kk/FM8LP6QFh
wGqiX4Z72my1CsHHHJYzcOSSdFM0k2FHwSApiXh6LUkzgHJtOqs69OgwODhr1ftuMCqxeXpA/42v
1uWGb6XCXRjNBqPHRpN91o9J7LvlRJ/JPMQyDqGId0woI0DXbfGIaxJs9ysiJOEt4Pi2YYHEfdU0
33ivnj1PWg2IHw41Aq54Vuzlixak55hx2Vy39C0yt2BbH+Z1H1EO1Gi0xI28naszBcpAb2WKFdm6
0OpVTDlKi8lo4ZYxeWfIs6O3fe9tBxuPbQJ0hL6xpSFPQtgUyD6Foj1OWoIYXPo7gb61ZJjIswIp
XEe5tgM1mcMeQkLEybfHb41EYen83/6vejryogH85IJqdLpoFIWo/Y3vieO4YEkxClsDov/SCacL
6ucKqKYEDFFqIQTTOj3PdeODw3ZXGts9kOn5p6bbX5fRx70qc1vU4FKzrTLyVuC0b6sr/RY2gq20
irFk2+coFNy4YNsy8ymCnV7aej5cr+zFIM7bb43LYmLi4rVUsc5v2iHy5zQxvWplqnQMroKncolb
sh4/Oz08nnPu6NlalpKv514Wyr9FY9NisxIHiuLHb4ey5tY9fbUqXBt2POb3NucmwGGbCw+mRbJc
u6R84XlPbldY5ZZg1jcfhV6Yibdr+lTeZOkMrbcIboSVcUipBZajzhyKXPMTL/6kt4dMyAcwpzyN
7lCqS9UcTSlUbAPOek20+LQp2aw+ZvhYQ2anQ1SzR8mAOPICsgc4YwZ/7cv7z3VnsrfQTHeOS1rN
aPDUbrsr07rEW+ydAawqn/TnL1QkDQReMlcbysX3kbovblaOxyHOYsuu4YHyeoh+089zE9BHVjvY
fYrcukgtT+5RvquvyrrnXaf+puMmYKSJpmWwHeHiIu9/il+O+nJloR7gZBX48D312iw+FlNA0Qwq
32/wVt9RafLKa5sB5uKwYt335N+oR0lWQLuFSKFT4VSPBtuuEDKC4LpUzzzoFa9iWR20in7EwqZG
7BhD6xEJpGF7PhEjaerHXvuw0wKJSP66GA5Claky0EsWIr2lWkdmwc41ESenyOqMN32wN8R5g8ss
LtF3Pc6qc2khjvCcRJtf64xDRO7HxbYmzLxDTlXYCdyS19Pcf7K4iMGkoCrBk1KSqeZYQouKKFLO
KcV0XMqtu/c73Ix39avPKlYXsEy0JpU2y7cmt3WWRGKhWNJ8HgqtaNR5xl7MRvqLe2zGGSaOfluM
VfD7y04bTW5ngtYFUAeKOqWJSZQ9VLu4ZatTxizeROZj2VDr2km4RdF6DSfByrqiuwticDBww995
Qq80kieGjgdf8UBACEomJKczAEsG+MdphoYhpW78rjzfGJSL2A5ZQ5dMNGvmbPAdeXH9ny+RmGE6
Ob6zQJbkQWSh6AmdFKcxw91DdXEg3fPLMPiGNi1IWluK7kWoE6Mg1mPbL43BeNgx/7dT00GqdN+m
q1Im8tkcrH0S+XgY9DttmBQ+rFs1Qq9gj8tkZSEomo1dtIuOQu02RwCRWZpcqTqfJikGALBB+lDS
/IyExdN5FVceJEd1SmjDal3MxarYoqJ0DxMBzCoZfyyG1j1fLwvO36B7E0TUJmC8ZMG/CnR0KkzA
YJ+cyWd45+9pIzin7i3N8tNcrefL739hb5Q2tEuntQ3v97/7FgK2YFxxWigePM+Ydk2PRy7JoekT
GmDeC0ysF7m6iN+Oh1xj2/kNKTwqg7xcQx8BOUcl92xnO8pDC6IlOSmLZ4YjLJzAVK/f9qIU6H1f
Vm+aGC5cAivE3bUp2+HjkcnrJSivzmfj9sIuDtiUnWZHaeQWU1F35G8jnd2y6Jz0LzNGmI3LiZ9X
9anFY6bDBG+4OkNI1JeDk6u3N1sw94vdoBDtMx4+YNOyZNzS0lv6W9TR2s7gwNfG0EeN0aywNy3B
DTcsJpStJxKt9neNaWUdX8G5rgGu8UxBnADWCwLRGsh9ud+Si6QuNWODPTV4SP3jDOp9nIb1BbgK
lRA2HyvYcrR55wwNEOGhwGrkKX5/fTWRcGJXNL6/z4WgkMuIuXM1dJMhR2wWqrrXKRu3n/aH0E+e
8Odud8c2ptFJiEQjOAGHvD16gonsZ685y/5VPAh/lPUJlWABk48to6qQb2IZpouKArklDChfWRi7
0DhAMqvkbOZSZMOWPgVPfbB0IUN3mZbcbuxsotMOt1ZrQ9cXlBPcwerKsHBGyfBtynk8GS4tNcuO
+GanPin73XhNvBu/MfTXh3d+O7HM7LdhFOI1h+Per2SzVTDj+yoF0ScvPAQ2VhiEfwdXN9QxemXN
ZIdOTDk59xPI1h3taRmZho3Vd+nugCRaJr9iusSTJ6JLEUUvzidWs+wnpjo3oKxDJrvWKKFO0FI8
FODjPctg5elSrPSZ6VAbE8PwmzN1ATU3/vCZqxxEhE5feXzSoJE/WCODQo6iRmtyFLlKeSHWpYUa
z4wm51bPOtAcZgx6XAN29TR7HOZxTOw2Nd2/nRwMkT1uz1UQW/zzun6J53scbthcFnzwljnVKPg3
S1Ki1HL2GILk/G0NLGzvovmfl/dAb7bnmSd407YOdaQVslsx1GMZwoORah4gtnhExRTVub57PkTH
eCHiPGGXeGaeWY6mE8XllsTsWOJ1ipWyfSieG2LW3HEc+OwZ9xVyo9xj9BRa0qJlBd5/5mnxJTFH
0y2rgnk/AIdY3tGTT+nEhijWpeLmint1oiELFAIYkYkbvlG+1TRpWqgSgoB0JjNhfdQVhGvvZfhq
uCfeVJOVgY3ioocxgECI8ddPN5W8PRqVsOqEkQ9UOkYtWqF3TiZeubdODT/qmKGEh9DKKNqZDvWj
/BiBNDeKuVDxjseYhfhWgujJ7rJq0469VXJ4w/G4n3rA5a572tu/07T74H8IDt0zQHazWrnre5pl
jZIwU9W3UYoyQpbPncJlIbMMx2eYnUGsU9/NSltqNlBKeramLSz7wrKmD6Jy8EWMCukmgZXRW6Ge
eD59OCbdZXTPZs9bNcgQv/kM7UDiLWIVoka/vfyC3Ahsxbrf9Ot4+lLKCZ2Bk2mEN/UH1Lbvmgn0
E3UQ1V/LCs8nKz/s17SpiwS+ZI7c0InH7tGka3SwkXAf11H/Skv4wMx5vu/2kdm8VjllbMn1neQt
G1W6flnnSbT5GaZ9Y7e/1nChWRsTgnM4AhJ1pyaZa1SHtHZetJ35qxM5CU9SifhdXd8MZQce8Es2
g5xeN5iVJXTDElF8a81IFPH9wouqjBnCbVTKf1aWtoIP0k1wAk7DGsJv9Mxle1aW+UfNQVjAKnLU
gD/M4KwBQTzUM2TC1mqJwZ7FuVUkH08DKiQhplJ27NYtc49mbZUSDoe4NJKGfulIshgdqY1/pOEe
75Zy98lBaDxlTFjOTf5/NQRNFzkqweA8zHsy9pwMErN1KdMcwGTLqmV3pnpM553qVosPwQVuOAAS
GHsSTSYBfoYgpnIXnn5pzAkm6d1mTnP4kB5YbObwR40gVgb+H1XFdB5NotbMxOGa1eRj8Q2MTwUo
ajUo+3eHVMHk+ZyU9YBJrNQM3ZAhNTpvUtWgOkvOFz2tMBTRar2/V819r+bud549qaZ1EIpRPQT1
2s2ai1JbB9faL0gkeLZ9WU/jjpNVskGR7Sd+By2biK5ZJbLwajC/q6TevW3gL2M7H4lBbj5NnR5U
zMjAVTkyAk0HH4l5QXr30j23UmZ1eKBkNR+eFK0avgT2FhEcZ/wfeXkA9bT53Z1LDdMEFSxH0vjx
L17DEAK6Ig/Rf+c2N8bOX9q7GdfyFRKpjp9NtAzEt0QbM4gOcLoL4UeTXK3nq68vyVbgd28CZHe5
f9B5+NNU/7WDl7Eku2OxHxhhX08vFdJ8oxqUzUnE8b3OQlV+nYlaS4+GML843t3NcK6sqyeR2erZ
HIgMYxQBjuy8pnE9klndNxOOEscCtqeS4N6PLu43sUcOGWgP1ANzJ1+gJd2bTZ49lAlZNQEDe4QI
yYxj8Joh38fLpyC8HuI5CVyzrKAzQKyG8qa4e9IOHVbfGMIyLJjFmoVS243G98e8TMdT7sg77T3l
qhhLP6Huo3I3REsjtKdHwBj2vY96WTe+Ir5RYvHteuiraRo7C8RxFh6+qUOPqRofk2ZUvjIrMnzG
JZn1HbD1UE9UHz18tQsCTleym77fkyLrf9MTTxtXatOCqYeLy944+H1gxeN+FXNbRpSaMFH3zS4v
CcCQFOIm0h5XXpRVKMIKPWsjkouE5tkxhpU+gEKwQaFxHogTitLtaxUGyTuRfxtlGcJVL43ByRQH
fLqab8/RTkkHP20bkVOk/bVWB6yCo6xiCqTlHJBjaqTT+QiXT0OunC6ACEqQ+tAimRyTuz3YW9gM
3BiQo7ZjiAhgPnUY1++8O3EEhM0m3v+jLCCrkocEB3/5RV/VfKa3U1lACwZae1fkUkSsI4U2g4HJ
cwei1NIvd2ILp4B9pKvx0WcE+80e8ed3rcjJkIPa+4HiDblDx35HOGyt4xFsvzJCXWd+VPHkjXW5
28TmcdysXRW01i54hSmmcZKPg8y2bBE01NksfbBMD5n4N0NeBp6/Pzj2ZpGHqXACb0EaMlq9yeGZ
FhtiZBkai4uCSp0FAZdJZA9YaRGf0tqebqa1fshYRF989FvQQ5WIrCYC4zA0BtnF1FjmxW7x8fV0
kAbymwS12vWv0T5pygrhI6fcuxc3IeXHy2Ud5b4XD2/XnvcfndJPawO/oZD4Gq7N5LND+y+Oe+d+
8dkB6tE7SSGcVU/OyYrm1etTVjeU9BoI+hdjUjClNGkJiMoQkxd4zFoS+D0bPjh4ifG0cqvmUZ18
kY22M7g3ASMDgXOaP+ToLP+GRclUco/snt7DHB3TXjcqJIlyMXi+4IipxA48K84xCvy5D/736RaA
qmQogXmabvOYBNnC5mdAuCM8YjFyd1/RT4aftRsvZrxsx2iZCZOiVT0suvBfD+5uHq2nAYDBCBb/
6dY9dYTAiBkP7TCFvqVJj5Bd0gAKnvDmmFvhJ4CoyI3A2cQQ5dIEuofVJNomJHcH7PPok4m3YFho
ktQneCYjZ0ZKUOb0Watxhzgx2E27Ig/DO8KjkI2EHyQLjf9ZhcrJvz+6Mbnll1AQA5mwt5d0L9gv
/IbfXA5ZWTGCR1bk3cxnOOxiwC8XzxRiJdh+fWcYzus0/sZ8VDu6pj8aPPfEKDLdLulgD0Btxwb2
SsCuLmPYLbUnTIoXlf8sX2Q8lf5WQX3eSMCxh1blcloj/kia26chKuRK7JGvJLZ0WGURWHxF2lTz
C1quqxbjyI5sDL2AJ/p4oXffU9/GhxSuLEBAVD5ol2lGtBg/UtkDERr2ZYLfTYXebUz2s4xh0Khc
hJziQwKausLTwvySrBYVnyBzVdzJrnkZfTFro/qp6R23P5u+kZGC86FV1AVyn7ryWWl6AL7gCNwE
+lE8JaH4DryKPRf5DVTtsDBir5Io+yJDAYbJilKvoMxKNlQjqINTAejbguqDBpq3/dYoSvSc/SKS
y09Wubop3sARFLtWkPYy9f11IusPMxgwSYi2dSmQAPDP/zR2up0XEeCL58DAWoRghmt1gL12kzUa
HEVRgphdPWLrSeyLvd2jrM23ZOvP5OuWftqvBEo6O+RtMNEdtlCLqKCC8BC2a7umbaowTu5oV0PG
sBgB1qBHXcDrQT0bJ7eyha3Q+lKdYpy5XT1q0EN6VvL6OOyxVbW9Kkd1lKUNkQwiaCFE7ZobJOjC
kWXOGStdgJVdj8+xG6kgJFu5qZ/NSAxc8Qcdrn3+PsvBYHbSz/14Q21pQPcBa2HkKueSN7fsIohK
V3zAD7+7CAP7RD2jh9Cu/nxLO3PMo2wTakYUYaShlILB9SkgCq5PAmqx3/yupfv258957WMZu9IA
qBe/ol4Jo02Wh5TWOJCY3HImIhW4JXfvQaglpFEwM1zJJ+Q+NsURueHvJDkpjgBEU1V+RGLFHOsG
Pgr3XGgtNIMO26JrfX9+Rkvk3iSsUrX36JvIZXnFSYAxPTgVokmuAOjB2X5TeESMWbhumeymzKKV
GlT6n5654INEnyj9AGwgQdCFJYFxVi50ympRv5VnlZutSy5O8QFmLQhIlq5tCVQGxhce8ZwNjvQy
gG6Trhb0o1NnjLyVC0bcFF1NdSQBKDhbVUeN3Y079CH6ycrW9n72/kI2c4h2I2786n7lx2oKZVgU
21CkJfFnuWZ2MWHVrzSxDl9ko45xUDW2YmxitFdtB03QEkp2ijHTZ98zihrutnK2fFsmvmMGxxR2
f+pIp8gmV3zTw9a4nclR3s/sH/Wuy4p/eAGfVSOBn7KhMgHmX2kZru+2ZA2I0G1mm+gv58kXm94j
/fIi4X+dywvGRWUYB1/fhxGFJxRkXNxlvnrxKkRwNsBQMrdQnf9fGdJhPB2PSY+OY0/NfiOsyM1N
VzzRkVuDSPGRn6JZBEqp3z8lbdnPoeMjAqt3XevE/arhEYKOJOnPdlYDsf3xKUKcPbtmnNI4pqkO
VtADVXGiV7QBzMBoSf9RK6rLcJwM0+ku9oizT2iRdC5cje+NtFhfX4e75ErRdF2S238uEfQU6NKE
CIq9vM1z5HXVYhdiuVdXNl86KMRN7dYzqoNFphs6+O3V+e4+3kKDRfIq4iMT1xQc1ZjcuikFnX43
DIXeR6/4rLlTj2jmFSlFKY732t9EPTwZsBm+p5ShqHD+D5s8oiym8kVQ8VTeLPx9GueG9pLbz3Kf
zUB1nlfugVXhfebXBgRAawLxPHlLbg9qLo821Gu8pKz0ePRDBSwTRpUL6KmvUzVsYX0RgUiCoNQv
LhDS++7QTEfNyWZaVOcu7sIWZtyiOterkki4YGiYMGYXMXQ+U8MqdHlbyFIFyqQwsMEodM83DNOg
R2hI4eC5fOeTvJgYi+oBDAcYABm60ecQeyRwKLMWW1255a4wcpTsFjChljDK04bRG8+xsyNJlyU5
OjItAShR+CvFMbFWbA4NbZLaIY1yQCbgZ+ITA5mSywtIDcMqE6Mr+/sAALLDRrKrcLibrfT/Lcav
tXUrra/9j0l/z4itDmhALDegDQuaaRHVTCpBaFAeipHoKtzvOoy01ANgv3D2ZzlntZ8Zo99JmSGj
Y2WSVFiVcDTKWsCQ5BSYrg/XV5AkMGdTJIFSiEU9dVGy8ayzU6qmdNlsKUdA6Rbxzt55pySG0Ryf
iL1xIdm7RZC51RPHlGFAhz4OJGXQkRmaKnEhLjyE/kpdZFSh6Z5jOPqA7QjhYCbx6gXfS5QqNN3F
1Pnp/I1CKUtHUB1qjBdisvSwA/D3bWb8UdO/XRjLx4Rzn/l0F+lMytePSqCGKE7IMo7yvmy89Moa
s/KDPog9QNiBd0TzIwPN3vNG3hrY1pzY1JkjGJxkE6di3kaDG6Ca8XmpLfBAS7ko0HmEzuSYVN/x
sSlWy45YpUR1A5m0ksnb8vH9QTGz4aEWPU9els5CSxINcxv/xGk7OKtZi5I+BT+YRCe6iuvkfUF2
+ar7hLzR03ajXEIEUIPrFOLEZQLOn2Zee/IR3iF0rvDAifa3peu4n1xKY7UlOshivTMPm49LzytZ
OXMDg2OqFASe69WT7ry9jGHdi2ISo4RbPgAwRRXB/Sbu1Kki7Pmq4OSo8Ccb08vbid4mWyKZINJM
ekZUd1wgW9tIjfNyxtUwXTZ+nytZ2XRyGB5wyQhgBWrpesFqJ8TTTaH/wx39nsZhYA7CTLY1zQpZ
SWP1hjcFnop/BOgk59hb2OB2cH4MVG+jgfDWfl7f6VCnZ0fEKoJ6GJOblOGL+Lt53YzZoCywohHZ
Ow/W8soz/s8hE4Kit4Qne3HkG9RgwSnlRrqrdjCepKxVdH+GONg8iTPZXS9KGDSLnFYha07+PwK0
BQRupZt45CFuX3eI7aU1RM3dZBzGA3yGZfwRbmqjeB69fm2RbFrhURQCNpmELStVmhW5HOuf68jK
7VkxF+y729ubjnwxiVSkk33FbZLVi4zwoTTcRZ7BHrdhSJr/eACbcPOSA1MeMsuSyWC8mREFoovY
macOPLjIZF70FgaomvQ1AwzXylDtP3oyT7lLOZ4Y/T8ijGQCNjAOn+R7Fegtboail20vThmrp13b
uKc/xclugBSnOZyeiZbkV/JpEvxnuSLAg4VPFU2LvsIiL9ThRzn0N0cYpyQQG1FwBqcOcknvPDc9
GCR2lokyRPAKH4tQK14FI/mApb6Paau5UBtd4dAO4zv5O8KkSGXPCAXvy4lQ4HuLmX5wesT6LRc2
Zdw81keeBN/zwKIwyK+zMKq7/dnXkWHRfsAb33LQZuFnQel9ZtL+ob8/ecIajwunmielxCraZeyC
nAwhec39c9rcYEzmYl6gUjwo9AYZ52GcVGmVwBtlKQipNEw6FJKff4qDHW/4NMzBEVHabdzog8pw
3Hnu+30m7OVOQMlftnGiD9AY5JtBUTY/FeFsVTEAfuJz4C+7V75WQCnwp2YJO3h4+zVJrQJkTuDu
DCmWobcgilXwUhlMIzdXhd1jKzIwXPm1OZesGEM3YPmTonaqvI1iXlYSgc7TjJ+ocAd5RbPHMcyJ
W+XMF2+FeTJsIfxy0qDcHgcEiPSm3AoKreHKWuPjnhzZ9w/b5rg8cP++5Vh3tnYurRmaiyfHdUO6
PuudDtOIXW5YmfiIU6v+MtAP5Br3M2zJ8gE5FtcKaJXTNmgL30WgRuhSzzdTclpgqZJMysNWXyh/
dAmSSvDkvLkxUEPOvAQzHQe80XVCzgNYvAouC5kn+XuAp5MPBlJWCTpKq6Gcjnk+j0VTrkot+XnF
CAzJDbyVshQCRjDH83wwJr60AFXumYLmnqo+uyC7YH6kgmj+/y2SLDBSR+NriQxcEWRZBYFt021E
K3nbSYDjx5grIgfdDW9J/X+EwRjceKMFDfrmZNhejZ0JJK3S7mGEWY9My3HOy0KAJCTgyKSwpIsE
V2LgfSXfhE/rcFfDvSLFrClKYQjW01Atcd0S9o4nKKzxLmgSWDqJZ4F3ocafAEjmkqOAzEMfVbzu
FX4FCcj/BD46WsiHkR47xkX45h5W3kR92AVrOd+MR4ksGf5f5WJ+DHtY7+rXyw8hZvXPARR1hrH6
NUv58jB5qbWKhwC3R3YVdZ6MdM8lYD8jOMfKkixH7x0dp8XU9n7EE5OxVAaSLZA5dID7FfroqZex
oVy+p2Zu1Z1uvlSKestuNVEOcnG1zj3WXU77rXBOx3bhRkp9ggeYFxDDmSbQoxDP2oBEFwrn5Uk8
959Q4mNFKpblHzRl6H903PHDudb2YxYfgOOD0Tit5I0JI9QYbiqZcr4c3CeL0ISHVYV6iLJQeAzc
6wawTbMZJ+Jrfdhq55ehmNZTFIt9xaLZaREurx5yhtoSgOECQSIjQByUpr0hepar8tA29Yd+oYVN
O3O235Z2Nc7eBF9yBT0tL5p4I4NDk/lGwy4GxuLkwGoB2f34xqD5IUFSWI4LJvJE/2n2iosIORRt
CeM9uyiu5S8GFihf/SkOvVdeCBMl+e3RQJnVe08ied1ZOWKsp4QdjfinIqbpdZRyrIw+9hWHlHjG
22a7qyJPfrs19QslTDTWe7s7rlMo5f/oWOUeTjmgdhWac0dCtUJuTt9uynhBfcbhoMlyjlJbPdJM
IFRmizjsbbVVFPYeRFmvxl7wENwMj1IgFsiwhDF+c65qx+ExeQ+AojZFc4qxtQABG2l9CpcV8Gy4
VuB6QrAk3nu52k3aJDubPWpLEWTWnQqXp8C/4FIJmtvxCenETjDXh/w8Tdtqd9jltJ+uJBOtwSId
EEp0bOe/93Q0LE1kRoE/68c/L71VBWvUly0n1XkVhbYgJgyTlO55ATKQY5Xc9gOrG6dp29BK98dl
ytOdPaJJn8zN2TzZgx495Yc18brCJcjFjvZZtozvsxZUSrmxrCZhLIDpfSfZqZSTEQhQ7t5JTd/i
tXDADcv4i7iBSceCNuEUUy4YI7xKhI6YrBKmXxbdrDnfahjDV4+zY0889Tk0Iw8nayuIsoHpbJ2J
Mqy0js+J7mT7U0FHe0AbaZGDBOQselH1zdLmRdg4JClxNgjHoaf2pdCozsw1qiOlKyI3iUhEhmUF
cFGfYHyPASNnpj/wSQhEpNWgEQfbvM/cg1psOa6/prveefaxVC7Xw+XtH8WvWGW86WCG+PokJmxZ
YeNw+DLDN6Jyw2z3MmZlKzdzD0HxPb5OGtO2K/reZ1lnp8WieqC7KweoH121IdzgDhKIb9exyMzr
cBp9GRPuN90PtOhUbkqcqBiKuqUIXUByKfCgMTQNtlL5dRkjT4nreCEt+0UcC3/RcY08/kyl1fcs
VXnE2xoaeiUT1v/t+bBX40coCjROytlo8WXMEX31JMxfOrOvP1t6BiVI6P7/xVwzq6HCr/WwqKTL
bIqkVgWMx+FRuKiT7iiXUwOOQ2L76IoLxf/fWQO8XNqiHMtvr4H+7U9H0jOTQrXOBu1/mlzjRwis
o88MmlykBlyQ//fYWMGvo/hdT7I/42FiLooila+HFsJG1P/3Y22ZzuDvy1lJKaEL2O+nlQIid9XG
4yEW7UIm9pGl8FTP2J3to0ohMQpHfT7V41GhBs6/ykXALWp6Fce66e/Z84Obx8iiNsf/pX4w/HLc
jOVxfr/BLCLx1bENX1BOG+1jwqmEhGfd15Im8pBWhQocQTsnFdeiwLGf+9yfaLkrNLI/kTa8CoOn
4QesCuCRRrmBjAE1PWJSyo8aSyeyzrE9RnF4E4krleCW/sLgHVauPzvtMiE7ndod77v8HQd6WGOX
ZXyd38pTS1ksyxpAQl9oGavCzuj/f5ucrBlmxIcpIZbCm7MC2C+2RuoWrsMPgx/CdPPeyBLxP3G5
8gznY0bldotbhO9n6V0JNQ4G9uSFdmzUGlkYLJHD05iX1HGrkL9sue8/UnIGBgVo2DuGgalB70Yu
W78OZoaXr/8PK18mSK+FZu0dAKzkb2efkAB7P4YF6OL/BRixpJaxLKxuA0dxJu3YLzwETFDEwZnh
HHTp7vDAsUQi7cVJffDG2HKtJYzPhx52aM0kOCuGmJzzi3hW7pc0kn7A1T2wHPoq5suPvwnxBKTf
1s+BJKbyH999yqCvLa8CUKSNSEX0ah95M8jyWXT+769i7i6WJTCZPNeC3lWHCxwKoWK/o6JphsKT
ZLzi6NA4fJGpoJNJ4S80sVSd7sfSCOBIGBlP3zG0Cv4CvOdv3e7bQl3E5PAvuFEtrbVcLdGstd5p
zVH2BrzsJSlgZ1dKNayJzT4GhdfK+MQ5Htg3tNhRgqGgDtEYlct7ijKOzAx+sKq9OTpudR3XQM1A
OGrAENupI35hnGgp/qV7l5oDY+V5k/6cpYjqK/e60IvQIvwHIFg26+bEbAREF2IXbN6VjNS3sPjv
svHvSfKpN20TWDxcER9Pj3+KqSuP0z6/oGBrf5qPf7sKMu3GBD/OutXwfrjQHWmgfRA+55vtJj7L
X15vLspjGWeJF1yGNo66M2QSEGWtJP9kuyHsWZC7/FZA6JybzERwVoUFLnABFH6D58OkyB+j82eg
RhLL3RhQYCjF8EtQNWE7sW31q0EbBn++PIzffhL0HYjiXvojiiMjXcc8FYflq1RwQec7rl7hzRtd
gI4nfkkWmCEzA8Ln3LfEpmdKDWJo+CPMCRtQJyGh8hOXKXVL8znJ95pmFqJ555QwgKAAPQFtKDco
u1OrPa6sPSaSCrkowHUJUyGFTl78omER0FA/mp7PcmLJ4hO9BoNhyZqeFMdq5KmwOH6Fwais1JRw
3VBukGjNVpcpTxPJANcnnuN04qPGcqpPPCK+hDR3iFfHs0ZG4Z1ZyeVVYE+GL0gCW1BLd+1+Xc6b
8zlSgJMiGpXEtL9XWJF/XtS+OdLU3Zor3rgwpD5Ekgbw6zTalDyzO33CapZU1t9EIFS4/T1lsNsI
iYiDHrr9OC7U1oxHfqyo+ikO0crJWschd3Pb22xSSoaoolE277wjSf9QuRXg7Et3d5p+S779mCH+
0HzxekHXNYXDSxsnFj0+DxdJBT1nH/ZUqEpbvM4kjVNZkPxOH0+RaL4mz5k42XKyApNK7IzgI7NN
jLw28hxAFKGo0L8y/croy17alqQe8MpJIWcdkXUcQ4CSdmXbdhuUUZeuzQXfOlMOeEhQ2/nXd/JS
VDPj3quNC6IUepTJw2AnCpJBJ9HCdHGTOgjDspgtyXN0kmtJXMk75Sa6VerZto8sVYJKO5YDtZ84
z9dmZCJWHQMLbh2TNeWTnbMRwofoNHsZ1aqOCyrBdo3qloMSALNG8lIAALx2qxTEp5k3YSkb9Rbq
oviYWSI4zwmiZTIPJl0ZhYGEllUHcDM+4PAy1LTZedNwZ/BipA13lVE0dPTkNjDEm6rAY2onydsM
baRUq2NrV+QdJ7+AqytlXDCZWUYuaAJTwwy/lvdx3ytHfHL0ZOCdQUJ0E4axORQvKFR4WzmmsBuS
Zo7nC6iwpRxRT/iFfyqFoj+WCp22+Wlctsiq1at7+8z7/udlB26/lOQO5lJlc0x9VFxJ1dsS2boS
bDBNOm1P/NjeCsoq7D4bh5eaArY42NlbqnvyxMEo/HUncF2DJ7Hk1xUcMwawckgsEbYT+GPDTFxf
MlRPPMneHtF5IlfKFPT4uJDIhe2NUno5/+d+FlFicRY9dE/uUpOLqJZPQYZ3Z5COYTuRn5jLjpuF
H7/7PgFKynpcLkaGlCMpDT521U+FMsgVbm/Z7CHTNaJmf1FGC81LKGHiqWXdo3FQIPqE/vxUogwg
V4sMqX3kDiZdWudKR3veSUEjl0KF5NTmoPU+dhUM2AEdQ5fJlnx8vQ9VQHp9f+KcnJ71bjx9ychP
mVhnvK1qOQpxB71YEnQg7v7FRyDBpleNhnoaQixNLRG5ipKvYfq87YnH2rcUG9HDO+ZO+AZfeKUU
zdhXtkyHZ1HZTEgxTf9wwQoJCfCUbB+WBREauFN7wwYrXgfqEAi9CHkARJBd+IKQntrmTg7Wa/up
bhGrVJcrFPlIiRsNJCFasZydlUz6hxarKwSy0bwfaPR5g1czd+YMgTcr85Z0Ba6KvtGvtdNTe9Lb
O7W0dSSVOMISGJG2ifM9T8Xwti+x4Fg9xiP78QQ2SaUQaSQ+yW9R8HTEaJ7QIP1P9tcxh0OBnwkJ
VmFjeR9EjRs/TiyNcNK3OtbSNdMByyQZe17oxQ6ym96P2CzL30kOi71RMT4bntg9hMH+Fno4JgiR
HN0Uk5gEF8GP4BrL2mr5VrnLPwJHvXMu5o2R5AjScjoKZWjXdv9to88jCyyBNvXWYDuc/hRVenHr
4mabQrAWpTgjILu5oD7mw9kiqp2Qx95KX/2N1xpw1pkPWUgLbXukX0Ej1oKN/cJnfNPsjUyzTlxW
8uEKFNL9slQaKFH3oLA7b9B4ig4SKj1H7niWQiKtDW7SLoTycuubX+yaZ0jrtG83g5Wbi0T5JNYB
b6WcpIOh8waM4i4LbnS0TDt2i74tMWbGrRYRebDWT/M2/lw4DNfuoebvp/bJqwmCLKmFVJO2MJjG
hM4BPA/Y64NYaBQ47IpNPbiWjENIm89L4Bs8+yMhkRSDyBakm9jJtNeo5+6Ju/r+HIjHnf4OYCAE
KitoDnHII/WHGdP1KqTJbBGWY4uLZIBzkO32IdPQ0toj55Hxlzn9sFTYfMgjoon8KsH2Pc+FXixM
BnX3Dt6M8UPaV7Q7wnC76EcHY4dgT3SPxHCmm3rt5WG9j2OVpd65UcGZoiiyM+4sr4SrT+v4Uuk4
BiX9O+8Ycf8BnWu82rIYEomSJSPHFV9fJramYUJDNCsEQV/fNE7GwXDCpRDpCdF2CZAXHNnH+mCw
5zpH9dOBTqYTZOH5dbwyRgCd6lchuQHpB5qSRzebv1YIJOPIyURwj4ptVpBfQA2490uu3ll6OKcg
xFl3kV1d6GhHfniI6kW1qvMe+cab7DqjOuuRt8muU7e2qgTVJqsIzXNHO2TpO6ykaQiFga+H/+d5
dH/m7CL6BssaENsAL1T7R/75KQ2A8rVjU3HpzXAkBLVnWfzCSQgGfnaBBQyTL/iygejLOtMTuljp
CW1eNk+N2vviO2urz7oWBfm1HNcgozwk0M3rGbMRF2nVZOv7ficV15a+ihmxjil+u+ZPqg2uVYyP
2IcQdRDC9TJi2bwEWe630NXcxpJsmdQ8YDXjzJuwB2sGR3aSwAe1I6lMao6ss8I9ALal5qK6OnzI
7CQtdKx7+glwoTW69KRRdyrqRqaai3VxqPYNm8X3iYcrZNiUr778OWormkQV7OY4yl0NJrFRChHk
9o8fwhKHBqpJv8Sh1pGqMibG1jiJlH7fRdhfbcEPfAdlgoN9ITk9YSAKK7kjMstLAf9voN34gGE5
bRBlbP7cxCaeb51hYFKN7xZUS3Qoev9ZBN+dSxlyUbupSwFZ4LHy/U2J0ueTm7l3J5JUtob6w4Ic
oDWJ245NL68b/bwi5/5JR6faruoXrgMvjYSf1VXDsEk1LvEoMC3p0NfwKq0LugIEprqF+HjOx710
JibYk+0+9EO6lGqddvuxsgyObvXBg/ww9JXH3g72OwgZWVPdCRenQUjDh9vvFqRhDtvEXs3RKUN8
Vx1ORcB1hgibb2eaHjTp6rzy3LuLN5ymynT9um2H8yAssXBbYxU8GzNDTbGghYUJaVFARZsAFAxo
FlD05w1+fXTChDUyiDpDynNkLpQ0P2aS0ZMXOa3UEebCfDe5eFzuIDkZyWhEYwwVdr45DdOPIshN
qtRjks3pvo2C2kKGVLjwZfMwDTyfF2FIPpYT+Nrz2ZsM0WvYCfZZPt4F4XYlf8C8OHWtc8dooPzq
gvXrkkd2xmk0HPefP+FoegOIN2jbtrZ1gUC4M4JN4TtreLn/SYJaD9q540vUVryj0Imv1F8m7+v6
6uvw8cNypvgASNcqfX5BjWy0+Y+4zZT/qbu3I1s0rlzh32Rqq3x5ppXjV4LJY3Bd6PiO55sQ6yQB
T8Q6yhauOmQFctU5ITlc/pRgb3mf1SAaFgtnLXCOyX+iW+tuWzsphokf6NLO2Xr+Sq9PEVp6jJS0
4HfuzEq2Y1kwhH8ki+V+Rn0zYsEyC9lJl7W6dKSaejpvJlNGkDcfNbHa7P6kVc0HP8Swx+KNyVNy
ZGM03tthPwEAU+buTsKjp82jHXRj+X8j6IpqRnRllbp4aDmqYUsA0RI/Xcjv2QfWjSU6XQ0mJLkp
TtaebfjManEfHImUXrrFnaANn74hobn2Dy3s5vZR+oo3SqWSa7GwerfY6ZtvazAcDt7SKGccSgPz
oFqLqyn4xVSbPxS6IUEUIrZtm1xqkZZSalzVJ8yyMPzqcbcSgfWJ+kbiPTWvpI5NWbOuYO5CVr+V
pzKzNKb+xXBnwgzeVZEj/rNOGXEzlQJh9gj8tI/sXBo0LSqM8zMnLgBfr3cJvBZM28Pk3NFq0bJ6
uSkVpBht0S29eJXsuPN2FZo0yaMaWY+/GH71ea3BTTmfoFMpxQULeAz2mIjXOLUNADNW/55uk+Ir
L47ARZGaCsQmK1vbYfG5POIYlUhU83VlJOptemuDCeDGyRNaCoa+nEeiMizeaSaoVwdSTLhEEZSz
HrdWuoKFToSLqaS1Mvk2gjscqk/fcNOy07O6Q0ajz4eqfMRpgf/I9Wu+8stzT5yCJjEnEWS3JJSe
8MAdrGmbwO/jC1g0HU6ovv8gqZeJ2agDcGPJOgABDVLmObEgsvH/3ZqUwzejnb8CVD/+15Ushq/m
6UUP2ScIzdJal9SldHi2pjv6yIc6fuFJos3i8fFCB5hWY02+B+0Ctz+tFiiyOmg26S/Ea67e2CDf
kNxQX3TLZtvR/L9+WTbyrI9XjzuFl5KOYWfg55axu84IZ9lWWJWnDouyLiuvR70IqzIdM4HvXA8a
M2AAgdCBRQs+Vr3gavpEmPLFbW2x5tZBmxoPMctR1Ga9bwNJfTMVCEBUT2M/ZeqhYYFRhn8v3LoP
brDSzl6D0cxA0e+JtPTrwyINgjKx9vhO8y3PEE1VJmSxwRcNNQ8lDS9xtcZM+MQW2MYmmmgSBDUM
M1umGCIJxIKggJdkUWPtpGssFKD9S3TasstBYCOJirIVKeoXgPx5LCEV24ltTPo0au7K67XBDSgj
mGid/0+U/AALgPUmsTRJTvO1r70uIQaYz9YCwsZ0hQz4PZWc+6UL2f6RfSupZ9ANmFEjejhYf3KS
hlpeHQlM2LDXyUFvfI1D48UwDxM59kqsd5l9oUluVUy/YEzF/ZDc3zlUwfnMDkuv9iOixN/eiR39
la7Qhs7w4HOs378YqwzrfZd41jOgWdVg8S9cnBs174dZYfiTCZpip0gXn9JVQaXm30t5k4LHhx8a
Gug0FsqB8HcM3Kutbf1hyoDmGNr/rmUgtXZG8DEv1dz9N7amBz4lofVWHtLPS+xya6jQRqdLlArR
bHQ880XKLjnKenp8snibFyGt+dR93O52y2pVkv7takXdl8Ub+pe7MiR33ynca6JkzrtoPcJ99C2X
euDqgbX6u0hrPQgpyF+eaTPA3Nbni3jEvimTLPCUh1iPl06kTwubQcvFYv2jXeHDFUTCB4FriXQA
Yo363nV/9E5OynwRrbTpLAfL9Z1la8GiypAf7ocSxtkLLH0USjkUVxC/JzuidCUQSPbAk5mJbVe8
v7mK3xArys5nM8SpduHX1Fjr3SFQWonSsGvTgg0laq3v7ihv6AofTjJZ07RB8ZpjZCG4jH28wSSW
1aqeXx5MDx0EtR6mFkfeY+Vw1JwIEREGDV8ca5m4IfAHMI9xeCG5SHdijMP6SRrQlUsF/plK/1tl
rIzKaEtpYPznfIdqnUx+M618ISsc0KSK0rbaQmkrUQic4YiJCv6ktV/XIQ0yjUR0iOSIrZUQ6Qra
vMYp5Kb5h7Gzeat1fxFhDCmPXpkqQQP4fgOH5hYU3lXImo7gSbRYGBCQ/YF4BXNHH0p4y8EACQGF
QwdnoTQNf8HR7oIeOCbS7ryDin9V6tBrJ1b60Rf8RkfxJjiTzOBrbB0XE/c0rPWg+3rLrq+A9gZ9
ZEHHs8AliqT/CGMZPeYiYHOydzRR7OICKeR3IptIxjttjBje2XPEDTxvd4QIjHzLom3421fPQVyN
gGky+nrY4B0/2XyHpND1AOyxZ37qeTF0i4+HzC/OesTXpPmHwzHSnbyUXSKr6rCvsTg5Ofxuhkc9
YV7DmaJGeI9Ki3FBZC213qjq9HeOHPKXEBNHDGEdaQJkGtRq7ylmE6XmSW/RiviVckCfRCCxqsF0
yX92dgurGXSw0QkuMQpaNSNVCkyUffb1Ay/KhKGwX2LmQpciO19HhZIT18qcMpPskUGqJrznLIo0
2D9TfZQmInPMEzA830hmO56DrqY+cjDf+wPjQr57IM0m1jWrcciUXq/VPjFiufv963RxVf4hti/A
Mh/M0tGLdAZlHO0wD9bXv5D+NlJGfRji9VmAA3NTT5p+XdkBIz1hgWfO8GZuridH+Y3yuh7K1nKh
tIjrIxSGl2Ka99REjezF1qJgCFBnjZ3qqxurlXNNp/sb2y514xmRIufZT4iZc3aVTCqVUgNFFQNC
qy/NTIj82aPN9tmZhIhpMtFiZdHs3mBwSYatqDRnxkVZE7zdRQL9+ZU8NzQe4wW16lMA99CsS2bs
gjcAYTuE9gO6TfPefvdwtf3NLboPlJlJOVZc8MeHUj2d8o4yTbUnARsE2Qks9l1L/HF1b+sZff75
ZB5xhdL3QpkLPCsQpmNGETa3Cz4OqsBVR48vLA4+P4G5w9+0yXJvnfjkEgAS1BPt0bIKTKe5z/PF
V9i1opeLUAQO6bsx9frGVNzF925Kd7fHJk47Bbd8jurxae8ZdEniFnQKeoeid+eywB8L8LdSzF9q
FU56GdZlPey5FOEP/mGnbhiIbf6B3c8fArrqmuH5JyfQPUBS1QQI/fr+9w8DVW3z7Gjlc9bQT1Uj
mMF5cAd907+z7vPJr08HkQPl5c5VVEiGmEJJflaR7pF1Ezi5+KWaxxCTIaim5KfCDb0GXg2pGXFH
dDiof1eg616l2a57pxykkhxwq96YwV0fM1fldDqrzf6PNulGTz8sZjINaJFY+11PT+u7q6aOVd7L
OBz1EMnlKuvhexYH3N2KoHzT3fYvks6F7bPEzBiDN2tBvAlozBpubmyUhxwdXkSK/bu4oB6+Qc2d
JgRQTeMv5Xe/R0NWp2TJejnYC/2UQ+JQS/YSYT2mk0hHwG3GbH2jH9+H74o7f+Vbu//RrxM4e1fY
fYru6Umex1HRW00EPOvsT9UivOwJQV84gjI6kcj57/k5oZLgjxOupPNPVPnfeCfnGeZpE7zBMVZ4
eZH07eIv4i+54W9k1w6IVaKWSMZGw0mbJQC2UAmFoiH+aM1M3AfZGuAn8PeyHcWcQ9jNL4UJrDYR
J5U7YMCrW6tEQ0dH3JPtijYIxOlxE52XEqDVT1k0g1ZwED5PsxVt+8eRFpKLzvSvKJdORgjB1+Lh
xbSBWx0RgjS+MZykH6S0wHlzHndPvDr9AtayN/zq01gu+7iQvMid1OLlYBZeH0xQEEKVmk5kpQkQ
3N9TPzc8ed8H38ufgUM/edJAv0mHALYp1P4wrD72I8RSwswCJQts7iElGia378epgPy5RilBB8ef
W7AC1PDJ4Dh47cXVjw4W09zZRu++hx+4XBMN2Q+INhPoqdYHEWqHQOsZx6RuvO20ZkmaNWJxXRJV
tTqn6GWDZ++Ra4YZYrcaVJjga233Z8Q+AHvtOpRHfs67NAPV/7xfCW0Xu9/CqTXqNvUA3iGFgBNg
1yT8SWO7lYqKvl0rEZTFRn5UowU/P2SPqcsFRmY7WlUMTYWOfIuU39D80eEn1nH6WsRldAK1/zvB
+adPt0Fw42tD5rgHt3+HdEqJYTmZsgBCRgCDZLx1v13c6Mqp3VtRmhsRklwHYwo4JX/sGGQ9yaw7
15wveYwOG4x+5FB1KabYrAZY8pbKuSRnwh+4DLg8Nn55AcAotunL4pmDCSIbAuA2rNFBW0rMyu7+
Jq8IMNLLzD8/Wq/5hMZv9Ax7nDc4H6E6tibAFjycTud2Zfglh+xY32/iLgIxeB7kyYQIpZNg1jM3
QDujtT7q667aYqTcSClqKN5KVDLVOxECZZ8r2+/CjWabCv0du80eBQNy5Slz9HNXpooVRhG5zBS3
yh711+y/xXeW5WoBvLGjcdUQBcSzG0GsP2jj0wuNKELmREEJfzXaxcUYOZQCej6FieiAg+LFZQpf
K6Mt+kYykekIMw9RtP0w93Y+Uvl7YpENTJrf8VznMc4ysnKzlU4qi7crXW6pfmYBrkAtswm3lWzD
bPKCPGzUb7plcopPLjGRjKpHcLWWaDJ6hRU22mzMYUeABRm4Y+BGzOzR8f9Wb4Q3+6BSqdiQ277E
3lyP/cwC0n4Og75pQq5zwvkU4co9YlWyrQXdm8rQuyU3aF9OsDo+KDZwzfhWJTk3Ht7VqHM2OvP+
qRwIFZLpwdsWwswr+PT/6RQ7KtmXKkITrSuq01I0b9/GKQwPOuLOT90v842GidhAXSV11NlDoDAF
vAFt0S1MiiKnKpdG5oh0iZlZLKdNUqD/s76X1CV98XjrqobgI706Ogqb50FEZUb6QxNxHmF+EWru
kD/Tyh6FeI82l9PksRWtesVESRgcREh2gRYqqZCtfrJPTV+1rwH8eQ+BTbi4YhZFis0A7AGOY8Oj
LF6w1u8jZ81cHevLeOgOrwQTCv/9iccsksdtfNGm47zfv+aMeizikDemgXPUJ0DfnopKbxvUz7G6
YSd6lFRO6DRJBHQbTZ97l9w51emEQi+5ii7ULu6rp9UgcPlMLboeuL4qX935h2rxCYfU85qvrrQe
qj6Iarjm4tnt4oGqIo8eYsxpd+LcfLAQzaGdEqHf6jMHP049eyWNLUwgCiDeeVdgbHhnqSqapa5d
wz6gqhi2V6hpoLMdjXiW3V8h5lBKntDNwL4mNBoAtCi1gHNEdmKIshsANJicNh82VzyqB0nAMBb0
1H153TDOgY/TxdG4LqHyDNYLLVMKPomFH1mBK/fzXrzU9KFhn12afag/abhd3TsJDVuRJw6oQ00W
rkJZ11WgPro/4l5h2S813Bo9IgarE7mhEaHsHHQS7u1+1Ni+InevHtB0gkxfo0jDrpSKVGvbWwS4
96P3CEm87ldsAH8nBVToOVuyxwHgQVuEDoik59dMBF8zwZXIa0w7GcZMmL2vL0jorA8P0HC8LXqQ
AqNFHIWxjqDoh/YrYObvS7HYgSEAzJWiUUZQG1tY3ebgn8STaN8BRhcnavN1zMarOnn3t3b8N4IC
yg9Ube3SHLW4UZz0LcGCMw4ofveO0pg8zwpBotw35KXN30DyH//WjUsnwQFDafjHP+FBoFcI41NJ
UhtpbajTR3fJWQpZmFDfd5uQnVy0n1XN/T6Qck8Q5zCefuIKtuMl4neTIhCXn2N0HUn5ktGcEh0k
OsOjUSGVtRwuXljIZ/SLMRenIG7Xxd30bnrImvhp1wsYzNhc0CgLLW7ggz4UVBPHioN0NbCTXe+l
Eh0pIQNpYv+dXIeR6P9LW8PQXdBwWN+YmyTFQI0gi7E0LTCZKf3fWXzcOmjcY7UtAb6+faJK/LbK
zjAIysspEATrIUpk2M9wVZEzpt+sbp5Vs1coWtZYesjQwmPbpTLD6uRuZbZw/bBY3mI+4qZ9nDSu
oGmbjpnbMf3hK99HM/+kmobiXWaM/mGrbuPeLpfyoDHt8U2EN7HQBPhDD06RzjXsPmBBps6KqcDQ
0ze59qKjmnmgvNznsSVf/UnsPZ9SSRH/HvLWnyJxM7vz809GZpFCLGQvFtu5IOvUInhv88ChybMw
f1FFsiHxe4MaEtwv0bNfI/KEAAd19wCSECDP7as+JFg2kpRY4zr+59cAF2ZY5S8flKn9iOFwvqDa
lZFWZSM0xuXc1U7leEqHfOvnlX+ir2HeGCPfw20lWwTBbDY+nCdr7k+dfobSbYHNEeJFrw2myV1r
Qq04Qgi9ugs+RLO5drOtJaZOvtszffYxYCj85L/3QoTAVCWuUIEZ1SxtBI/00YqgcGeRzmNHy191
9AZ4fCzP/OUxSlgFJNWzCxZujKuUv2hikv2ZsQ90lpHA4cdGMnAeqa3x2Y92yVaQo61IwATbtB1B
X0zkTZ22y5v6L0Lk4K560DnS9u7gbGZbQK2TEhUVL0UeKOoXWh0GhQWXcAhwpJ8xLOX1IEuv8C5u
l0HOpk70LFX4ZoSsySci+3EAeWbF4AAp2bff+ZQR3uOjMyRuTlqFzH7slBXw4AISMncL6wMxZkwR
Swk7A4WtphI9Jrkunw+M97jom5+EwUyIsmCtIh4Vsx9xCuknITBDK0DzlSLoXL/Nts2AfK9DaBtf
BnQJPwOqHk7dkpVFrDYfUYCaToRML96eGXU3ZAtbp4fOQUvTUf3/Hpmd1Dj/OWXsZmxQd7KJtieD
4lMS8EfUYoVE6FvQu6MrKaMH6cpWReq9gFvrM1r9yGgwjCuTa6g794rwMTnE2LcFBjoRUOYETKIP
AxmcfSdmEQfPnIorh4CRU15zjmiCI5HpVPucXgbkHf0+2oF5sLILEjkAhBtstNlJzBc5bbPo0Xcp
7LO6gC2XSVygT9N6ViOfSwoFVsQqIAx06ZF+cKSNAWrMSlYCBz3wvk/S/aC+xKWsylflPJG5KcAg
AJd/zWMPgqM2pdVsAa1gPgkx1S0kgUvXJvjAMgDqm9eKSKyK3ovN6rj+0cJTG5/Gy4/MaKzz6xXU
5vNrJes8O+zN9cB8ccsEiJostX2Q/1KNC5uJRarjCifXrxiHD6onrIpiP/I32bpznpvSPRkPBbl1
BDa606dSjFzodVpFJ+uXWJk8rYa/Jbz5bZVREDnSrHO4PWq+S2v84hPNqtVVv5dEeFuccVWMLtH7
6+MvFdBmbIN+yEOSNGRqpiI3Gd7zy9uMoWrunfUQvQMABwy9c0/qOKr/12+SANxouKe6eKNEbj+4
tNn82peEBDbVTpOr6VLdjnvLzarcAYUAeYWMJhEPJ/6fD9I5s6md2h8zI2DJs5HRgrTqc4Zy/MtR
LPEvMzPyCt6xqrF3tUc7b/pFIGBzwJ1B4scfaQBkIAiderxzNq1gs5gB/XzJ3+vWblKoai33POK7
qfhuPBxh6tQNDXMIAiI2hVvSjGAi0/LVpmGxm6Rxnfji44c3iF6fZkPEnxSHo4LY7IAas+WPhaUt
xKljCAQso/bhrtv7ZIOobjyrFepINvjovfJjZY0Y1uXF9qd5j36AprCRYT1OVPa1TDH7NFMDrY2S
F2eydeFyiiJt4wsmLlNPIZYCB1UvpOrvSFqfR4Y14rvZfkIPskEe5ge8O86UhlcsAbhJHT9RS8hE
om6mjzuuQU6HbW6pZsWUFhpzgfoAfuD01P22t5n6Vo9tMBrQFAYW/7CliKAGN+kDLmV3bn0ydOij
xSDvKm462SqxbifwgmZUe+zDJiIqpto8gFHvpV0mGRjDeH5eqjQpq7aAlBrMDTxnbLSWoGv7/KoK
mUv8MOBwZFK7LZBV5TDaeSUSiSZyLKJ/vG1/pTReKvAgW+2/lmNsWiAAje3A0icB//TV1dWgqo7a
GvZBHpmKjTQqlCeBLXQJZmBPkk+pkqkEer8SHCBe2XptSBYXgBAzH9ODGHdMswR96DHF1qfhpSKk
ejsWalKgWgUX96ns5NP0rfGbMNrZaqZbHcKXpWEn4Ebw4mfyl/Ah3Ffc20nnYnoUAbIRn3+cLp8/
cWDRI1PQOzVLWwUv0ZaNpclS70olNrDEvLl/hpKfgUMWUZRP7rgWx3lC8ZCWILAb6F/3uT2dOU8Z
RXOpZydDx4nB4Kkt9kdbDzRi2NNJ8IdbWoth7J7uHJjA8vCvlh060V0wwhd8CLhuChhpYpq/cRUY
Hs2K+6uq8MAAq7XqdMW4rUQBYMN7cbojxpa6koo4WxIcmDxMy6OMjQYgRyfDQNa0E0k6VPPx7e96
L0onxaqQxLi5PkgixU19TdQQPwE+qxmwwUGDJgShrOA+5wwg/zmL1vevuK2doHqApuEqNq6DwGhI
tSTFg23G+JRH6Youwp2CPUhEZq1bai9VvsWlbm/OmgzQaBQT4HSDrbxFzSifmTIbIi2CrjXIgquy
DU7xTp5Z5JzkMubttDun46wRxFlNw43S8lh5MmIh6Mk3M0L2YZYHrSokjxV1sk1aygtlrGOTSnlk
wcd+E9otvLacY9RYGWMkpvou9H5YsJSF7Do21tYaWc0sOWhKWl2rLYklUO78xu+ic4SCSVvVLpev
8TBQ2YrVHSThfXtaZtYQc/rWR2REhoGh/0l4xNeYyq3SePdWEHbxsZP7Nhy8HkhB9L9qIzrW25cc
wJ6JS+Ofy0BR/P/DZyQ5hh4lC9g+GxKX2pmFoJXMOP0r5JZwjHqw4/48tRb8UwV2wneBAuMyvdwl
OmpSkDRFZtR1lYyv3TM1mTLthJarxBsq1swmo20KBEqQTzXrYLDg7eSP9qx8CuHjDZmPeriNwcih
9TlBEL0SGt60XmSTMCAUGiUeLvLbtAiiPIa3gYSYtZG1YZfP/gJQ4sCvNfrWXBc4dcVMdF17hL6H
dugb3jd5Rk+nLdLmJUWMbK4TmKHw09LHR2cn318LcKxB9WLEMUK8SXnqyrqzJTt39gT+x03rXUZq
r6LdHhPtsJ2Y37ubit12STOGYOiazU5YIWfQ4xVpx3Av3ALYV+D1N3rCnW5zP1dg5pxcvBLatREi
8qYRtA1iGhdltEo1cChb9CPYGe5hsT/4w2zFOScfUh7SffgJ4A5QRSHB5md9D9W3caAklgu0g425
GZ5c0ef6pKZ16JhHT1KhDhehNchpb27a/HyWaiEJ5yihObeXfZooL0K4bcOBiIPtast+DhJDFhL3
ReiIMENvzqXMqbQq8mjsgokM/qykYkb+KuOOdSXpVBdzGETok8aAHFGc3pFim7TL1Sr1YR9jJYE7
JsMAt5RqVcFFCnJjbPbNL2Dl2xfEw7NtVGjsn367MfCV/k+jTD/eN+pqPC+W5BtppIZ3LK5XkGpD
6us8/6pek/2YnKXw7qeB6TML9LThy7tt0NCDf876FY3d9dcuDqcAISaGO3OjLBEs0wLwcpfZLVxV
hCTTnVub2mEHY8u88iY4j2NF47XClA1PCFrGCpARfIOcOFGpIP1NrtYwpPhlU7t8Hh2D6Kw+pRpd
RB00s8EdfAUTu/IXPcaPlALkh6aVxngUoKg1qQ2UwMvgoLA4fgURyLRx/JvbSsIfm1pbaEACfslQ
TmrDTp7FuDd5WmYphwB23FCLmEbYNOR/BKhOI6SXUyt9uuLQ1NXvNlx/XUaI83vInSwXdyZ7RSVU
e5I1RShwooVNSu9x88zE/WL70J3bjSziEam8cjI+Smme6HQrAYl/KW0z4ZZQQNsSdpBNSp76MH1c
kciCmaL4Ze1HLAWSeTfot5zdL4wtAB7Bomt8OgF8g3EbyPKw5lkOadrBOgkLpxQYavevMGPH394u
r64TeZsz2JAUMaSNxsBtzwy33o1XvKnKYpFFM98q8cwN54j8Z5Jhrxxntr57HjTDfxzdWbNKKGI1
3NgccAK0AKVyGaZeLkwiuTWUj7YmQ+jn8MgpGD2G9/IUPhjaseHmdbI2okY1dUI0lU+QCXCnLHqj
7Lcbf8Exu8QqZ6HbH+QHKemxrFwP2A43FtBB1tcQOO0z1ZYAUrV9WaqFnIoN2r3vL9VOdB2//4+b
IBAQ7CodT/U7vTomWALWUdW6WhDdHHsHVQT7H4c6PZ6/9KJSA2WYPycq4AQlUDvRURrylh46TX/p
9q1wxRnUBRUXmik1Q1KffLkL6eyTbjKywMjA/KszmHAjPxpSrLfdKrFU8i26aIMwz6Z/9UxULAVi
ADu17FHVw1A1qIN5HyI56QzCt4ujEq08jxEQfHhQa6Iw/+CSdKRbSqSQFywLYh7GFwNsEcVFOVC6
KttxY2YT/54635JvxaSiraaGIVQTd+JNJCMKR3UHNFYF05qJiH0aFjaQg2mLNTCDKymXYKzRnXGo
Mwn6g/Ronk+wypOBtD8ktvmOwxMd3anZfoIgAZoBCeNb6irtdLEHWHd6p9aPIVQ5LiqCOkPSxMOD
oFVApylYOvRg9mJzKcGphxngtdnMUhLJpAIxcopilZ5Itw6vxtPklsm7+8M9suF7JJeLtM0g4LKW
pLySOqod2B7h8p8GMOjEOtMPU9GbFtWspImq1a6ttHQKus3KPhsPbysSB1txXXbXcSCxrT5iI0gH
66BGGHKIqiffbR5pgAnBmsVo4ZjGMf92i4FQEvU+FCpHTZJw6fih9jQxgA0Oz6kpHJBNv6BorU/u
dQKj3Cir58H8kn3YzFfjcgb/Z6Va7tW7nEr1hEyYx1PDmwU62ioxQ3MsClPzhzFdXkfMeDzGaEuu
2iYmgvG/Zl2Oa70M2RlH8yfTbv0b6AWSc04oLCcz77cSOhRqyi/gkgT98NxjSeuL7S+E3F+QG5V6
LjIZtInCcVH8YcfQbIwcMXTY8UQBsbh1irl71+Jy55gCJ8kzxfXLH7qpyLRuNxbH/S+WfJW1w5+u
AF1IkbtSfOTxJAn8rt80FMA4YWBEfYj9R8X/wM1UjLMJNERBF54sxlwuYN7B0CQpbFVX2++57CTd
bE3yv+Qi1HcRSgtVgnrsnSxQxYmysmu0sWcCDB6W6vWL+XcNQSu5MgGFsJj3E2aaB+jSV4v63nMl
dare8eAdkACJ+WXEUh1UCqIjhEzIQOGkCvR81gYMnF3iLiLAVcqa07Fx6YO0/vPmveIm3+V5KBDm
njm01LU466PQQRIFXWERcm8NAUdht5W2Zr4HMYpvB9IjQbvyJeypGvHcqKbpc8Bb4lkKdZlDbZio
Ga1Gy+gePY2hHKkxDc+c5t38BauuZwENTf43mXyLyO4U+59H0IQQxaIaKZ7OU0OGoq2Fyn9EWqqj
zmSNzGNftEhGCkNqBJg1QLdoc0o/5UvUn3RzlmkJmNiZv0DQdstYp46jtR5gBmJ0/GjqGu4J+H3W
7zYtCS09vQX38dBOFqv1ZW7iiuUIehEHsapHlTL5rdAdKgYHAr6LlyRbySnl5ZOCPnbjnNQccNng
P8rsGqzI/AeYZi3/PBFcIGQGRXv0M4fx7rLQHKQ7fMLZArX/Sw9rRUQ7cUsvNtjXttpHNPEnAX6A
L5b+U2pPbCQZ1m8l7C1p9wDxxCMminmESgmibGU5iQkd36aZDhtbPE+Kd7dceYieRdKeNVafT9eA
RPrM95hhbSAWpYLy82cd//awbWV432VGlIOCT0JPU2PVxL6t6/FFT7CQDwCjVG0epRsF756oc74B
OJiMUkjcekoh0VtP8bsAcSDzE/l/aPUDTezrOvScq6RxvmiKyW4CmAhIUuLqkWhEg/FXR23bJk8F
9FXmvcQZRw9JCSUnP3YLXX3Fj7ADE1sqT5EDQRJ/IyD7Kh4tAGOEDNa8XaxR8My8QWn7kuC2l4KX
c30LByw6jOF9KX+EDPacuPUUUhsEKIzI9kaA5kRz/tVzx4+FRoEujppKgn05lw/JREH/1LPWRoJS
YRNfiyBGGXcnpztS/r6B+kRjjt/JCiGm1U/URjPb9gLIXh3iUVGFL5bWQZXKkbuiNEOiKKfIyh7n
tXI4kZXRaREglBEOp2Kmy1Dhs1MDdMiWG0fTJ2W6RQDX9bInCnes09vqmBCTrhxi9lQePlhNenyS
T9d9IT6DNLgrzqxDu2McBgQ+6QifSu9RoijRenLgDin3Yi12juByX0Hy5bEkUJhCtl8Akd4a6mGM
Khtx7H+hO45ETBpYMEgtexFvBpJFtFU76So9lOnmmAYeb76ENft+U4qODnCqmNhKNhi04BNVs0wh
bVAzOHIeFBRY7PWMJ81TjCgABkfjP1kd4I9ZBPoG6tobRH/r0bCoJARMIEX0o/kSO2aB9UIIlht0
P/fmZS5PzSVeAvfsMxET3GAGW5mwSgr/Tmzaw27DE8tP4gH7xVeMzCvPblyKaojawCUFVdenkEbB
CiAWHOk280MIKguyxWZrZ/dGT8gdnlWVsBLXIp6SMvnTM+I/UpO61eTOKdAg88vHMr5URvY8p7hx
FaNfkg4GnMD3JRIwgkcY61yYQwLuYQxbat7LEk7zPnSiJ7r0dp+sP+xjFI+nFDnm4C04BidUP6Gx
HrMrvNuXQTmyMH7eMDdfORYLFD+E5RNqTFOj6Xs5Sta8LBHQu+RE560qALIPYb/OEJrsLQ848PM7
q96RkBBCzv1uRGaFj1ZZzwtuUp0VRDRkwZJ+Psv54K3g5NwzthziX6W4y70j+aWnOQCUiALi5HhF
VI/D+4FDkWB5eb3RZbwbdSG6M/vI2ESp0gBtqdHcuGRV9o9YvVFDxajXwzbOOxLKUhQ6+kP/IIsU
C4Ujkri6Oj6mSrRMUmtKYAoK6ycAw6E4MGFTG8tFYg96+2NM6tGxozHoWP8CeF6jwncsp1nRlUDD
2L6xoeZnID7CxkGwGr2Yj6ZWM83Pm1d/+9jlW8nwZDXrUr17Eo1a2DLjWhJA3fP7zNMkYyzok78y
5SsxlaxxzqQ5nQuo7qOlJG3Lk49C86/D+ET7RU5ta3pMLsGfzoLVs/oK/sY+H8fxytzbA7TeE8oz
CGEr3+i+BWuViQdHc7ACMDdgQgM35rrTU3wDOsepcBRitRNK3bNcWUGBKoBrIFJkwh189XS4W0Wk
/5U4aIcj5qN0Ieh3+fLWRtPEle/NSogZN+lrdGvS7EqNCPJYagCPMQtl+RQguH8GBZl9Ea0Yk8n9
4yxOteRwUU4Rp18Hb4LAXAu79WcmnnBSoIHKAUMhkxUmh8xTZjxrPv4UYr5R749zi+IONK5O/BLs
ov+seNhW7hcoeo+KCzI2sltU7RM67gVWOB5Gv3yQQo9k2WJVos2accVKYCzRSI+6LPmOEF9XilJJ
+Rb6Gxr1EtrhqphatxV2WcFc/HhaNoUWdkiIXm3AfZ0MzDJVjfYsue6801S0HTaBZqoLXOrMaW/O
1JUPN/x4L5L+csllXIK/gFXbvI/wc2jEqBl/5p1ne/mLcBjFqqSR/4c0gFLnpMPpEvLzqxA2dHdQ
DDCeZ0oeyl24TeqR3r4RG/aL6LD9puSseJMhr8TbggqeVOZkSWKnFdWz5sPMbTI8IfxCMjmb8OJn
Fv+xmL4Qm6tq+s2HEw1lyo7DqvJVEdpjirYQc0aTBWZ0dPZPKKqSRa9azXdetQ1unka+xrcAXnFb
XsoGdMx0saP2i52S1tY6AvvTl/OLrbd2sRY/B9jN7KuALf+1OQ1rEI603NatoKY+ofC/QBWKvPIM
LtkwHajHhmGiWxhNL07hUjUuA8d/GVnqJ6n9n5TBvBoqsWvMueDQukLNpvFHGM+SYVr08w7W4I0u
PKyoi+h2jt2fu/Md7SRftqc7kWYzowkVVidjBf+utIrym/WLvRp/T9EY1O44VFF3mcyfOB0C7lT6
QRgobZgthCi4VVo59etPmAYdGA+Eb9xxpG9dxET9gVBVIvhwAJ/0KUNaaX1QU+pMyZEd5mw3rVa1
JVoX9kzQ/66N8u0wQR8s3sTpLF5ZVbtmOYqnQJXkp3aNuvgMEU0fliqVu3M/1HxzEwKJ7CUw5qM5
PvXt+mRSf1iGngY2gxglr0nzm+dyGin47AvSrYmYB75LwTRWbA0rZqPWrj5e7I1VqlxCb8e770iE
uW9y4jcObdj28yVhb0nIngfnkZrpjTWVjWpCnvumL9Guc9fcSlx8G53t1rjgs38OO9d2zLqIk8qz
JErPVVgyq3iH+pBR8QYXBnxwj8rAQvf9qV8BfYzUj4eOjL1MUevZCIr+jp9TEhUkA4YDkhnXvef9
FQXnrjiQfQwfHrBsMhE3UvDEXx7W4yOCJuLmjNShnl9IcZ/MyyxUyXkag37lLsYVpUFjepRyAwjY
ZLyYEF2EKEhMJuCL0tRxjQi8bJnchhBP6e/TgdnOh+3A/L+DZT0gdfG55ox78m66D58c4VY+8Uwa
CH/HFuoYEHG3w2nS45cyIK2U5Q+6bi5fZB2drHX0jC3/BUwheyhOGN6QfpSiRXGMQqMeoFcox5j0
cBZrVZp2M9vdyxDUnHMmbB50Hazzz+WKnMWW47aQLqoUs98Qpv32+8c3zXZHNu8ukJRQDzMB5BpG
BJycsbmGdOow8p1S3ohng0Ks3wIaND/zjTbqwKWtxfkzsafX6M6DpGwak2xXxVXEtFdnRmO4NgCM
63kV8sVsG52kRaf13iCan0PAXZll2mWjHej4Kxb7KNlNCdhnuLjQc5pPgcXdGdbOcfKLEgzJwkso
92tKur7cUP3u4bM5BFlEAjQQ3EW6XlcqCigyq5WQQ1iADwDxhhkSzT87gH5R7EAzTJdiXzL8yQX4
JIpPHVHjFV84gU18aCcqwt3u2v6FnjsntURMKuHS9hGDUJ59y+qEisf3YYT9oXwV2zayPNJ0sMoR
nDG3KZFMUFJ1RKUg4L4WcxPiOswTDjFyP4Pj9D8wHVx3grFe+JOyv76Y8J8fNd9Q/aQsNQahduTS
Nv8KonS1Ry6Zb+itxW0TsglCJ2n6rnXELKHbp26npEWGuKuJIkVXHKpbj/vZwGlUzDnSU+V+YFKK
nNbT6G0Rq0W3UAp0Ev7le8lc/+FuisauTHrG5NeojCQg58Ob4upPw8SMiJ8Nw0yCa4RatzfpU5Th
x6tOv2sIr4XOGJ0kKNeGczlBgaDfU8bn18IvY2W4phIt0dNRMAcntLGvp/j3C605QXjJx8pRS3Yi
JIFTZpMD/+x1aIC9BDnxT2yeMCMvotKjRqVHow7aY4wKy2R9NKgTiDg2hcoTnJVKKvVFwNAU+SZt
kS3BOa3VkUF6M82zUcRavpYbOATgUPn38mPMgqiA4sjwXiEVZzM/IByMerKkcbKkAYWZ6BckXPbd
b3AdF0HysoxJCaK5IaVZM/JNCicqE0KmnfbwF+5JWsseHoKH6BOGU89g1UYbN575NJef1PnuXBro
SkCgeOShgfm+eRt0tOsa2cWhhQ3W+3x0qsWM0FIFZveIriT9g3uFVUkxmHLJK1PIyR96gi0yKPxY
3YBbJwo2fBfxo/DCzUxslCr8wp2m1QMOgETmE69vfVNwUmHWxRfYgRHMHN4GnTVcnPpBZeWx1hph
0qP3Xl5y819ADDgUtlV/FIkNgM7e6gVZyLulZer4kMoQfLGn8Aiwx9roTl44cwk0rc00grhnv9TN
yWdeGx1bhvHUn0sZCqwZ+QTea1p9vQu1qMoiKAex6gaJOKpeHgqSEiRiiTqOTQGnbeqFafltsI7n
O+yYRMpH7CHLqO7VzKD/3d6lsSfMzFoHvsJYQxwoUAB1NL5kurtZpL+6QmKd5VsnIQrVBmgd/2xm
EBkMaBNDHHSGDUb0xl/IfSJjibjz2lsHs7nFsc0IsttDTtKXLzWkkL2JvcP2O+Wz3bBOf2bLs7QQ
CWvs9AUFZkG+yfS09Sl+cjkRQnROyzxYOcmsK153iSE5u56N2SNuR0BzZkK24dILz42X6rYq16tH
YF/xmihaX2kYY2d+cLNKAY1WfH97TUw5EQM5IUqiFbwWlDbNmwNJsQGTJCRkONSL1ePVQNu1Am+t
AHNYUG27gvOnFoPhEO+vxqL6hFe3tE061lf+CwLcN+jYljsnYRgnPSC07Cb1VtFNvXVBkwSKEfds
vnNgfddAjxCimlRJEZVqwgmj69iNk36HNKb7gkSvzO8ySamMm7qjjbHH4nIytu6bW/IvZVVLoSnl
Zwa85rlBf9XOoGcolftoCAojamP+703pPWRXjQgwcNDWTXnlu6vPV7brunC1j3yRwKwt2TPMQyv3
oYE5W7FEGcSbULOi1z24QrjdQ7kL22biyRYC2A3bo600YZoV6Hsk/wBuskOly9eLgfVWe8hbMYNG
QDpvN3LtfU3dv28xt9IDzO/yIhVFX3UE6CKCW1NRsHSV5e/vWKT9orl6pzfF9efEVKCpzLxhVzRn
jEhiD7tOZwdm2RflZpx2Btg3K28S6/3nQT3SGXi0tQtHWnSzCJv8QrSeuxvJOdMswh4fJAgXvyF6
JNkcd5hIrprAY4ET2FAO7p2TLzCQNElNDeiL6FR7JWG09swFnjBVAtsx4d0Ane9LShZXIq0BlE9E
UAsKzuzt4iNV4NImHrRuExvYw6AA2o6rpGUdTT+YZR/S/RVA08CHahrSdgMmWFUwdLKT1Etw46O3
v0KYlOitCNHB2cr98UO2MCLzpR/fn+zJyVTjxTTVcBAG/v2rrjEOGdNzaUr+ByL9UQwDmK78yilP
RE+WQXJBdfgv1MDUpwbX7IHZbDJX8hB5RFij0gK+ORxYvytbtf/WYNj6WC8NiVTk6zk9kPYWZJIc
4k+k5BkWwxZvLbV7bDp7RndPz4++fmrXClfPGxAODHz2AkOsuci+PPbDu+A598ISz+klqwLm9Nmz
8fSgeZGgw1dl1ovo6ehmmgZgCWxULyvxA4C37xjsH+87vj0VqPALTf0gIg3eAsVkMUhg/Hzmv71A
e/po2+rm9HhkBwnTfOTJYkIJLBz1BG8THwvQJ8WIhtFWGAeQll9CM+zrAGrQZ5J3pR2sR1EgsAud
brHihAK9awu0PgVN4CuiA0ehw0OdwJGZ62hSaQsFvP5GqfwqENGHJ6OS9vuosLS91qXx+oLJ1VT6
ndq0mxLGwMnM7+KTuIO/i8XZqta9wcprnQFZDyh5N4zlTYqBUc/f7ybsyAhyLSWIKuZaxZR1Tupr
593I7CdT0BEdS5CffhWKblZDBKtZ9HohS9n/WrXg/xj/EcZTbG8BqEpGmoueIGzqUn/i2xcfDsOS
nRjJX20CDu6zfXR9tZ7yZphd3R2dxfSws6FN/n+MeYBIeEAblHjshpuTiq0sXDztKjb6H+qEOoGa
imv2z0TH8s3ljIIJY2VrdxHClrAQzfN4JFL7dODesXi+eiKAahdn4Y44xzYHOQwpWipVyUd67KQh
9HsajaraKLqLRAKn/e4goyB+xcxFGf9WmYWZUVOEEF7lpHDYmzPrZA7T6h39WvNxpGvr4hqrGkp8
ae6kLJdyQUiFiogu0aA8nvCYurJrt0+MRYNNLOLR0jmBeF7T7/IUrljs/nyaydscURJb8VHXb2hZ
4aDNG0Nxgz48CISqDYzprzJynpdM1QyBE5cn6iD3nrSH0CnMpqpSs4IVsu9Mzb3XNIB+dlV2ZeAk
GOlE2qjqz8iMOCmsjkIn6tfP7z3xKVozY5UNQSDNh/qeFE9I3E2J5Xbx4c9zNaCljuQoRxQk1kpn
yejVyG82r2HOwbjJQg1/ESdskidVhGLDD/cLEV1pKWGnxUKcmCpUSbX3FdBySnWdhnwFHys4UfFY
opWocDirq0eXBr346f9543YbSAsQSHDHLon15gaUwqmnQ9ioUMmNGjlM1LIs+W8TmbjdpUGysv3U
nXzc1fL214qhNO2MqvuJw1pWBILklAwAeF+3cz6uIN+akF7z2xO1GNR+RkQMC+/hJwmfvSDT7Vtv
kMuz8BlGQN9aSXoTvATGdh7mnbh8LaqaGg6yiNe8GnZEhZEBm+Cn283plYhMLfooV7GswQSqyaNi
12N8HiFX1xxVAVdgucKg22sKQcOEEQ/zCX07Q/y6/4JaodqnfE9ZgFg+mqk8xzGoWXXrrRwFXeNs
YE83tjq3ep4zV2CVvcfnJlW63i5H9DnNu6Ca3VtFLHv8tkkR7Kwgkq8u5nC4QEqx++enNRvEKt5S
yUGl5gESVyX3SZLOmWCh1MgezE0PNmojNV0RVAeeT6YIt1ia2lsJ3e3ER8ixrcsCJknBljOq0I0O
dylxgVEHOaG29vsHp2irJfFY6EAl4u2UqAmfjpmNTZcQkSDnG9402pnSCheOxkW2HVQnP9rFlsdo
Dm8Z3jA9qmIX32zoi1P3uN5uWQSPZqcUzPK9UHKppPnZqS6IoDzVVMdSVFvBIMptWkspP8XU+DqE
AIrlyZQt6+GczuKAOlIxPOJE7Nwh+5oK5uc/TqPPuca3U8WDVqTNBsC+eck+nZ6ayOUYzrcvWU/K
9+ih3XYYUVkaMsVjWM114Fz+Xm0CLtHPf9IcuPmXAMMhxdi2k4zJG4KRaiNMVJGWpnIKGy/aMrHx
seSEa4wXv0n0O5GAa9IdA7PNcvm26W0nCMO/UxMFRlc5ms4GldL8R6NPfka5ZXeTPBxeeY9x3sXF
oJgtLndChBjbKdcvOloTGu5m/QX/y3Q5EM2ne5jESWWLr6ZJrvgkzAqPmJV3zd55TVUQ0Op1qe2n
L9Wj5BW+ANLJQouodJZI9XSi2WrlAuNZ9UycfrHtFZmuIJH4GhHJAU7/CiXNXStv+/Wbn2BNurrJ
d78HTN5sU7SpNf05DnyXe2F1GhdCD2nLVrIGzDfaboCFE6325BHBh04tg3wXZ8KMytEVmvABZLQ9
tZlIu9Oq8LYR/mgIjLPwQCCjeBAxF2iL7prKf4NE4W0qZRKrmNmuyhpR/imB8+XRLdVsZiIuxmkQ
PdNmrDg30eZPgRHemAez9Yeh6ez6Kc+hFptR2fKoW4ZwdFuNZgVv6QrzyIUqZPJk5b16WLsaaXYf
lyIFH3mSjWmBT0oxXALgDAAmsZuDM5OYsC3cmlwfZDYv6EtuRXVIWUtD4yFIjmXHzvgLIbLuA1V7
OlC61QvCGNUCvKbHPMF0YFhvDtWSRftrxWrq+qmNS88Bt9LOL2NsqgBgJLcjld6iScWdL94cTSTX
YsWA39+kzBD2sA9Gnv4vmDUFBK9p9WgcMA/+bFTT/OzcbZwzn3FovD0RwRqKEQHY7bb4JkxYpJgB
SNN8ohr1Z2Eq2ByL1r/PM0u1HykMzuDfi72WUVzuR6s6NioGN1T5rFtekSPe7CqASZcnOlbpbiux
G6MWajynA/VX24F851mCC5k+4JmS8pwhc12TEH7B0rFmFEH5DCqUrTXw9Z+ajUr+wdp8GXy600UX
+3eL5ZYzPO9ent8agMUkxggwAS/M4rgk0mrU71M/9080nx65NMw8Dkdb9l2pb/zQLgeMDq3qB2K/
BMKYn370sbW0kwAdaMDhiAxDlgnmsmMMgn3DEC1C39l4YSbDt9Mj/1qFFdbFg2EdYtRwchKlHlWk
ug4B7HecSvtnXR3786+t2pVUJ6DnBx6dmUJe7Fe6BBq9JmFU+NkGZFkppe621FTdcu3/As0Kqbpw
wlAYt3F16hbA/Ku8DI9nFDqxd5eQVfZdZo1CEmgEWab/660ueiewRzToAxpoPsH/jvi93L5vtXxI
AnzzH4OHaInFLQkHheHmyTAPcMieif06oQCEspVhS4GvXnpBvdAuweUaV6kJDR5rAB+CbZ4p75J1
DjysdqxVxUEyWj8Bufuc9oVSHjW1z0PRiVlIFBrIrOv3EgMEnBrjITfE31YcT6wa3qxTxTuZZ0m2
fPC271U2uYjrzo51g1XMyUqIIAC/Z69ULbaxvpFgMZ1UMbUmvw53Q2mhv9kVtmveKSMUWsBi7p90
GKNLLDhs933RiTPbaMi+WRIScKkbZs6GncG1NNaK4RoB6F6tPbXn36sJtaPeJq7bqWa9+6rY7L7L
6Ni+y4cyicp59+d+aLLtHOo8pZ30JLQWGyvliZUr1H6CxaqwYR0pw+/aW3ExsitQfxukmbC5CGu3
hz+D3z5yllKB3n+1AE5JuVRxFtdVKJr7O1Za5StE3C1cm0sfLlmUaEJImKwdZ9XVdwlVjdTGadbP
wrat/o4vClUoMewX3L/oCEjLnSt+aqsDviL8Lkr9KH9axw/MJvPiGZVRCfz1ppZ7ebywIulP4lxE
lN5r2a1KczYHcxDts67ZXO2k4cdcUwD30h46yIxoCNLzy6qS2/U6k4tXN5KgAnD7/E6mrdrIlSof
bklgsIfjo8XSkCT43hR00ipuo9aHE6MuV8o6L2TR9uH1X08xkpYziUxCRDdtGSxPuinOS0Owzn5m
K5RK7NPhKKfpxSYG9pHjTcUZv+LNa+/0e4tQd7kbvxqTLSG5PTBHeWQxJjPgQwcOwpKzOPeDOmB/
TZu9GdrGA8bBtCJxDpOL5bGzOIKNmn1S95roKiMaSfoEZt8CRkJsJPAz1zw3GmwjDtTuzno2zzl6
KKIkMJT6d6Xmay9moaLNkwRixrtctjyGmnX4V4PVj8/BYDSBlRBywYTta1lj1aF+YAeVGjOvT02V
sDODMbqijDor2Im2ZJSpKnfyvPRG0SjOFwAHkuRfL6Dwc/oZAMhSJ1zENKRTDhK/ze78GtivP2H5
Y8DdC+1o4Q7Xd9kvRJAmOr/PSLg4X0GQhutYRLSSLaaqvoidxE86jP9DrCFHUhJet6Yi3UdqwL25
8teHQrGNGqkZGXpBn5T5OZXy3Izknoaa1+CLvzb/AvwnmlE5KjUocR3mumHMBOw3dNOO401sAMqW
efr79hE+zFwamluEsY0nQnOLLPCT2rT1h2mdackihiSoEAQzd9a0iGlZocB+kHB6dfWMvkoJGfY/
RzMIwQPcZOP8Z9yvXJYsIgyLo8FfJTgQYI2w/kseUXOlcn6yCYl2fcKvlgXD9O/H6YQzOdkgD3EW
2E2lS7bt7m9e7Aszw81v495+Yh1s63k/PC+2PhDD1P8wm58e84xrqa3jDiorQBun32oWDHF20V25
eTUWipWx03W1Ir42uwG1ZhOz7V6IouWeUzRRf1oVXe6JBVpt+X1duMF245WsVY2JyhiI/4CdkiKM
Nbz7QWYOdhxgQeKUVu+qtWyNXEr+mj91Fu1vNTQZIY0FQnK4bdyO+PTTdfG79624Nyi3d6rOGdD0
YoN4h3Mk1AyrhVUl8tdfidcEpbMHO3J5b3QIozzxvIMxTvk2aC/P2WTDAxV/Y4scOQ+HgnHz39Tr
0i9h1bo6IsIgzsDNGDeC/Y4/WgcC25Gq6a/LmkSgHOnmfYY5C2NCy9pTWYto6B6AU4WrlW06AsWh
8P9mGkw99DFUkbO0G1efKyhTnrpvShfzYVqlqwFfDFtFhOgWbbNOn8v6Qc2QZKqst0tlh9hfpLqQ
PvNlUHYrfW5ikGybmYZl+k4Ppi+rCVB13ci59abYmCn776Cupi950pOdP2qpTpSILsK6vNaSSoha
BoOuwwS03XOvyfGpViR50q9olmPGOOQxoNU23kmbc0Vi1nBUFvnR86LISf+lfNrdTk/7JHDXyZ/5
EOafKozfgVL/1IMtDjXYZeYGVUXlilK1d/5zTCFSva/vAxImIeTm/qdRyQ15MgNaHD6jluq9ou2B
yWMArNMaCcJvxChmlwl8kJSzExt1Zsq1wF+o8R7KpKtcPY2YCr7C9Pm46c/VtjJ6F5RcVrsXDxyu
1NpiLPVNHxAH8Kc5K9NB61bJUIoEZbih/F5aSF2Lwo4uubtnBCK8XZ5RY2Yi+B+RfHZKzdFuHalW
eW3lT7R0UeUMsv00mBZ/MTa7UPMEiZjJHwQGY1qGkVOSt5ZrGpTsvZPlbFUsA92SatGUfGlGzJ0c
qvbfGuvqG+fijYN9VfrnxsVDNiejqd/N32JMeqqZUIDXbzAkcAu591LAB3kObKkNejgfsYFD2Qf4
DaP8k9dq2A9imPKaFsLOvY5EHLL1jCUX9VS/Ia8l5XoudeL1Li00nmKVWIb+ChTPKDVjkKpwpJKw
UOlTl1nxfU/XGaym45IFqEoHw5ZDzx2Xki2hfyzHVpQvskW4slV5YMVWKa07u0RV+smOgfUlRARD
EjcON4btzlGU3S0oJBdaBtaVbvOcbPNkMWQdHmW3O93KbEqlZPCqyp81PRprz9T4AwFjPnyBz1mR
8v7tunVJJqwY3Nl1S6g/g4JjrZCP1TyKQM1w1My6W7Hyx2Ac1+qbsTNVkWb8nJMu6NSblplp66cc
nYlTTKNWtk5yAko6HDwV5KsymD4Sx0mHIxU74iyQ08owEo6qI+0SVeO2KqIC4auiWLMiOSWfXRz7
mvoyZkWiaBAICRh4ZotNLiU09djp48lioPY2+glYAw2x6WoEDDh19YgaLe0DAmcfBz2QwVYqd98c
2kBOSomilwb/3I0UyNWjsxNPTqA9pNMYwRo4HRVUAz8ONeo5O8UyYPwHnvQHpV63RvX01dTNiv+J
kno8K+Xt7gJ5sqc3+d16sE5fzbSotim2wZv85SEPoEE0zJAmRQB/6OHJskRO25uBcVOH1NsSIlNa
M5yM/+RNIO0DUVqb1QSYRICph3j8R45w6mPPxTEFkPbCagjcaUoPka0VbqOMTn8gdVPhpjU4yJZd
oFZUeWCu4+1H7LBYsbJPcL2IPDQ6vaPrHFWpsd/vb0DgjV/IdCWgSuauMchGC3fh4Q6cITAWbxsW
FGHaE6iD4yRs2QOF7CbXlUgVvxaZyDQPN2oX8b6qTws8Pzvi3/wzXfpnX0JPEa1+fY6LCbFnzKxT
XLziJQaiKTjaBxfdmPUDFLKtAH4KzhGXjFjjMjvQUpGUX/pOd0xjgnP65J9UeT6GoK4kUBVASBHa
8WeWnfRYy79pymwB2luG7wtOzf3RIXQ+/x55yDtgmfFFN2QTMCLc9/lRolCtP+rpyLPIFBWYTfs0
32i69k6/oK9r8sgCdbi/uCWa07kiTBm+xdtcLSAf1QBzJDDprRK4DkaII/zpgAA+EoY/zVemKb0k
qzOUo3rxfHvSJSYuqnvGfg0PYWIoF5DiA/HloXviX8NUoBCteYrQleGxN1C4izXK7BBob4aYYSed
HA3l82XEJHCPzMeWrMjCvdLVDUPPuU50OKzBOGXILM6WIJGuQdA0e8iwyq5gZ3c9vjDMVjTr73lq
RPUYjGo+i6azUjzZmF5pzTIDpoeDt7Z7h21fvMxNMrIVymkB2uYKz0JWRU67GZ0d3XpNahOYEaLp
07Mkwq5HCC9KptyK4HHVQ71zz5E8hLHw7ezwVwMWI1G/XnqY85w6vG4lSm+Z+P2tctzS9HCJVklS
+Spq2IJRchCUxHNyJ5Z4rkBrgG2L9PVXBDkFhLOg3Q7E1qfG9JV5GiuMidZ6KBdE5iBs3UKU/G6W
gk6udHSOmsa0hGRfvXiKcEhMVb7xssZcZEW1mgnhQSWAb9vhN9bF8l3UQrnRw2hubQ+jYLu0Dnp/
hnypUO3wRiZiZbtXmekljSrigTGLG9bWHBsef2HHadFPizDTInAZC/LzD7ntjZG1oZbcqR1zndAv
0hIlpKi0QlZZLY8ZgoaGTWlujyZ35eZdcHFh74uGuxq1wxA6gbPdaKSshuDs0w5Mc7Oad/Ni1/YR
d5cD9QLLRho01vAn/j8QxHoxsAm3njehMdKSOXgY2ZigzZmd/DI/iwDP+f5iRliDCrCkdeAMSmGe
3k09Orh5LlbAf8MSkeO6ro5xHqmScPVlrEg+/cmEZlYTKySsgcw17/FhHyGh5VeRAF+qHfSEhRct
MvjirzB7sRCUGU6zpzrMOhA9wlUravVypSFokeccue91/RUwiTiCMyS0zpbqzJmIjlUcDThVdaqT
xBtdrMT4EjaBpM7m6PLej3kDkArrqyk4mtirS7IH9PCMWQrWX/rfbsNqgRuFz0M34V8mZhvd7g1B
BbYNrHz/rp2G69hV2zDh0iOnYhsq99muYZa4h7yfKUV+SGSHxbj532AKMDfq/tYKxrlk8DUyrJ4M
CdlnvryRTqzViNPLsr8QZCoezt3txa7MTN1JYdhymNk5uEEzvUyZ2ghCQUoL6Ly3TQucqE47p9Pu
WNhwQcxZB6KaUWA9TgZO4WEXm8QtVNIYlAi49DxdDrYZ1MnjXngdkY4Ms7NesYorPW/J82FBg6ga
Z49v6bzf+BwAI94vIby4vOTS5pNpe6AVJ8EDpTiBQ9wccGO3/8FvLx0b6aWQQZWqyf7x5Bgy0JcZ
IxgrE6J5Qrq5caSytvNaoSVIwnWp7qNJQPHxDjsbce+ZwnP5bSrdML1EhhgmM8/iWsF4sxHFMcrY
OibtRAV4N7NLi6x9QU+Rbp485DJ/KTK9pWONUCAUP/fpy4RkdRg/hb9M1Cs6mvMJdkl3pxLMFZ3s
v+uXoPRAshu/gxmq6dBxco3/EB6dF7IPOfPmMmYSeNPqYYbPpoomQUxUzi1H8orJd0ZQRslfqtus
dMOAcRsSYranbuKSL6G6oTfeDkgUz16y0en9HqU/A0UzEOPmcBKNv76SCox3hzb72hlZkxNT3NMk
oaRr0de2Xg321oyUpl6T74oJWigC2QuK8/0vm+e9H+9QPXf2Mo32zV1icTG4w0BL/NkCpJD4bZjD
9E0HWg1yaYHVAFxkNtsQRUch6KTJTzwNFfFN1F6rYw7Wzj308+hsFLQOOM9S/I38kXGiCJ6zeZOn
KJ+Yy/wErACoOGNwxRRSTHyC+kRvfMLbcEEMk9fy3uHRFgD5BD4ioKrGKFXl2mCjFkdV4crB5W8+
Y3Fnj2CV2bz1CMTSeas8NPwccqLEqqLCcOvsY/ZX+YOl9TPTvt1yDOAHnmk2iIvDs+oFt2bvz6x0
2nRyHy75xmMn+ODfLVqslSmx8vlYEYDZrDUlLSSnwMF+d9/zm668muovQ0sCXh4Gh2nJuRbH096M
K4UyyNGfnkOCtc6S81QZCJ4jlNzaye9MRwkIPcjAEuK5vno0ov+6iwUDg57qfc2OoOO04bZDqiqx
QGHyYnwM8h6nDG6D9VYOqKTPBmRnriR5wQrtmgxyADNMvem2VODKxJoypbGyRmMKwy/xQnX5RmQa
Cr8ayN1vUYrNK6jCRWlEjOXUsHM936iwk2aMvGT2bkzoFNIYT6HPgnpc9UjABx2zby3D0iFvtu9t
7SK/MCuveDM1gkGTPoucK9+JmUqk6hHCcrukZsKs34Jeb3nfj6JycKfDDKr4RzIK9r92Xh5bBgFP
ibF/BgCniTGMnSCuoVPLDmYPvuBOEWM2zXaaWPtSgU1odu1AyDwSiPZFw5abJ29e5Wigs2P58AhC
ypOvGofXfssdKbpRCuLQieiXb4hbHGw4+6Y9MlVN3bQBcpiEUUgZbHVDFdmLPOqosNi6UDbiB8/f
F+q5nM81rcxZB4bdCrpoczZT2uYol9uZ+DaBTW7cVdYRP6b0/IiiAUD26ifQtR/LUPi5o7eD2G+J
sjJ5/JqFCYfHSJIelVLRb2LpByg0zFZxihMJ9UoHCMaTMjSj2smLm6U7Wqk+S5sJr6EuHf5TlTDB
XO9cwim8r2BGQdR87kP1jk7zUmzhhtxU6GYb/6Y02A1htp8t4j3IG/6HxK3jUIlxP8xZ38GuP/6f
Qn+rgLERfIHRwPNA3kW4V+XdaJuOXnuflQxkuqClGZKjs7vrAEouH0NFClpbBah62JwRIO9mudGd
Ir0xq7ZMgEfSH/XJbiqMHAsatr18Nv+n/sRa45xOJv7gvf0dGT+vyjxtBbO/CHmxoG7qTWKVBAXn
6s2IStKlEI7RjYSob9Ly2DmeM055qBqhiUCpHjxfKo1fss2m3HN6w7qcj6Vg7htPibXGi9vFUC7R
uwA8sV9QAn5J2QjM9RxLnKvFDSqniWzKwTjP3lMT4D6tyABLmX4DOckNeqbqb18eeWMytJo1vgTI
IqF4HxPPE4PJbCT3Ok7yho181n2sl3h/PtILziUmMF/01yX9sQnoSOGYQswGCt+Q3ePhRjmlr+e6
4np0mrKNTmups3Tzw+vI0OsZikfrEV1KqBCM6f55Lo/jnFk1IclTbdjpAoiMPdKfUXLgeHE5dTLT
Ra1SUu/421YqDTDtsJtbZUJqLnpVwnKvfk6lsqvlg9Tt3rNEjrGGtev3gy+1l1SdRPKiDYT4BWaa
z31jCSKVzzGp1XI+zObe2iGwWC9KynnOGLu0lSDdZ2wyd3E8aSiIwwgKl/RHGIlw2Lr43jXG2pDA
J4vtUTmfrZ/klD4K1X1usGG/nqydi6MfUVPObXUSkiugF6LDlKCuh7s7gw4VJvuLbvb/l6jBAKEu
b5EF61KLf68X/xUPuhghispZIRtrYoZYJOwPSq7ovg84zmxX+iqyynUpQncCpr9VArLhlnRWREdE
pVkuEvI1oZbsIR1pWdO3J6qSGixJnYePD+1MYPbgbv6HmKlRACahuul3d0UudL+m26UXmwYxEyP8
wm7z/eLtrQIAntTkeGZVg0yPhIeJ46hhCA7XR/9WrYo7SyqBtGuV8RTOYG+YrkXeWupMfA/l75sN
8cicrXm8AXExpfM1oQElTwxxX1V68h2m0rtBiFskNeaghSetqSOk/MSPBS0zLAyt7OGJjau+Qrlk
lHv/+9pqM1pLj6wJDI3YlaIqgpOO6VlCgWXkd5lCX/D+qJtAHTg6WOk22yF7RA8A3rNGp859KAPq
p83Pp18yzi3LRU0zEXnyEq9vKJYB8xdtNszl0EPoFpNyDqTmwt/Ylb9zG8oVy4TWCfvbY2r06UQJ
FPV8ID18iaJcc8VCRPhQ/yGmG3KUopFEU73gd0piFCOpGsC+8UDaj37vfBLVJG+iEnsVi3yx9L/2
ZuZ3m4GZ5cV/+TSPVR7DkLsqXWmWNLC6EFcwlHK2+JsEcBVKY+TwIDwk/SzvbFKfObsFV02TfyRy
kgrdLJ6+WPP+tmEXum/B8zuwuUKvrESASTSWGEwz72ZP2HtTz+IVM9qLVONY1s2UImVihW8bU1Yr
ttyoiAUAbJqbVxZ03jCO5EWt+H6SdZnh7ZfXalNjRqFtBTzzomgd/XvM7eTo9hVqU64pKQocnNSY
OFXVGl9pRIU+6uaAyCEs7hIYuU3zRHcDFGPm0RA/O7yeakUYVnRrShtWdIEyICQJqJD+b36JVVrz
gNx36Lh/lBSPCZ9TXcWJvbHPIaQ72F32eiB57Yhz3itQ1yZ8zR9n7NUZr3GgSecO64Re4qmN2C5H
WMXf4jOEHUha+Aq9j4m/Ln8/gfuZ+zaz8N4OhX+UuOk57xIJrfnwcW3cJXihHfhIXIpyq5+45LZt
+P3wZhQ9DFAAKpRlUO/lArdGI3wU9PViYamYMOWTk30nqfocAdW7+8i+dDKyqjDV+qsoGKu2zDli
y0Gjzl+LsQynYpgF7b1GBqi503GTrfAxJvSdxmzIiTJ8+PWTg1JYgEK4h4dm4E3AHxWzBmT41TRC
JjRNMCs7L/RQYUkXKClsruJylHkhGE0OubUqFcnS4hb5oF83jIbfufp75XzQTn02EWdMf4gcEf74
xpmcY74a9O1A8e6sMMh1+XT668fkclJ45KiEDjiR8fxeHYofnA6AlAkmtknQAwgWmG0Hzr9Q1kvI
SoXLpkMeoEm5cYRvGtiwD8gufW0Hi/8zams2OAEhhD6LslnjvKnPEf2E/TOJcm9o5VLCsB3KmrVP
2md6WdxWdPuxwBenWcQ9SSsxgrODCT/VNp+C0BkFjfPsTlAOfImjXD9Bl4NFmNBSht080qWd4lGG
GtzIeL4cZ7ZkrgRpCDfsyzF5uJfxvybqP6O9ggFEbhckgbgXD4642WmRCxpThVO7PK+GAKf6Ub/X
x6bedsRQN4m9e5XmpqFd4jPiYypIhJrNHSnqXhlp8DwYIItn1atFUroODVquQDGy53mI6mfowyoe
k9z2Q33GZOJJ+a97Et0iZNM7ANacFSkiczyqBxaBpAKmwgj+Qv2yDOO43Cn/d4Vp+93AdcxLF3j3
dDBCAwIO4hsj2Akawdnsd1c6/1pYFYjjmgLxbS1l22kJFZ6xOKuPc2D0Wx6FLQehh9vra+EQwObk
ZjDRq/OCcQY8iD6hYWwVl4XC+xGRzgIkL18doXYJbbcwre9TfC6NuyZ0efZovAYvQp1cxDuzqYdy
8kjOtwwN3M84t3xSIW2VUW2JmkOn4I4nZDEUR6LEs4E6gaeqpf4HStHNjRyR4KTep+9ico6nJBa0
NdkLGn9Q6aphB/8HHft5DwZujgHsOdEG24D8juOAdTwrOTJqbjfYbMd3t4vIXYKnmp0py44W17MM
0vQH/iv1WOb6UufQNDPI5FCu5nDliRI9rX5KU9mGt4cTrLK6Ei5Z2liZPALWfCIMJS1rjw3i1C3U
jEsb7ABkbNXqFGYt/muKIUyxZGgd7gXMp6WtMhZau9Zm1t8opu8HBRNTNlr4mpWwnmSRQoMjLUp2
tAAzUzAi7RQPj8Lsx0h1xihaXFrGzuZKzPHyrNyuA+6nGpuNQPA2STQqBrnyk18TSKpDYCtGm17s
G8luqRXmVKr/AwBzw+KiBta5Sz6ELXX/4Mg12jQG/+TgerIl1rojqW+iPr0uw8tG77eVqOr1uH9x
JOIDE49UKisilzM/ZTjBgiwRHENdy8X0897DukBLUGPnVpNKvm5LlYdZzDh0sFYy4HA2dpDDRub0
EpkDAW8eIzvm7M/BqSHmsj6as0kFRqj0Y5aOivnvfX0vRZJD1MZsI3jQYXkJHRE/sHOv4UrCXyZi
EjO35RszmIJhNc02AAqlmPQ0CJg3hEwfxt5IBWEkcx+ArZwSkC5LGUpGeb9lMWZO+LzIOUDcv2yL
N36CS8w0EIDHkOhRUDyFRYKFin2QOnHXwcFPBFNV2sHOqHybL9KXGDYSOnFlKwOGf9juVliGx6OY
v/dNl4AMR3hRqxkjvHzNWZFbrymBGy395Q4opmR4eryBhj/XLHmIYMWWTl4yhHtprvJXtzFnvH0j
O6abUetx5MbD9m8HKyI3w9aqRfe1UYm3D1F5QE+hWqkMsltcb8oBlssK6TkxkOQAxeSIGUDBYlXi
LN3h51h6n0/BnBNKYtrxXl4sgDHqM8293JxtFI/7utBuS2DkI6qX/MRgR3lgyb+KXpWdwUiME3RJ
PdRqmfXZQ+TVVX7RpCuRKrfGU8rXrXC+wZAHx0faZWH3BtatWfwVRvmuuuTpEy3D5y73U3abhFKQ
QR/V9cnqT6HMbA+N3d3+MJFWcWBi8Eb0ImMV9NgkvgBOJMxEpgJwTQ+paaqKqwnHi/mLur3IWTrR
MEGqc80+o4fMt9fwSIsfYVKcIvsCJwFO8Wx1lBmMNp0vePllnotMRdFfEVdsaRfxZOMkfdL7Y/39
Fhoaf7eCkNd95Drs45WlELHH61eUmkjyCqPLJc5sJMNbAHpi+WLS+5kn7CYtHuxZwNY9mvqUYC9f
nPAkrpX9pfWXEeexle8x5+nMWU0ie6e6u+rpIAnVcwDv9ZymqvIxNewVTJpm4XSoz3w/yb2arBRN
hyuHtmRnRVSYIRy6+KOfuygiCuIkRaxcrF4zVyM2v8K9NSYDhNP22o3fYLWfenjukte5kBaueUsX
DB1kRn8UUIkV+jBNknZ5M/GbnC83Xn+JMkdeOeoEBukQaLc+1h9KEBQD0IPmAGZzqTvu8IBi03ea
bxMRtC2yarrECyzMHlPqTQAxGS5kPke1swEMe8chp9typ+r4HxgP68CBNmziTuje7DvvbLFmuvIx
D8BNSaNGS4DZ0qkpKLvArRtSjTcCI1WS77KGXL2l4XPHYwX9NG5Dlds95dRLPg1i0coh+EmhVqrx
sxYMtvbENFY0X0jHZngo2j/cRJ/Bpc8zaJnAynlRRsGCu2MysFWKLxUu/ok9q9B8q1W3Avp2CeFi
o4pRgux3NtocyUs8yAUf2vfYWrrwXua83wVQMyLcZtR4RBY161lc3kyjH+KqIDn1BT8vz2O+zLGp
X9DPNdFip9WRlanVBz4vg1lQ0LHWOIBi3meI1hVKDS497STnnFhZhinA64/DEgh8DV9WvzQQ7kmq
JArfUqhxuzVvVvTnHBRXhwVkaSh7JmNRZKqSuw8wlHOHjQl4sMWDREXiynbp9pb4LQjVdjMWgCmY
YqyBrzH4lkP3fCAL7gQ6Wep4NM1DzjiODHznw/ri686/re2Ora9ZIJYFL5fc1XLbCSRKyrssn2Cl
09lrCTrPgYdUN6ZZMbQTXI6L4NprsdmIvYOKKuapUQU4iGPtcCVwLuVu1QcODDppZoIe5MV8bycf
mKOBCNflcUXUEpZi+w6+xo8xtWLwAlp+/EW6zMhN+NI+RI3rOPoCDEt3aEZkMCoXgyN6B3sswnZP
mUWvnC00X4fwoW8enQXgRJSXjRHXEJtLRR3eGxuiFMkv0yV9sDrJDWwG2QDKYs3191bkkS/GVMDe
lzYWxXhasy4N/jjx+cTRXLigbmnRSINIC7kHkkHUdXfjYI+bTHJfNjVogrgXpZcnvUgUBNNvNlTg
T4KXDnWtYQF09SvT8lDY3kgHBGi7mLVjk+U97oV+dX6G+hsWu/8nkwwG49xRHZZ/3gbOCzp24GBI
ryxtU1bzi7kx4gomB/p6GFAg2uxSc0edOoO0rAQ0dOTIkRC/aPPlsT+qmGRo+oP/JfsIoxJMNeMb
dC9OWOM0isauE3+1eQhYEBB3G2b8sCtjoGRQmo6ANkndMSUa1oyjugbEvn7rf8N8qqV3zBYBoglc
1xuLv2B/OvdUONIA90e/zKk/uOmSz4JNm2OgpGmICntTwkRyqPjdgz+IbqmLYyybBQfYAO8NTzYC
2lnj1ky+CCaGABdZ4G+zibDWjzVVT+BUpKZcu9esg9cjfZWeb+ble4Qr2bh2KkBQMqbdChB5qdZb
/pAYgCTG0YBtOD6TGY2pxLYjtJMI9arVbrxXroMyzchGGzQJgvn519YQNZRsv9Q3/F3U6LAV+EkC
veF0kQsvjNYv+qajuWCLmuwNOVlfcFXcuh/LIcWMkOrjEzKVgVHeBDxNKMn+kC+yUvR0wg2Ol2f9
HqeJILDRJv+1XK8rrrCjDYg/+HBV/9Ht165EpQwqvGE0A/8AVvfP1Vo7VYAHu6RaE6nutDDEaPty
xebifyDxg3uGt3aB3QKTYgpVaBaC6EvO/jN8FXKYiEn1K/j1qkuAOJQn2EiOUfPEsVhYHgEjONNP
SDuRPXj+2uVF8OpjPaMA271kZGTEaF7S2TBo1UQN4rpNLFyJEVvqdEqf29E5mNWea53i/Co4c3mA
DUJqpFGg6pnpXPNOx73XrNxhfMAvWJNwDcZuKR+bOGmf/402SxQZ/+lJzRRlUVvrrht9TqDlt6EL
Ky+XWWTtdbKDp7csHkBEC931V/5TA9sonK9/i1HnFr8THfHuZHbZyEviOfVn/mVakMd8nID6JO2r
aFrQnITkE6vNfcVkAeszul+b3yEuxM+W2Jjw67UnqPYDs7ql3SUr0xnHegKA9GCDKAZ1AaMtKlOD
TiSAHdfL7MKMASgOgG1BDkl87W3h4BeR3fM3TwDheF8CfHpj4rkpy4mI9ri8jfuXfxXq5GjkS8E0
A8ZCLgloI3Ruw0L2dQr2FHCMN1O6BWLfL19GCXT/j+BNrt/fFKAdLi622X1QBAcCYbwAmzixjk1W
fNmogdMpHCT6R/b0hbEAvQuq/DPEi5v9YuDDThT0tv/D07fa299kqOPn6VAn9FXL1R7WjHepmpP3
JxQwxSNdUy6hev9edQdkdaWaADj44pnHBKngXJN4k8vpcIfUHlBr4B7CG7snvnQvpknZ4+ZcHhMo
DLCR+4Git6GknwDKgP3TjmWcIK4/aGhwjESI4dbRkp4ampjdSlZ0c7lgy7ABPC6v/VZoU5rKPLrd
4yHsezz3L0LyBsYjYOa1c1hhtDtg8rF038OtXojj8P1yt3bzLBMjKxFGwUK33c4lyRopvF3Qo7E+
V5Tte1qofOTFaVgONrBfm8nnmbl6BVNKZLgNnDbRro6/sJWLF9jfO7PF40Car8D4mwqnK5moksNF
6WhrHntZ8yyT+b/2FyyBTTCHbeuFqgSjFL09V1aOF2fWXzaElURsPWCGP14+ww6fyzAYS/1cThwr
vFIuUhhcenqf9FllUGA/p9Yv3dNl0ZQ9G6WRC3JHRJ6Os0aIKH/cV8jGEeSroJqMZhq3N/j7EQ6q
qB6fLYagwXy6sP8cDkmKmIqOVH2/d7eJ9IwV2uFYWTKSJ0IXjEn/XgkwbYnlraYFKQR/WjroPPl/
h0oSpIJEDY0LPXy4HHCjxNmfJS4r8Pb3HmgAfGUSYRyzgdN/lZPwZ+Bv50QjY807p6fz4liZLYqg
fco62Y8hXLlaaCge5RdDzqMQ7fFkNyur1LRj8PMpLfPoz8UvspnmjfpAxRG7rwR/sC6//zW14+vK
q2U16OJPV+trvhCHEJMFJtvVr57J4q5AMZt9EpvrtkZg7OhfQ6lAd/uW7NHrdjhslOXfGZ0cgztL
eUy1aSGiKBKB2B6N1bXVLLdHPQEhJHVyAEBy6M5quPsgKRbv4vtVjQfNVgMgwx5ZvhKOZOzVG89T
s4yzFlS7EbKk+WQD8o5fsqdx14IMLv9VjOh2SA5Z0LXzeyE59UyGwfD1A9KrQ1oWQakcT7PXTbuT
rJz0Dr3dDY4Pod3Tcjv9QPGmivQw8KlTPEuz8/z24YMgDB/kZ2P8pBtrF2esSPkQFufot8JPI2VG
3EvSgbxIDyGhs1xDkP5VmuVy1Y5xa4l1npo8uHEtkEMRTe72oHkPLtxoqoWvvuc15tIS/sngVO0K
Xk2KoilwUOPT2BdlhGFzQRUfmJD7yapU6qUqqP2C+m1vm+wtpeQJApk/N/EADpSwwPrImiklO9Df
qTMkTdKPKCQkR18YVZCN/AU6WArBGxh0aTXasFeWxTlLHVSIMMDSx4MifCo5+GMjoaMkrw173po4
209tWImx8dMcytSdVKsGBVAdGofH2NVw2EiD2q0NrgjEPEY1hg5ncgRsjYEuphj2iws3P2XetIw/
APtMWf7PDxKtic/bXig7MpJCqsVt041Nm6FLJFbZCrzojxtSuNdiHYCHMMZ8j2wPMpg4aGyDKQWf
cf9yOI3hgLNCbqI9dQaZi8EKxFcOK3K5fmEEWrET0D/ENY/mwKvw4aFP8llr/7WYuzlHKGApQT9P
61GbGAebb8hE1deqPh20jZgtxiOuaJBFKB2xNMnnDgSnyJic7NgwAK47GjVfVMT6JEXe6MUMgO3h
u37cvTEjipP30SIDCLIv51dnBeIWFBdFtvo9B69g8ZSGfP9AXlg7vNOlAELqvQ+ceBalknKWek4U
5yOSwpqupYIkfX+C9EpLbYbOku7QrIf1scV0DNAoB8MiqrEW+DT7OG7wnDkLZ8vHkQ2kpvU+BQEe
4SdzX3Z5UkwF6U9FsH6XPpl/PBPXwwGSXvzm86iSHTCsisYC3Jxcu3s/O3y8OXImC4EjzzzD1VaU
iY194hLmp/p2vqhYhXnp2/Rz+LDvhcUMdtd6lvgJ7FbZz409cHouAVYhkLkHr4AnHK9m+w2atTG6
DT1fQwKlrMzDl0JE2TTMS4oiFkhFHPqB8hHie/gZ85Pe3LH1whCYPjzvG258RtJC49NfJudm5zwi
LkcoVxKPqkfLz5In8lIvxZZ9jTjEx27o6TlnPHK3BfJY2VwnxfOlLHuBF6IPlU7fBr4BZbxw4SoQ
Fl4tG4OJ86hPOISGHnQ64Z/X3VoXTn5yheVdnUDRw0IE/Cn+KUrH7vDVk3i945WQmxwS3VCezPvi
eKCmRgrXdqT82sOdHznuDCllBkPFvHg1NQiItVDRm9p6VyYKdLmIbFE56aR49kXucvokb4DGe7MS
HvddsI2deeAQEOu0+bi6Krg9F5HLnsSdWWF5HB/ZguKlYVWvc/qNaYm0LwBRTLUUdfmZUhCpGVMe
P60Z/H5RnP8iBPky+CxrkjRzLLhWd1KbKVim+BzqvjDPDaotfMl3NrMxSy1/6K17jZvxZhAGfiYH
t/mpTudTrh/sxbwd0rkTT29E2ZVRk4UAWnKMR0UXCsdgCVtuvKnUJys7vST8yrzfYSyT75nbFpBh
NXq9NA7lUIxNNtQjG7J9QFHqhjV0NSsE29tsn87/BQDEQNCSVeDNmzR5eG4/xZsdJrYPcyVaZMNK
7Ib2a06I35GEl7K+DkANKjss21e4+5uOIx8u07l6sVbP9lcH8varnvSbk7hOCu/Faq9tDJehj21p
M0w0jMn8qZw7Nnq0CRgu9MpC3SckqhN99C/iP8Gfq9OHM0Nvs0FmNpmSU3ByvKWL4Ak8NqWo27WR
3cDduvdkeMVsyzC8xz/xY6VfmpAnZpJNNadM0uQM8LdTQmAhgg0SKzOfXoiZiGVA/+raqxPZvT+m
1+BsRJfAOVcIMwQ8m8ud0/oboKbpmytKD9xzaatH1Idu1bGBW46jhqZUt3lPXnlwBuoo6hO2KFpx
7vtaWhuyXEwRH6yG04L/PjCQ5wU+y2AAmnVFvmgjvNJXKWPFa5FH4IF2cjhEyUHCZRB1UJ91HscW
VtshCrbximd7gC4e4j1bdqzDx/YXKPyNlCtrelc9n65M+QVvizIfFtwFzMAKxfVygOhuktdbxL92
uD4fYF2xKj0FAieh98SnbnKUHsr+6Vdib0A2sK0Evn2cfDN6h9E3BlrTLDwfsBBDjf29kuMyd4EO
gmOAzUY3Va+3mPn3h/5l2wp8riT28i807I9NzorSmzGzn0WjTid9GTdHvWBv/p8S7ci82y1F70Xg
jHArLQZ4zx3dcYQTG8tRmwxjJ+N+ENgk5xe8XhwSBo41DGn6ofUTJ/BxxPnO/ROpKevX9LVNdSBb
2zeQtkRnR24wk1Xt7X4ZdqQRazjkN4XcafpI2whc7BZ4sKdx7fKWmVZZKvutuROPCu7w2fjApx+d
bFgXcekW9pyzByzgPtck0ESdL2LZnV6/vpZq17Ne4uwqApLYlTFAE3EiDFXIteCgrXclH3evZADS
RcvHn1SNqt3tZAabitNIJo+lvR25UKtxSrAloj4Wv5R1xDa9bzD5vqX7oEk3JErfscmcdeeyJQWK
HH8NVrYRUzkeSU6R1toN/eWJZXeM+IOgFCemqeIfLSC+2TO+Oa6tK+2I4q+O6UyLikjqd7/tTp68
cAu1HGPTh4MikH8CSzT+gbz1+76iWii2NCCZY6UqDqkQGaZEPzTXbygZTkRiYaXX2jj3MarvYmKS
JoYe3OG3WUHcw60eG52XStEyQJ42QWWZU3vOmcu9vrM9kxLifN/JkpiYFmuAw3GHw07EuDIB8nSu
IX3u+tHj19nyoqkJHE9LU7Fw9bWsrCkI624eQ5kSMKrvufTGHRC1mdmDgo5vmCsJrM2YGuNZ7ZYz
9o0qzNeJSin13AtYy0zNsr8C1uVSBQSh1azIycD19qbQISPC7EyfZin5uvtSV7rLN3kKZsk1Ypdg
/+9GmoX05YbWV+/1VPkcKjjha4Lv7q6k/rWsYr5UZOhVzxKPlQ6llpqsEKcsazshJavx4ulKm5P8
wH/PH+hd4QGK5wZVIVLlw3Yom2jgh6/c04wdUruDwOpc7zBxZR8FDb8BfHr73okXKofK91vj6J9Q
nnd8m3qQTRCHEp3Iucxd8HgIa8Hwy6A0FuD2g6bLdVo+P8lW2YCEEpHOPXGRag8OikUggzySYfAt
5id79n9kupPGu80Hx2NCEWCuhD/jlnkPZievemy9VzYdRNnkSfeYX/Bp3hq+oq09LULu0jfgSUDN
twU51JeCj7eO9cg2Y/xt3vGaXHUMhPCL4UlzEgDX9RD2OXqjJ6jDW5X+LGthFHA2AhF7UbLtwoci
X+80ZFqbT6RQFso6oqi7z2CJKGvgj5tk9yVzDngyh0kQeUWOjMI9zxhJ26T5Ay1svk+3WpYnESTn
kZ0UucDy7R900t962iVQG2gIx7Gk52YD42CIVuIRPCMktYZu6qzdnmHDXs2NW8/AihhB8qkZhOdY
D95Iv3sm1kwxOKf7FT+IzU/pQ9qfdFIx3bmjGuz+X12tk8UgffQX7wn4Btw5I9UL+FdqPBP0S8Ol
fD7dz0vgkKP5nkFXPRPfXlWJEl45xjj8RX+oT37e5S4PU/rquKO6s4LN1+STcbBaVEHXrFMpEwG1
BRtCDZ9aVCjbURyVARn4jRbAr7/qIImVoACT4CxP4c/h+lIZePSvPiOtt81Ik0nrdckay+Obe89V
xOSiViRhf5Qu0Bw13mu8CrpD9egCTtdowFnomaFUMUvzxgoAdl0zn1iHxei8aehmXFJdPU1JEfHy
4glID26azRJ9OGL8Lrw8D58kfFaTW8gFvCTaoB93q3JdKakxn8n5jbI0IXunshjOUPlOC7W+ZVmJ
o70ZJ4iC29HCkHTDw+VdScH8f0nVhwAVBcPVo8/jOWQbfE9xEm5e8wdAnnQRGH4ABDqdQl8aKtJG
JsGsASZ2hJHs9ZanmuiqvnWm1MnoupwbEVWR/ZouF3aXXB9i4+qO2F/mXfEXBM8o/ysTnfEswvwh
sYgQUUeJGgVZlnq4DXF9eeDR/jCcxTYLv+hLhjYfSzIW2mVYfKPgU2Y7J/mpU45TL8PZ30VZYey/
3aws+CHl9mt5EA8uZjLVYb73Yzn5/ZIJMJo9FN/M0Ys2zq1IxwF9bhIAVNQi5YZ0MtYRFAUzPpXL
XTWi434oZM9zXaCTC/azdZIOJ+vIbUDVT/NGOWzIg51r3bZN+kyrOEZm2pOwevfFEf1Hw2HGZnIZ
k2fkGAz9St86G6qElQ13ftOk9UVDVv81pY3/RsKMsssMos7rTIBLpYz37ZghEMFAx4hQ8HEI7BKy
UwXaKy/Yz2pCMr0WV+T1jlwl81lJPjtW5h4bJjJpX4lbT6aCZk93hAbFE4qo4c/n0rHxNLab22Zo
rIe95LDHnaTZuC2Zyw+3oHPwNbDbgNUw9cmmyI1irnndRPkFjYMmIM65OFeFKIznqYrOuWSU9kVG
1IioQF9Jkhz7897sDULCd7TL2lE/JC4uM2eqrjsROlOG/DAvJtIY93IDPPaMGmuzn4r7zecp7Ayz
tUgNZn0JLkLbOK8H714A75Bk/8TZAXfyZIxV2eiffgaM875LOBHQkjDE/wPHYTc2AtwEvIFHr/no
NX8TlYDbAd9EWTS5vth8NdWGRiAW5AI+RAyYkgbu2qeW5X0PEQTKz8W/3571I9JXasZQTT2vdsaJ
zZRBesputdRqYVhZElPsYdTQIDSvwEJh6x8zKL/YBg0SGiA3Ujg6KVAW8SeYAEAFVcmykfNEEuky
bRPmJ7YqnFeM1P9D1oump4/IPWR9jXxYOzVrPKUDlQl+w8cnWGown/e/3jpXgpNUV/7dG4SuwHnE
iF+8sLeJVoKtSBhxRsyTf4aO+4jojljpiiEpSeKER9VCpqzDqbpuwYdNiEgBIb+2G/5Zm5aGL+6q
8TnYXzesxQl7tR/KSoQpSO+fUYCn228NH0JEVeXH8u/o/jj9aiSCmHmcRlegVpcJ71yCDNC2ZnqL
1LKEGMKYrPY9wJ6WSXQXOnJfHzumcUeIps92sBSDhsLoTSC2IsLsbamEx4TeiT/ojps4UUysyk5M
NDs8xsC/Mb9fF+v9Wmo4rClIhkyh3sMzWv6uGAuUJyD3TqKJei9F3oxr1WbQ07DJgYXowcH6cYT1
FA1ydANX7XKaFVxPw7ce/6WeuKqbOzH2kHYjGMPkrH8eTvbE5AEqd2fDOuU1ZBZnSYiLuD8EpALR
1q62YWtdaLBsJbMWAAi008cWFeJXoMvm3L6FpApNEFM6sS1SBOl8xVkXygIx2TOADoiFIWWZqaqN
hzR8BgWtk0RNNxcnS0FnnenMTFdB7637HZhfuOvBKTfnh8A7EkTYE1JW2qRUmWnHez2SJap/3Llb
6zoltV0U0qk0GdxL8BuSXq0+mNtDVOXrADlQo7YdVrvPtrrWG40PCU/jydBGR/srgq53LJmUfM4F
TI1+kk7gTBDLLnecq3d+Yk3VC4ZSNwAkrwkNItxxJbdVbA0/hvydrkpnT1KtsxThvdPsFN4BiLwD
0PlmqPCdodp3uBKkYK5cgn5qIIwSNQNiI0uvubRe2u7Rp9tBOnmkD47if3H5qrFKyvVayifPogGv
wJjtJHIXtWnegaTiGJPOPc3O1LyEPNagPZrNyX6IMrqmUL6NQnWpa9rxmNDc3DfF+b4TCJGj8EVd
9Po3GOoxUoayTpF1t4oTtOFJpIZm/CcGKyU99G2fmn80xLAlHtpVPejlv2J73+ram4o0fJieqM90
yRM9X9fcQxZTPD9PSZqPOP+SqMyOpwGK0QFHnkVJsj2Yl4sBqPF1KBEt/y+2Zp4HqTmPuLQL2GxU
rMSVsXvAyub9RERPpA+tQYkeDEMRE55o7e+IAdrVvEplHX2g0e+RHie3JclfB7CZNxQl9oJs5p3w
Ln2WXZNWwelyLoae3Pt5iFxJtORXxZr2jIk4xmBRAE5s66pmzbDJ6cx7CCpTgKmT/nXsby3YC5Fs
EA4XgK7OkHpoTY8MRymZ0aYRvfKKqH7uoYIUwqcwOBkXiWWFKKx8+LpGGB1xpuTdzJirDTbUnz5H
tno13PGpyt648vl4jlU22hm5Q8IGf8m7Qn7BOqi/3xOowu/HfDcvjnhkIE4QAsy9fEJr6lIb9RdD
xh2FwnVscut7KviIRpLH/ZKgUECowxxpIsJeyFGis9aMe73pBvklCH+FrLkPJXhfH+5mGkGq9kcZ
Yk8JlPoHSKc4pF2czTGGqbAsP5mnZ0YvZslCpISj+4x+rKk8m5pQ8mDFXiz0VBQDcQZXOd1JU3hp
N5Q6O/v2TlHFnlqXf2AczKUyuazGdJEMO8ILlC7XDxp93ocphzpgGMmbTDkdvAmX+TdGfMQQSTc8
MQ9/mJfsq61EtBi3gkQ15JIoN0ZCLCE7inO83rg3qkvaYPY3e5N+IayiMCQUQo2vNJm0IZx0XDaZ
0OZZbWVM/G6om34MgASF9bCKDZpAEOB9nOE3XzgT1saX88tTuLvQNMa/BUL4GBS++pDQhklE4+cE
hfwf/OuHHluvpS50fb0uPBoi/88Wo1YtxfCfFfVnVlzjIqyr5/xqHKDWvSNU+Mu/xfHeH3pHBtTL
8DWnysikEt11s0Ga58PuVaDNuVATE9xHN43XRzZx4Es8KYDXlGjm5uC/TYC0GRHTCTxCNPpapCSO
SkeqvTV+IXlAs0whoFQRHRfRQVvgvHDqayofT6q6BxDg0vBcoS7tLue1plJvkb1WQ2ZLgTVohLQF
8zyohbc23XmoFdLLcr70y0VrFN0e64yhInU+NO1QvsOJPFWFMt/MNJHr/0M6bQ/6u7Ss01JKR/Ui
G92isNie/Rel1FsB/BRY7PFD24xKbD+gbtQhZxcIarR00hqc9senF8P5QSFCcOPphTaAXoUAqnko
3kuPcN+YFajDsQmesCUnYvhGRocWHPvfI/wFb6eQVEkXVzg9UunVE7t6bU94v35Bt41HLTPO0OyE
dC9hY88PFuxYIoFhTyzXkdYbRPKT7LuercAJQuGS/VdgEDVjrrrQd+cL/lEpBhNS+0vqdZFfqRRR
PuLs2b5017dBh13nEaDNRLaMnCWHhUy5qq/0DU5p8MEK2w8Ba/kGgdeEeD9Um1zYaTZfchC9ZOZ0
cThxhSjjLqeqlBO2tSjbkBhGE+cLBR8mcUvRfbwchgAjyaUVAbEykA5sSgOm8fyKXGovGjzG30Cw
w0m7c66N5CEjh72i7pPrjW5D6nGwjdPS3qKMro/QaFOeVQ1cOYKRrJyh9SdHPLONx3FMHOCVK6hs
CNHUE3MzWH6FCcxL2sOS/l04evSy1Q/rg+KjWFA0EGO1Q/h0a9dvSsVkK6ln1QDuVGOj2bt8fTPn
KkS+G3mpyKPveXZMMQRtSmdAyKegNPr5mhtSHGaPtpv7vzMI5iTjUTrT2cB1s2INrwGi8OoNLx1z
JrOcneeZWqtFhd2Akl4uLjOda/hW4o8MUpdEZuXOehLB2xcslfe7R1vja5IkvA+MHM+jN4u/1Fpn
SWFPNF9Lb6TBl8L2UYyO0Wzc0bn4bqesQp10DIeHWzR5faQkDwUP6yhQzAyGjlswVXOFto5c0bi9
ZhpajHCyfEQgeiD0T9aFzoVYF4BB8r429ZsOe8c1AE3p+UhG5SYVBQcuVq61quG9yZ2Mmpo1NHwH
GiMDKj0rEv4Rs7+Uzhy8c9ON5YTNKnbzUHDZosPY+GmmcZNHmpoufEbJHqHxhpFQpRI+fadvOths
8BY4zkM0lDF0RBuz0EbXz6fqi0G72P4LdMSWFriY1JGI33gYTDVacoXlMwZ85B8r3MvWCOcFxn6T
EIiZN38WhxwY+doF1iusOW5XV/8TAtt4OiP502r/V1dEJWaN9KnUQ6T0bDeR0WbaltYRSNtWd84a
Hj9tKZ3DwkuFpW04F0DkN05VHymTLbFvaSgqrmlQjnkQHeeS+tMwNNsOrGkqfJYvXlh7jA+oipVc
eKhTkjvXLwljq3rt84q6aUuy+mHByUSf1NfvFFYHw7I9k51fdee38JFw38oFp1rD9ESrYCuWd7Bk
mXzpPx9Fnv15/AmLddYxM90q+8UjJijCgDF+XZv795mnWov/ulCc5Z89g5QuulZ81VG1IRGBWZMY
PaRrMH9WQ+ktB+2WfgwtbjOvJC/l5c4he5TcTID1WdUy15ObRw263k040eYXrXkoYkuJqkoBcO8T
JPsKUMmFXNOIXueMIanDOSZ2b69Y9Y2uK8OEqk9/pF+XrdluBtPTpux1YwLw3U5xO/gOxJMseVJ0
gy0/awsyM2xUdi2slztEPgs0322fmCOUaUDYy64jxP6X1yqA6Y9cjKkirwIaYFOgTBTT+eUkPREk
gmNewx3s9LFYpKrVhG8z5b7QtoxRkX/4Z6qIcj8q4EDhuahADNRW3l5N2b8EHnZ+jPVfNzqGSOFm
d/hP9Lg1hmPV212s4mjgf8GfpTqq3sBlitoaiP4bgK6VENPXuropADtIS/qCNHl9+l87onmqaaMj
Xnvtf+ljC5H7GrntWFu86t6QUXGaYwoFNGNAMz1DNFUM86CEKMjwln9z0ms4n6NJ79pXfM2eR/Dp
88YHHlkYkvD/a4BF4W5HwuC3rGMiLrle2cTLN8p0h64qCVNCHe90WKeZ3SXmsmrxs4m+8bSGKS/R
ZmZrnpRXmfctXcJl3naKPGNqlO9HYgS+U8lhl2bm6+JiAOuS+OdS7e8SSE8sRDc5gfOx7QaiCB0A
XO6Uzd9UBiaZKOhl0bc36Lz0gVGJGzVhN7bK0D5Qpb1bzeN4inkF8hO0PzUiFddqehN+EcoZxxam
crv5+tmWd8Vzii2dMmB7/9jUwekMZ1T3cu7Jg+63eh3/hGIR3gSCruQePt59ISOXwEGegGqZcTH+
u2LRyj8AU8nLHKtr/xzbJbp0vENREiJzP0K5z4dKbA05qIP9m9yzNbBDeBZ0HmuhfWiuwHnZmexe
uErJ33YasMPDLofOBYXFfLCMAOUQGeMV1V/eZZX6YTrfoa4zjVSX81fvAJ6KfRib9gVxE6aoHq9x
KpmwFrFYmYlC2G5ECEjRJBAIjtMxd3uvHPoePTpvrCDdgZWfkBHFC65bZoqlXisy1rbhCBQIPLOf
2jQxahPpzSfJnqpHmKhaapPDwZ+7GFuTQzWEha0exnYLykq8IoZ/r7vFlQEL5BD3plTa0WITXxmu
YuuHLsLGbBQWjgCUPw3lix/iF5I0J+EjurUb2ghfL5cElZyTFvEkZkUw02uLUz1v3ls6lER+iTzo
EmLmpZq1Cc4y1J9YNg+DnVgY0LEGp8LyNtwSc7BOde0Opbnkufi6n/LxSejWKjd/aicsxd2ZtUGl
ry5+S1GkCE5xKzMEG5jDQCV/QWJp6j+4WC4IbRFYIZh4SNgusOXA+26uzwtec3fLG5pMcH5TTws3
h5jTlHdLvBDTX0d9UzT4NxcrWDgXVs0AsgbMP1VUMTZPf0xPpePE6l6VVOjJScKuCtgGznSbiayH
I2NNjk8dkQjqDnzkhjdArt1QmGWwFga4zrGM99V3v7W45astsolRTsYrAhrSMB2s2BaawwIvpNmw
Uk02YVAi6u2nlvE1LrOnWNaQ3nCI80c2E7sA84RdYgKPW8Z4W7j4pZNwt/s4Rx22Askmr9UQxgBJ
SMv+lURyMRWXwRa932vBcVMAX5I/wtdPD6t3UmqG0RVqurSFA3MdjDAx8R0y/gW+WCqGUV5rTyWR
S7EsAZUXfQhdRN2rWF49K/7uT9IY06IZff2oP0cXqOWBeqCoRnwKn/OrW6JD7RiuZnS6p87Chd3f
W2zdl0dSfiTc0X965Ke7W//sNDcn516V+pIwqW1qEfdN6XIFst5+3yhqqKkznPeWPoP+SvN9NciU
6tNxgbFjkvkkH9xXcx/1Ehbty/K8OeIQfbjuo8UQ/yuoqHTc1GiJ+mSl36/WvOJo7pEexsMKxysj
lv8qojQUbm8umEOyghMdPYcPAWV4Dh6nPdG4MhDl7TTwxCO0jiR4Nhxo6PkN8E36nzFbrupgSxZi
u2XdLMmuoiZfwvXyObMPBlSKJ4hFAvSLmS0TBURe9GyrupkWb2Cl4Y7v/zfuPm5aMvTlV8teYBL0
KksKaIDCD+HGVp5TATJIAXFwzEyDOYwBEjA5d7nhPnQ5/rjKeYkb0+i+YMZpLNu22sxzutoMKs/Y
mT/xsK7I3yZsV6UrvOR0gXjqq5XjZ6CK14vxuNRX/5+Dc9+xbfSzIhBHlR/CEDUauKzJGfz3XmsB
7BxdM+bqG+8u74/tCyepm6nYooyaRc7QOQH0LDt3VEr5aLtCBZez1KalZYG/PtvXzjKa7KMHfV53
cWFWIftxGrQwr6e9DD8TnUvO6hA42xx/KoF923OTRacRdfWYRZcQJJDli3HCuR25UqADwAYrrhan
a+5ULH8IiOABr5D3tVdGuRJoHFa2OR9ZK2bUjP6FkPtQX/YCav1xse76Iu3VPfN0cvSFpNxUjYXc
MdzQgLfpylDfuiaNQ99urw0EFc6Fnqfk79Qgyje29/Wsr5NFxj2bfRW8rzd0aygJ7Y83jveWKt/F
/aWFcsjPZxmRZamXZ/Y4RQC2iM7iAF/kS+1FbEU9nyrLkD9hL0iVAWUbRPZpsFb5MPFGRNqDcEFi
qoqw4Ud84xSvnseB1aaTq3wc4M4Zd46KWCWClSsrXpRd29q9AWl77/bOPkg+kCv81/3vlHBWiCS8
z7BHNz8d3prZviUSo8YpyukFIuL1/5QALY41Rcie10XzNVjkFj9CSw+zbMkZoC5PjzkvmfUUFCxH
wyYd/CQC7GHv9gzjs84NGQEDqet0ckybnHENJF6EY0yz6MtlUSQSo2DnJjCsBH+Fosl0V5wsF0t9
fNRlHknfO3fUmpRg7ZE8dG24k/o9tV5Qmdbay3DEYqA5dfB17U/apGCXzWTeGTyU9/nPOEZehx0X
cy3FXGL/RG0Ej5iA48myHQCnHPqeMiN7GQQHse/HJ0we+Prg8HMZS4u0B8oZuSGjufU7acweeSf6
UwtBy7dr0R4j7pRgF2o4OKQKS3ujxuXSeY5NMc2oX8W4IcQranEjrYt2lV1vsR+c4wOv2u7cI7Lq
1tk6GELtE8LXR33AWu384wCzfKsiKC4yHJoOmnod6n7q1QfOsdwnKeasSOFvR/Mi10pXhfmfrVq6
hisAaJ2X8CxLSVpwlKnklBa4WTO3TKZ8iZBTe60jEhwn5OtKz+SvsKCfMQs6+2lmrwM+WZbFPyBJ
yiBjcZ6Z5iDguxezhpG7/DVZmd7GGHgTuMI8Vb4lJ9fN06EsiFUK+AUT6XIGjdH8/ewXV1BIA/lk
1r0aRKVWEeCQGTjkj7TONyRULYipZ44wvIyphTfxa98U78/08T4AHdsTMTY4MwPgBMmUCMnFgLsm
jmRGXzS+l09T9NlWqds30zNucOYEy0OhWZNTIhfs4FBs9mYQtRDU1EKMRPcNiBq4nAmGtrklRcyN
z3MIipeEkrhoK+Z7OXdeTVAhB73/kHgQ91MDRd7rxpVy+RT5vWpoaKa+Oq2xFY7/RtVHgLezjo6w
FILhBiIVclv94oiaMokQTXqFP15G6dcr+6+C8yMZJ28x0ZpH7z1c8K6tZXdVojxVg45d2J1wAZnJ
K6o1g2LpaRKq47CxZpD3kJE2INJmBPTfrMDukwyhhYtR0/zlL9VE3PlnBuFK0NHiFENP/kQUCZ4K
YGYy2mPGuMXXrvSRbQzNTlGcIZPXe3W8HPSebritUYUTX6SNY3W4ykdIvxIGOinnNAeKl/yVShgQ
f+PcMpg/5u7/lYDWKdMjCI59gE3tOsWVsIpiUSwhrGkBCj7mU3eSgyXEQ54tRkhVYgJUGUmG/LoX
OPNRv/UHA3jqxubiExVuq8ErBxyQVunVkIe2ghh7nn/lOd4M+dUSJUlo3bSpgMuEJrCx93U5UV2I
CAdamunP98xVIn980Js0nLGvOns5u6gR5LR6Qw1F7wpQlN0k+wzOschlSM7WX5NhoGzu4PgI0dU/
WaHREn3YKGSncGB8DIPt3JFD/VNiQKkJ+WAfbL/cueyi/swxJuXi/LdBSaDxaig8if2yHmtqEl1F
pm7ey30tc9Vlg6j1RXn4lgE/FNVdK0QfJyKSJnrpt/svCAGpqaqWLrpNgp76jeaKgd+l3gFgMbll
9N5UFQFzys3QL0K/PRKBfW4/ssFA0+C3KjnlJYJRTbv8f5x0oJYyFVuKccn8YTQDT86bbM4V+jY8
awamDs5qViYp0Biul+OoWqEELDLSMoLrVwHQ+OxiDZPCwTr4FlmH2vzWwbZmTEvmvQ27qhaPyEVd
Iv2/DUrThRLbPllPlZL9x/XS7WnvpwCEldRxsZ+FlEOIa/6AMhN6cMVqVHL5BJpepqjGcJOj2YuL
GTj37gzJ2o0JPKvvVc+pePMHugBFzT/thZadC5PndaEalc8CBxBLE02DaEeLOTFue5rTmAYi3UEW
knsa3rGffAiEiksKrGM7zcBlZw/K+KblN6cS/sCDYnbePn38YViuuK6gRGLnzknWyE9ou1B0Kzpf
vBsfFg7R6L7k9ozUYCeKRGtzGgIbxv2HjzxfjbNPnY+OECk4RsxybWmFQOyv3ahOL0R6QRpFFsyy
i3Ye0XO+J/6yVQFMXdutvUfybm+8be1Aik62OA1+fuDHomJ7An+O29Kjud+w7oX0knZ6Ifcisu6a
5NRNFyl1e//OkXLJAdVYn1XYPWGcbrtklKj0h3dn16frMYzLmc2o3gaUvlz3+c2ZL8IVHldAYgz+
uxJLmSprUrUl1npF/9wbUscJIWzUjVzSsDnT8h/VSAox/u3BmwYEAw2J6YHjC8k+nUdC4KwwIudi
SIOa0Qb6FVuHPDkUV74IBKiq3V3eiS3+/+ogoDAOYBNplJhQNuo4zKmw3TZnqqQdD1b1gwM9AHYd
axvTexHSzvOgzsfDNZmCE7UvFFhYNc1gkT0p2QSR7OwQgG6DEs9BspFM110cmfbgyoIh0zF3i5Mq
TcmKRSwUJ+mdbhl3ngQc3J9mOjXxDObJ8SYD1zU5pdUwWLAq0e404z4PYf5pnTS0/6xd+lLnEuwl
ADZ1hqFzrqwHILV/sqnOzIiM32GSofXyeZAJ0xi0nEC4fF0ak1gwEvS6KEaIrf4tsLQDid+yc0nF
gnSn1NjqwWVoP79pL+/eAgpcnOnuY5+dF50C6LtkWqGdZJb7t7L3PU6tKwcCJAtpozTBht0ZGWuk
dd604aRvkKRtQtQQnEri4r074koyL4hCNqzUA2Af9ZbWDo3LzzAzser+0aLGSjaot2YmPsmfxK6K
sfGYd/4rBMW4iUyaVNnp+fq7G/VQFGTWPjM7wvtketH1TVhbqZ6GFcs7le+qAqAl6k70q+noeOte
q2sWAf91qrHMhA0HUDzfZMKtcEXoEhgvaSryQ1/ZEkgDsg8GNBa/JzzRc2fc6zRzRwlWYVkKhJs8
QdtIB5g1Ou4r4LCC53cKoJINZS444L+gXaUFkach+NojCpiRtfFvhxZjSI5YJCXMfrMnSlwzdZcw
IWRwPqmQAX0P39TVXRfcGfUMV9T7J7q7ADLOUsGSuEznVZ6413oEnz3Ni/GnZ6DzjGgxH/7pPWNU
Netofk80m0Ifv661p4/Fy+emN46jquSJwGS+k0Zps6EVpGdjPnUkOBZNiqTWXplgByqXwpbbp3WI
YbPOtz3VYUvRe67N1KgAEYwNRB2AZXV+dckiCznCAT5TNtTJRJt7L81TnS/lqpKh6/jR90eSOJsk
Onf+iQbMhe9rJyfN1FnY67t4n89JUg3+1gym6KgdhMTYYKkhK7UlOjSHr/HLT3Fjo+7GgYm8K8aU
PYdbMXwqYY5ng6dgTHhn8KoaYSblLNQKe8cmtGEovHrIUBbBQ/ekYOv3mQ4qjxvsryUKM7rGD5DW
MkVSYxJbzD9ek8ABBygiRRyzdmJLrPgTB5wx7eS1fDMbKem9xT5UKK6yChYQbTRIEYSm8REY1bdK
GTb8ax1KzhmFv2P1mwXl9reJtH8ZpdtJ6hs4yqDRdNMMk+yrmzl882MCE+OLF1Hz1HdJIF5tSWVm
kotaW9EbwfOdyQ5xfvHcIXB05sqJiYXp7uh0vQR6qMvPva9bCUM4ZfcUsEFvHnUHKWrIWYEOjDra
B0DEm8wfY7TQrlBDOZiePW/6KB/msHzvZ8t3MIHIN4lHqcXedn9tp5Pb5SKGB2TglW6Kev+Ouluh
SavT0buBt0FW0KAUJyhcXHivyWzulIrpQf2MjKD89xZbsVPfxw3Z3gLV2fBCxGtLa39/hl5+gzvx
HsqcZcdIKkjzlwd+lQq2xdHznY7X4+iTmBCsvTQgd01ttUwLHgyocw74jRZjCVNHJ7kguxhZB1CD
TzWtNkCderapEHKsIVj3lVzw77G1ww9RqfWBJrxLS9CGErItrH0tFTqjxqh+x/oj6jTWcPrsc8qH
aHvqcwv7ZG7A9wy3oBSq+v1w6blElwXO/2U+KeYB5hIFwLo1i5B/UNbrEvHc7eMFrTaOX1Y3CN3Z
2th0mBeN/VFQCWLFD0TpllZk/Gl5bB9pL91gwzvLsIu5XXiaFNjZYXErXCL1HE4gYSig56l5mK73
Y0R1uoi/s/VMDGQuxxAcugPUHY/rzlCNS35YB8t/iy6+zrnN9sV5hHk1a+QdeVJhpm26k3duFaWA
wrKzwW+4taa0D6ikowFL33cY4gIht6AEH2U8zaKZFr5vRuaNSvRfO0F4YELQfukqMYPLpmVw4yRl
wnz2EXXTYz46P0NDHptpvixAA35KIPico54ffEPekVmprhitTX5mWhwSup50D4HsnDgxhzKCM4T3
DMRQJUsXujbTUZ7oXzincyt6x2ctJZ5y7KjbkzCaR/36iqHg3ybNNEmZijpVkVeThBLcEK7mc7b9
VIUHN8xi+Q1UlK+Ek/IzdAdjvjQiwXtTTb77Wjdhc3xt2uQVh+QG78RZ+4kMGfuQLZEJAh9WItzI
8+oIBQg05I8EQoHmvXPJU8v9nEv8aZyo/bYi2ZEroAQDKVaNCep4c3odYql8iauDFByX40Xx71vZ
AzS0OxpsSZ4Q3FHsux8KZUYEiy1BWsUOoLzJuxlhfzxHx3Znjxv/1ioUu1c1NJx5QOlWM+ZU9fmd
IRcYNp6obsmtNMJfV5Jyrrxgc++zX2tGQun+GY+BjoZQmWMZ0BWh7m3xkvjBObb5pl6Fn6G2gDxM
Mn3zAABwTnqRQCdR1UPgC0qdcKKmi2J4Sj4pKdtzlJ7tVfKP5WWH1RmLVCoyH6i+XqCJCLpRIYQC
nyLcy2H6kRx5tinOCVVE/ap48gDP3UB+zFRlSgkLFcdVoF9pUpMA2C8APP+ff86F/4Y2yPhYhuTg
EKo/Tm1D5kJBVQDdQzMNHgp1voG5i0RCbj/S/Uv+OUarx1FozUkVBxroE0odpi7isKx7jUgBCVZ1
YUiGjkK+itElKWKaNuuM2BkilM7gKCav4QtMtJ2QSHU4U7cMPOkwW/bxzHv13A50G6jJ9v37IsK4
ME1XQIQO4swg16aiPXqdL20uxVNnIMsXxumV/ZQepZZK/NT6MYwRIn6QEVE7YpAMT+fciUkKgjmW
vt7NdklSvgTuYQeKMsSzXtIvvpmvYWmoWdD8hcCEncX1jx/PitPzGvRM/GTrIBwFV2Hlt/GXa9o8
7K2BrcrmLZb8CoGFSgkOC/9v/QcL7TyyqtJxI21xMcnmFi8VrwWWPhAKA2chQO414WaLXzQhQz+k
7nsylPlpJYUJ7Aio2PURrIluu/9Hyv5DzLaJZ+E8QLQomd8FvqELTa30UCg7F/aboqS7coKrC8/a
kCXyrTaJXSe99HwBUBJ0S7mbUR+cGrHAbNfFCNHbgm0WdWvELBJitGzldE+SaNsIrzfPcPpkwRFE
XG2R+CoAuaLGrucWfE5SVlrmi/ZUt6T+pYwTQAR5ifNijmHhcMdVzdqRZVHD3mz4iW/PJNc7sLBd
9xGCJR1RBo4uVy23xOXnQ1vMoLfoGiADDmuYsbTLRnVbV/FcoC9W8B7CfSWAQdxlNsnVnBJw3lgJ
dftF81vTvy/oePwUZVnAmnEqmFWqQJGlgKhOkzVkSw+SSvm/JjhwulVeFAP08C3G5x9vmqvxpvKI
SCxg7gRA7QiUQ7/VybzY7XAWIC21sXNjPUCVuYQYdlCeXU3Qwp/TbUgICCvywiZW0ncq4lC3zDdi
Zb9WrNCi5WdyxXLWbCRarLK91KN7oj9LUwnJ+HPI8XkxwyCzbLX4kR2PCsW1kiB/y5wZWif7/gkI
2bxzBuRWNmw5htT4YmeKhbICQpXKmhQDw8xBqmvckTz0++JCvA9SXekP3VkJrgfujavHnxeXCvl9
t3rIsLAiSlFjjAMLfW4SOneLS4lAZm9j5S2sf49xfwa2yFIgtulTLMhVUNf2PAawya/M1a2XlYy6
zM+DggB0GM/uHIoKUtT0SIBR45jUVNBXvwVrGxFdgm5oSRPUswbOE0FPZxXKKvv4n0enYNcRaQU8
aOjjfKCI/Y2jb/EEYQCHY6seFUXlGcyX0PY22wqz2lWqvU/uYK9cPe0qF759GgfkQlYJpvl2Gw4f
JPq+1/hkodNlzrnLVW98iPvoaGTqpyfTR9jk6pHPSB64E44sQlWrzNe0nHtnFVHtldPKh0DLuZVk
isphRV3J33aT3s33cbglODE5r2IRjd4+UXUMWwBOGk1o4PvsHherjUC7DKHDZsoojrGPDAKhnAvJ
mKK8ayfNhby9e8Jue4iyfL3GRPEEddMJgaJp+oHxok4qtyeG1O2QjsPCELzXa5evSFa3ZJLkl54t
kpcM8z2RX+z5UbMsAbA0d+QtrLzh90PCd3wjrL2v1xp5FeeCMAhdE7XLqBiKo/oCcimsHfIFRc3c
0yi2UPgayrtvOD5uS9YDNma42Ouzn+Rdb0gnsboIGCdbd6lgDNwjh78M3EBXTP4JR0X7II6/bDlU
TPEFzdPrTrMEU5vhnCibhoFFeZDGYRomjOfcZF/5cBCBcUNI6I0JQfVY6tYngdOyVBk+jhf2CdoJ
eVLuUce9YJ9XfQVmv6aFc//thbel+YFkcY0ShBO2DlN10W2Jf9YbsJKvD4oaSafFdS3DbnxoKGSc
W95z3gHx6JtzO4MghUn13DaK1xzj7e2aNRa6Y+Hlf8n08eHLZmMhs6XMo+Tm2YtSEWJPFuIOhZO7
5m0QhiV8rwCWnfcXN/domEJwvZzgbKT1pxLdpZEoNQwPO78IdxRZvJCZh5IAheqAQlMpQHI3P3qG
8tOsRPBIfAOyCXzU/7ZyVKIxIKMyvGWmsPxdG5DfAaxbro9t8Fx2HaYRqCpBXHEELhchZ2eoR7of
tZ0pqDYzaR0vwmfmxuEe1u6HNjLPGyKpjLc8482ZoFfKkrUrdt0zxV+aSooYtDPCTPs7QuoWSlUD
vV1oLbshatfMTS2b91UubMJvm1shKtcQOu06GcJUJIcaisdYKv4wuEj7KihW1CuIa1Wh72BbdXTa
fMfj4sCqa9pjCUFXVW4kwDyAKLA4CwzQCZwZitMRCMWVrLXOCsrJ6KP/64DK86cyFUK/v9k46DNV
B712MSVbg+s2VLu9DDCxUN5SMpiG3UvJiKiWQlUS+XIT8WZziTb0xVRLL79Pmjx5LtcSlcqOUViV
4g6OJ/0mDXfZqPl7fZbExTJ3FQOr/zJWZFFVJtTZNj16mi5ZHbeTad9zHai82xMVsxtzYkLsOY4P
6LdXXSv7Kj3m8JjxJmmoQNkJx72kk10qskN0FEmmPmt9UlTnoRuMFxQ5fuifz5BU8YnV6wJU6itW
jPmP/JEVzwIAhVMVgtgTSy0mJ39LaBxATwvTk2qFLXuHjEc/Eu4CRryEiLNJO8yg27Mdcsv2AWhW
5EHHDeNuJ9O4U52bjVi6Y8st5t4+UjfZcJ38cd24/qut3bgyTcM2de7fy4xdOjNvIi86pJOMyYUe
fBDylKXN0XlG9oWM/E6VEsCF8mMZwd2m2500sDT77QecFGF96J59Y9jiqOirRzICHqRdYROcvxCy
HHK1xs6U90xc7CvjsZ8XBsZllyCagJsbJ+UI8AhbMZ2FB3AK1f/23rYpkMH17ihMvKERG80sws0q
dVJUWsiPro5DIhi0+etcXhUfYH5kniN/J56lZ5/47c1IbS0FhJNTx5GiOfOUgkXiCBbdv64y1DAo
Dj4iPfS1awQRHh8XLEE5ZfSVfZXrHDVaMbtn6Ious60k6sqRpi/9iEZaHGFCbIrZC0dLSps6b2sv
sJCBUA+k+T/m3LYtruPXmyEtoQ0/kdECJoboIf2AWHwu/gpKhMVLzHXD033eAAoWM6YK8oQ0vNM+
ZVSFBHmibCAuUTvUOqZl7D+XPBJMwsUeVYakQLYXxnUQiUf955kZ6XWkOV1MSBesMW3SOF2R2tWc
aVA1WkbcciRo1HGvxCPRo/Wl37iLQSj2K1rF+NiD7O2Yanp/a/Bg/hVLLx5Y2BjVfsyEohObTh84
pIsRosxLizWarALKN0oBkRN2PzYT35s398lk6YOu03WABXHt9heFqdtdIAAT7mdhygL0Mn08xmz9
8XxolxwX6W9kv0veGlkLdPGiRjjFtR5GSJfi0uctFO7WUp46xF3HiTWEzE1/kHd4mBVSg7fgC4ZM
C4OC9HkFta7544gSRgIVQ0N2RG4jaiN/tzUoOtn4dct2skg2KDOETKCBHbiNmgoO33ttknsQLrAZ
PjTljanq+vjIiGunnjZ2YHgG9oVhdZyqiIZ/3Xer36eZYg8hMf6Ar+zDpUrZKQCiW+Yu0ry70SKR
7CrjIm9PqgwXC8S6woSfmW9qQi3cxBxdX73BrPcDNPMEodwwQU5iqrmg4Z14Fv5Tgg8gSiTHsp8P
cVOMb7EyIV6qHjxHvzFtQB1hVW929yNBryhgn9gbAjzOgEIDFN+tF1Qi0EtT4Kx72MiIxnzO9l96
cZO7Cf0teq//jlwmKiya+K7ixSmblTd0D7ktaLvG5yVQjtjvYB0fuBESKZVbwLEm72ApvJhnu+rD
8VWqR7LTDXFoWABSynpLJjm4D45HE4rRlYg3gYNDiwM6hJGSCMT61jHFRqvDIH+TB6VHqDxXlx3Y
RdBanCslCVVlcmo3bAt1bLhseudSbpSQnJuMDSo+qRTGhRhutMjuejpEDiDXqvryySPccYLPV1JL
FdY16nA3PBpZcmyQnrxK9Zef9d5JSXw7MHClOF+XbVE76Y/U1L5XSBxoTS7COrKmencIt/FeU3yC
ZVd+TWganiBlfOf+4mDtSTZ9C9hc7E5emL+PIKdiQu1kAR/NW40TdQrHNeG8Ni52WAIMEC/El2on
ELdlT1+zvVXOvtb02SFbxMsmfdY9q/r/+DYI/nZ1PcpwgHchEYT1Lz3c8Od3gjs5Ihoc/VjZlEBe
MP0wvd/Mov13fvfW0+ZJkvmx402cuRbV/OY+5Lbwmtgf1kIexQ6tqGLds4kOPw752uRl/AHJMmhH
9+6GUW/OL+CLOkPQlNWO44noXhdW5iHRUAq57bEfOeQmrSkDcYDI+qnngYwkBvxtQrS5QbL162uX
21gtT05pL7SKM2tZ1PAwcBI6fU4vHpWNSAN1zr74CU9kxIOzfiEr8f5xkwRjdl2KEiIwM6xl+HKg
AWH0s8++pqBF6RIULkAuiP0PHZJAezf1Uj+g2AI1r3qWxX0rRfJE9gNHER4lSUpudscUODLC5JQO
vpeCkQbaWArbs1JE5NnrpPkiRHARW5I6g+q2bsP2HQ+Nku2YAJkuNWu1EL8cra3LErbGw0rVHSDn
DYC40Xn4wNt2XFlaq1C0k+EodH0/ewISJ4TTlC7gYfmsMau0BHG//y5ImDU68VK8bK4NsPrtQJ7e
j7pb+jDQXohAUxLpwOIqcl8wdUODcTt/9XuvyQ4o2MEbuHkRXizgErm3gLeKuLB1E5M5eYEddmkG
HomLqbfJVfC7hqCw/Vs577ovWQ7v2xH1iexM3N6C9vwLh9/8mSbDfjPvKQ7fZPTnq5HIFQhSBuMM
vpiwGK8t5ZwlqOyrYaBkcW7asIOOqoyyRKWELY2dKDUitMPdLDE20Nf//MKfAO/85Ul2FyvtUxTL
znRpDMo7N0vvGO6ovrJpZEKPsMDu4uKRURelJWSbaMYiUx47Xx63lNYm/OuSgslG6oL+mOl43oWV
ycgxepbMuxZ6AF8EptrKKsZsgN6R9X1f30hw4YWc8wBg0VJ3iHAdZRTEYbSdbGy2nDYu1negBuZB
zr5jKlIqtWAN5LjwyIfLSNJgsutf2SblLC+bzOMxDEDJqitRjo0zr5eXRLVhwFtrIg3t2WELwukI
PC2m+fzOFdJeAgp27eTQnwQHdDys+Rqjek2BZ03LrAOqorckDAY30oqfpSUmi3fo2kN8FDxzL3ov
P3A+hxc/gYQUpHpL6oLNrQyb6Gj3BxMynE+e4mL0gb/P8+ECUCwZ4218XExu3DYzHghpTSb99YbG
C7idbxPbKxdReEMsgqkdP7cdxXEfJSIRuqsx70xVVmgXMkgahfM6Z4foXIoCOykGI4wErZE148r1
R28O/4An3f4FAdgAAtWMOCKDD3zbNsITY8/SAUFLwGitNdB1/+0wJ+rV8OayM/Xo+JnVp2j+01X5
oGI9MCYJqdi9EZn/+lFenapMUdZ/aEd+A1QW6+mlM0jGMRz3BE5NVuRBXMCii8+5wdoF2mSbnBO3
cGq9PMBD/5e8fMYZqNgC4sI/FMmHltrBhvPCkRwXXf1FvcmHnVewvfnHyPFRVurgP5D8Y/SN2soO
CxftpCcRcw534C+iL3qw9mEyQk24pV/O7soyEcWw5yoajSDc9+9EtP3EoHRluKeQGpEwPamhLUko
Z9LRipQY1VnF51awYw986D5b8SJKEdSfi5VJQvR30DmgrFbVHQU5ZhrAcQNC86QwxpcS/IAjuDIe
00NCJ+I/gjt8U/VTc0Hk2PcPkmMXlhORi+m5Jq4EZNtSGffeIoXIxg6LSOxXmadX1J3P+XpQ7XhT
50inyt6LANWvsiPU52sLfD5nHT2TAL/LWleo6rh9XGpzP3cx2P2Ltj8ylClT13oRE8tU+WsbV0GS
Di8V2Ey5imwcpxEuaXgELRP2PKFV5JZW0qPlJTILmaUtqyPlElwqETd7UEW7vBJ8oB3bXbPyYzjv
gIAcTOOR6zyHBuYTdGKWheFhq9tkk9V2ZhTmJfzGRidKYpiADTigNHz/+JdUtOM+ESEro/Rv3ZBz
GXdL936E64qC6cI4OIimt8xkkOr9Xq6duYOK0J/1N2SbbOAp4MdIF6Szv0NQZMLmlrqjMpSebtLf
U6DDgvK4AuA+z+hDC0JqMRc4FaDJE48tSZBjlManjmTBQlr7rZs069vyzy/GotXA+SzfxtTcDUTi
Ua2YaqD8yUXyounGQqez7EDPf0FaNQaRwzMc++H9vIMvlSCz6rIlLCmZko5PAtXxiBs7MXgEPzkE
sjfyYCOPDYFlU+y6LBUiss/BhGA5nwcojjB2PBj1forczii4HZlGhUyzQmWdJxX/y1a5xZhsPQs1
ihm5IKTIzOrC+Ab/oIPH/HneaRPDh84+43a1cql6qTOUKhfsyRnaKYqjQaOxFjEuWWeo07v3wagt
aUAMKor/eSTsBHOJnnPZ1wGmj7TDmgZKJ+ccvtoRtg0iDZvq0I0Tgvffjx0XkEiIdrgSJyNn+JTF
550onY7vB7Is+od64IpPlVT6Hvk7hBRlmCLdjlavSRNLQsYltKP8/cpHWIpk8GWab50cBb7nUu4G
symnpXdRd29asBjGEpSAzaqsaZZ/EYNI4/GBniv9o1NWHK87Xc+P8OINtgNHlvgGgWyRx8e7OWIz
2C62cy87nUSq0kkEQf/iffTz/1IfsHUGlB6LI1av35APTja2qWU0EJtRUzCc0K3fripYoqd9UzCJ
L/gka5NVACXyVZz93onozmWefAv7idESaeCfyhqI1Z1MZCWZTgXlGXpWKNc4GbL/6EwSpA+A9tcL
Pie2MC4z7U5G9i4zgHoLEPNLRaSKVohuGayGtsHNp/473QlDo6Eh+PxjNqNZLHSPM0KFGrfm8EUL
jzk8EXHFA6d0Q7bM+3IlGpFX2J5DbPLoQbAdF/3qJFO6FrOsOwZJQXG1wB/eKg+ald2dxJQp2PL3
s9zGlgRO7nzEgYDnC+7yNdPVS+WGE5xyN56eOxS2fZTGA4zoGYohbLlaZqwSyzph1L9xpBd3E3Db
esyTha9g8hLHO54KXOtRRmuYa2Jap3g0/rgrLo3n0LQ8TQzITGqQVcEuMjpjqKYb8/g9ZNnHmHIJ
X+6VrEPigt5elzYplT3CNd5EoytEpvza1QrhlMOo7iL/s/mFKUgXeoZXAOHpcGL8H8RCiSz3zsMY
XMm0KA0ZWHDnyztq4jLMNJqNLcTifAp3O3WX8AiwyXinqDhLrvpT84czD3xEVSyhpClMG56yHQRx
46zKwAdsXNHPz+/AmRbLcfEBglRxomgRJNyQ+v8oGKfTrxzpzHEHiiasdY0eEeo0B9t32Vor1bsS
vBvRt+AR4VBT20FWtNdDwQ9CPK35QVVmjF2nv2pDTPsku9+atRHMnh541gUuIVq77zZewpEx0KTZ
+wrq55j4D5W1X484iPtPk2X9GHMtImRI6pyV4PhQPuYuchFIHhF3hvLxgQSU5S5VCxrrn8S/fzX7
RKyb5Hu5sTJDh2aY2+GWbNOie5UNgtou/+g8KzJ7lieglZ5PI1d8sKeZa+HwrQHnO8jdE3kCGY1N
tCwDYyVhe/LbpVz/0m8/gEdJSEwMExo9OHSJEOpwyoDd5ibez1wOeVVBHrfbgc5LfZaXU24KM/Oc
FPKALAHis8aqfx69YtQ4iFWtfCWLI9eb4WxA5nK5+bx6f0ve9pQ5iQRV1QzCAlz1BHlQT28HqYJ3
rUMpWCrDKYybr9OVYbtpkExxb1kSBbWTYqR0U/uM6x/dREG6e8tD7KVRmxsKk8t5TLjloIFk/8ZD
RQeNvtdSwLPz8GHF7BSndq0hzhiCMHAi8/IZFURT+Agxd/AFSn6Lmvgk32nPwoEcwU6fiOYXkBjQ
VeUap8/q9eABo3KL9WIDPaR+KlFMbhc+OIfj6BGSxZxelxx9ft8b/NWJMU5wpKC74xJUHQ3YzYsN
Fa9F27jA+ftcnhXBgZmLinPPlUBY80L1YINxeHMoQYys2Phnx2Dym44Uqn0rN3hTxqCnVx9wuYSR
aQaXFdLnUldvWYfp0eI3qtIyxdiQZhc4k0V7Dtg49tLcXYNO6wptl7EZwTHshlmFh/ph1TNiWX4D
hSA6dMqjfx9IFe2PjHbypa2/aB/E1oWY+VdSalid3eXuU5dXFuN+8k/W4eHxHpgL6F5v7hYxI7X6
xdIBDZ21HwGSRnooFhVEsTA3cXyLDrTAooroGKAFD+ilT7YIyX9ia0SVd8VGr+3XWmC/4ENlW+7P
9RVcP2S4rWepceW+UDqD2sBmSWX1Ef19H6EimsyXb9WWNlMBzcIcIg1Cn0x60Uz/9zzd8F5wlJfS
bMh1HYV9tORw7sfX2FSmbL/HGc+zDrjPdOegTHM/YF9k7hp3tH4b+YriE6dR5sg+bbBl0uMhmbw2
5xR6MAje+cMaxxX5+bfuSTbv9zSXR3OgVxDU8aJcU9zDZH9oQAn9/0hev/hZbJTizPEgL7L0heMG
hgfv4SX5mzO9Rhn2h7/zqJRS7WXg2kjcDaXlVFMgHe2i8cp7XcVQm7XqDRM+H3zjy3PoMJyVm+HR
ky5I8f6is6PtEhADtRMqMinPK4U4dK0TxcZap1zOcCKyl0buVJsUCA3Wb5FTaUfX/89BzMq2kenj
WBDTdWWRDX3gTy5OV3fLZ0qMRgSjngkJ6FXXlSX0IgLmFyTFsQtdrTHQknNXOG1WrPPVxVOmkZsM
GIsZgeWUpH5X3BM1e5HuE8MzCzE/nOcGURru2wz/OZ9R3O/zkQxwSk99/4TvmLllcaavIGoeJz+l
DWKQ/dQH0yMrGsx4ldLAJ7cpzagACjSedxMTRwocxKClE/bKhe+zr+FJXBWeMlHKcKoT7DTLFn47
NX9bjyBVkatWub8eLvq6H95mMQMkj9mTABf+QLuwzSbHBc5nCfVWwjpibgSfs21Ve2J6mTwXb9JT
aJTA4eOtzBoqVkEdJjpCr3CAgschFYKx6GhSFXqMlWA4H/5+PU44HClYxVc3NQdUFkSqz1/lCG7A
Q8DXOauByZ/wqAXwfe6LtAIPACTvFmoqQbHFUPOwKU/qSUETgJWTlacKpPYeNs/NqE7jB53m6c4+
0THPWCys8hr7VBeaZ0aqodyfmZLyYcVkQvXfAA/w3QHMh1Gk4fQ1L97c9/vzBixfmdcaW2hsYXLK
Zm8e7jSRI16B/pRNIheaVHAUDVYzC0ZPJsRcefr5pxXnDsu/lNyoDbkTXcasYWd1yrS694AFQy33
3TjDkKuUSgHRHO0Ct+76gX3W5RiEpY9TPtedRCKYN7eBO+2pLqXGKI3SCvdpht2IZwFI7r9Fa7V9
cnXVmdjZMmaXP/yPQovvacyKsNhxhpDdXvMaYL6Lc9fUJKF6vqO6RLhUjZ54PA5xcVfgveOLo6ZY
qvd95pBh4xn9DWLKkkvJtO9a3o8ZhxIYPqLywl1tfTPZLuZyFqU5WVr6ekSgilQFtLNXz/utve4e
xnon+5pXv1+BhpvIx/xDGeSP0aY8IIV1xhN5oa2xPJ+uqLOp6nHOczx/zGbDsCv1qVCipOPfPvNx
FlEWG4sBdLxmuTXocfcAxzpoEEwR6IrTeYOR6luobzGN/jMXGbL5CBIXPONAF+bd5V5nIAMzbWcI
W+m9x3RZzl+//O9ERNDza6e9BaAmfjzEWNJERf/+yJePdNlzs6x8vcIh0Xzk5K7pY6/HUAaVZAVK
xJXqK7jFNRTdPCHTEv+uMC1aX9yppzE4UBJSlYo11UXT3eqKOpietEXIFHBt3k05t4Emib2MmSwP
07QahDpUgLs0WLHc+948WjRH73SPfpm9F110FHanbaBL+YtgdkXd9kILh3Z3NEHiuMTLwYBbv1YH
4dnSV7O7aIuVTnvVO7rbIzQfjqevjKAe9CDniwsSDeCihNdrxRYkm5BddHlU96bTrd60nkucOGSP
dK7N81paQX9LLNT7sHCwFbhsfdGWHueAT6IkrPscKglXKxaw/87Y5CXuoi/ZBCJBTzsK+bdfSmFU
AG/d4nuiU0hRH6kXnIxso+FMBFJPCw/rvY0t40FeKLo4h9uPw4sv4kHf6ifte0I2o+e4bbenhhul
3U57M5Czz+YCw3vJPry5qu4wb8BTJPWbLe4Wnuh/3YcqJoIeO41M8fkCU5MxfhGP4rrHsISWylp1
YnWQPFUbC7ujtqMNnWgli4KbLFSlGrBjLKzN4NpEcz78W9VCzcIqK1X25Pje9W/7C7DnxiPo+m8x
QJlsoTb8kFglNV9DkLf+an90Xq+wCA6XwfWtNsn874OBV7rZmBP/4DJfXYwcem99Cf7RWiAigsgJ
CMC5Qc9mgB5uuhLZEeChdXR572oHA/X0q1D0Mwr8bEyB8cArI32LoMGgAqjtAcp5CsmCvDJgyTBB
mppFFlviSzlrnkjEzAba5SMsGZYdfdaqgHejmg/LH+E6GE4JD/7hvUm4kM1QfeBw34d14qWaycdt
TM4x2HHCqWrv2SdzblSV8jjYwMf0BRhKIkh6E2jpzulOQQ2R9rXsAnmV1s5/r2ZIxzr+peDENILP
79lU+b8eyt1cmB0Lfb99LjpKqAmitHIyXNzQxBLis/2s31Sl+y57AWAqysMa/9DdhGN7DRUA4l8l
YnljrU8wJV/H7OP1XQaPHW6b8MmxZwUIHIAMTkVz14Z/vKP6EwF6r+ugBxYRKbDrI78DXzkQRJzl
Vt6o+9bZH80zYcptMbJOt/mLBt5Khc6VczpNFcp1TkJaLkbdkDtrcN6COIUGUV5mzUF9rRSWrXAp
qjKdJ1YcsCcmAEal3JUlq49iUDSJRBwt+SB5BEVLi5dDlDH3yHqzHzOORubLa6qlYourVKUqXwWM
gkzZH9lW4SP291udCDvtm0V+reGnGV7K65Di2VUIVWr/uR296zeb8ChhtBcjDZ9JgkN19PuGs8Gf
8lOzZ1tV+Lb0abc2Jh/O2xmK4mvvRpRelIGoWw0BqtRQaDmO1dOOrjnk6eY1z45yjEctRdnyvlSG
PHTOmGEJOAHJ944pS2w/6IYrPednTFY+/ujb+1eTanxqMI+jZQd1UcBNfgHQeSDdOjt6cdyRPdOa
k7mBUKuuJcFv3jLUNCy5+QU2ELlfTjPX7nr9fF625781Yk+WnXUl4vEnVD2XSsknfj41Nk2ez9rZ
gqk4A87HARypUnQ6AMM++uZCULSWJOOyBda4Ilej8R7HEtm7plJno5+XQT+R46+SWAR2UuYCPMVQ
7grJ696AV5/1cVkJuql8oMuT8fBAOWnBIBnpDMVpBntj88Yum7OCLbDTU1SCgZyvr7+WTMAKay6O
XGNKN3/hiL8+yuoZtZE5USMSLc6U0lqlh7vJP7BWHWQbnXPuIvAZ4cuC0C2SpPCsfQIDWBJZ8ctu
F1MQxVoCRDa3loN8NXrl1rbOzLNPWhSN9T+Do078RroAfk0PpPNGlx62HDpBOHyOO1hqs7WDDz0h
5XZlCFuE3NvJ5GEjOInB25UlHe2nAGzwpVS3waWpomsskyZmLnPonygnoSv4Aw4Z32d370UhH4a9
9TpcqEqldok5RVV4B6PjSxS+TVHLrZR/QwaegYxpOlYyV9u9XPKOw0+QfKK3Pt/K7N6kTDXrdEUh
R1/z+moAr25RCtaQr0wl3VpZedOxfS/4tlNKypvh6Q8NbiuozqrJfIcB+MDxYOptcHYvLIdioxWt
7RNU4NRtPrevtyyk6Z8cZ+R1kOuhbAA5NB34cJ6ANg+2p0SGDBSO8v1sB7er9kKj4xFJWGvSX/xl
F016vUr+e4di7yhBjWVlintcsQ+X8Im4FtMYHAjWZ3mMtBAMHTWDBM74mND4TqxGxQlJrM3VavKU
QvkKySY2gh5++CymD6o+7EbIguTIuSTnlXC0Xv2ZaLUIhaXToV0ioyY/pbywUbTlqeU4iEoBOXrz
1AYmoixA5dM3srJTksq8CD8tv0+2+KFLQ85JiUpAs51sSPxSk5x9cXZpJXYl9dxf2WwaZ4mgdRmI
wboxYJd7pU6pgVICmEW9OxdCDW3joH9J0a7AGxY86cIQnFXANwVg9a+POEy0IMaOUlEr+TRoeVe9
7i00AIm1xT9SY/MWW23g4MSCCgSCTakCkLF5OFAVmP8459P0BtouoyucJn473EuafS2PZ8y3HndL
t5IKMXQy5YIKVXza/S+rLeTJ5+Q5ELbeeI5dmtBnhR4crJGJZNKNhv2ZX6pPD6s8UVEirQmxnpK1
R2pow/ipueoo/+gxI6CVycKnFT9dfKWzA10ZmZibGVw5OIorF+oaVpQpYdzGr/dboJ7MM2rGOcuI
fjkcfBU2FPwg/Z0FidOdrBnVeEnVm9kHGszEQSXTGainxdbmbx2XP1pTXlkJ1w5VKIMTkbWHUd9+
YGXRk1kv815GgmB2O1WNk61QtsY+b9FGokNWXSNyKWEaPJ1qeZT2/4SBFy1Vlm1kSL3Bgvg+vDoQ
Q37diUJmpO7xbJCWTrLd6tiPYHE8jgbnGNi1x9d5HUBweRqa4A+ZS/ekKJgdmiwMOfmdcgFitr2C
tsIDqvktV3x9AWK2dsXVrgsSN75lGOp8F8MDfgdqHHUwfGRjyaBq0+dd3hfmBaze6lFZ5WdNzNJJ
7Tq2szcV87SWVmK/HaDIV8hdeJN/lH91xDv+vV9yWEe0WTfF040tBb6zddJ5l2kVIme88qgoBfzw
xbVwd+tDC9vFQATwYJBI2Ni4rtRwiIyWtKOxzq0jDtZ9GsygZU7FCoZQFK6KjTSQur2NMcHn7DTH
Vo8PAIP7/PMRxgmP9IwTU1pqcofSOMiH90GsscyG+fq0Mk/r9XaCtm3t378mQe4VjGGIAi5Y8dWk
jNzi65Amb/uqtXaa0TN92LKUaGqvynJyCkH/vugBh0W1VgpFkaGDd2fu+JwSAwCAMa/nhchmUNzn
8yi+DttU7pO8N1EXFIzzlG3NWZluko5toy9WVoDOtscVrygkMdrNDbtL4kjaySVKJMRjSvl2/TBP
/3e7c9jw2RmVs/OwjrXXXjfDdGS1kKKYIHQ7yglO8doZgWvmZGp2ThBlrVybXtNqpwJrTh1RlLr8
eiB+yUkLBczwIb1g559xA+6DwI93v2BRnIbtzlKFAJYO8wIx51sJ0WUTdiizHe2pctZAJLr6eJfo
Xy9ASI8DWuiOp4UeWZ8cRGvE2ZE/AlOFNyc70dZtHyfdVz+hOvGKilGo2pHUi75ZPVrv+bJGmKhN
TtSLBQbV6n56JWwAsopXfXWNmMp8Bnxu1Ff5vachDXa2CaoYqU55oUeKIbeZV65QX8JEJid8Ox7o
R1QvHd11gHzwdFlrm+H2MKcBnYbnX6gqWu5MwJwMhMYeHPXZztqYgIeE4NVG3kqwR7j4aGBtDzAt
QfaQcA/SLK0ixdzDZvv7lZAr8k84z4f0dorX5S9y6S8b8xD2CWZFarOju/4mIKz2mk2mHRWeu8JK
jPRZI0jVsHyZhovAjEbNV4L+x8br5yGkq3D0yohvPwAY9eSeEfqTPTaa0ptsoIMJGyLEMOqj5NSN
IG/c/rdrqWYzMP8gL+atcvAJFlnerV61D97W86CKMol7GMvXEkKaZBMncnFg8UzDnjyaEldYIJ5Y
JPJJJjsgI8XKIDGsy660UKJTUduLIPevhhEktY7SD0ZHNYU9LGjACd62Ql+F23KEwv5jhp8mlNpp
Ak8yy3biH12xT2LcDE2x1aM7xrqH4L6ZnxtA44sNnJ/L8W+gaAOl7VqabCxefrPcdPa/7fG8KuW/
hfj4AEf8UF3hk9iP/Eve1wRE5tbdKtitkm68jy/ZamCX0rM6khulRkw/JyoBgd3EcbuCiMNXDBbF
B18VWfX8dyz7wqlXOThNCxyN/AerPPzC6kv/nOFQRvP1+WwVO+AcTd2Q8cUGZdEDoKpWqzmobvYv
UJ0uJ5RIFLkuDeZs2avcnI5WSKOohjdHdxcTEx0vOd9YqrcGeb4CgmJLPq/U6Z59Hi9biYlbBjVc
fpYkG6CnvVbxX3wQMpnlK0xMKlF47N5ArBmNGqzzL9RbvJ0vngDFpXxJKPNheefW9CJlr5XqoITw
Fq8WSGT8XZK3NKSq6erDzMA+2GhnfWPBunhdr6H+vksHk8YiPDbBlHZ5gXsj2WG0bKEq10xDsYne
VupoI6cFFaWyq5pKspjtMkl1Du2A86JtE3AvqXFYwVCf/HweCbbWPFrc2ptBGrZQlGDX3UrBbJ5R
3iaflunlsdgPibyoZbK+SEcu8povs81vQE35+WcfBQs6loZ2NOOXwhDTO4RheiytV2uuypaD4RdU
qtzP6DP7TsJgAsZ5RS5VeMj0Luags6EAF5c1WWkVPbmbHB/t8fTDvQ32pxprODfpJdDN182e48Pz
IZK7WGE3o/0zFtDbOD+Le+l9yfSm+F1mjuB0ptsc+L8xtczjOwKX/xkhxrtK0eWVRndAGN5Fyale
IjO/UEnmnSb86SwzUpaXJu0I694bqIxYWVrZAV58JjqWf24E2MEcjSHKSCJic7cy7M0oQh2LYD27
UtwQYkwzNACvL6HgPrgQfblyqa458YDfM8lFnYdm5+/pB3phThvfSja7BvPwR5BhImReqMNTkMFb
nG1TJoHcDCj1WpuBnHbmlZn1KIxPCDxuHkSyfUnoSGC8evxmAm2RDGVzg8AGnrD0SogVmm4hzOA7
ziOlow/3uXZgB2gGBqk7PRPLJX4Yw5q52Jm0TPAILLCbqmezdum31XsigMTt1EflyHDsx+o+tYrS
o7ZQ5Svt0BE18PFo244umC9ksFDPR1d3lIFjlbv/u7x6PSQbwAaEUcL+bkg+HRci6VsuR0R3gt+H
JhELJOTu1Q2Kixx89H6ENw8J2HYVys+VIVGi0AOpXICW5YIEIfmvzJxgAll3RVFs5nNh4SwAYeeg
S10QPQQbtXNi6ZKS6Sju0dCZYXAjntjAea2VRv+L76Wb9XZ+SutM5bnV/1PUKrNeQcBw8WDkA8In
AmAFB+i6zLypw2Gef13fg9v6llee0wmSCmF3K6ArojmLbqs5pCYuTLgsvnASUWpvIJkV0KBlj9/A
tDtdMArrUxVQBpvCQ06Oyb/lMx+1MDcrS5tlOds7ka4iNtmANiM6eUGk4pbbi8kH5e0kYJfKOBNu
iEDRfnADbfgHd7su1cHJXse6hk7oAq8mokuNiT+BTWUofT26bITvWjF5Z+cVJVsQ/w+UKropOj/k
Qzr+xdH+tqa1m6Yzxhvu1gqsrp+gXfC0Dg+1QykgmzEJ8VjStYa+IWkhlnvWoW81xWWk0WJHm+ra
2MzbQDo2tt63hT2+EmDNuP7BbcxAMTHKZQwNATptP6Tp6LX/Jy34D3Bqv1X7xqEGkCD4culaAgva
H4A4qOi8ct3b9687amTT1oQ8RhYFa49NSLydDq7igGJK7WM1ug1v4z4olpyuQJwpVUd3dZvelmWD
3uTZZ7lK+9W80Ev9Fdp3qq6D/zfZUjbkDlfxPooO2laR8NN6kK3g6AZtIBsBCYTNhpOGF+Tv9dzV
diTHyZwyUHnwQPDUy31AteEHEUsLWrPduwyhOgNDSyxLw2AOuRJD32N0VT5fhAybOfQNnd+7JOzF
QYRWjo9fWq/NiEtOmtjtEirrAr9c/Y3TA/riLmLSqmcryRhuFNVsWCeWCUMIH3SLjTtuhpBtqOX+
0kYiwhl8N3sRv0tr6efKwBnQfeYdaC7Ees9PXyYBo21Lx73oIumponZ+YRIzfO5rInOsaF0A/XVp
3Z9WxO05IZT05KNZukXV12kYyHvYTwlwMzyrR6MoXqlXoO9Va6vYJzbPva7A9tz076prA2kqdsok
/qhe0QCaqL5XeSNyt995J/eGILNhtezZu9nS3t7iF8SjVpCuRO0bxKSFDlpYxkGfRKSmCjIBrBcu
NMRpPvlptNif1G3TB1TIBggOJ/xF9t9rcjnD5S61d1GBYOYpYGEdtcYvSZh0J5kYZGFW1Y1JaWc9
SGA+8JqGdAk6HW+pzvpGKh0cYnfJFHYVev7+hwwIRh6n3JZm3x0m77UmQ44lKDx29+7nxn4HwZV4
D+3nHcPr3kaZZek/pibrQ3x2OTPZGPhKCToaKQ/MQ9/cKtuDBEQw2VwJJB2aSRf20ZnkwC10lrpG
nj5Xl1a6BLRJQXlac7iubgW48EIgNQ4KQ/FRY/dJWZs6y3D8qsBAW69kD23awc5YyxMg4dTf247U
Z7amUgbWWTfeQRduDTiP+FCfWQ418OqO4Vo9bnuozTmCy1QMaAXfoglxMQVmu7h6wAzbFqgyO/Up
tEdBfWTvCya/FfmLvG+baIaeuJytVSZJRbPCJ+gDgRPqXOO20ArZ9QGXUfoeJKGAwEG5jLE1efmp
d7KYI3XaELsVtcQeE6qbURsrcQIkSOOhCvUyT3acpBysVqRMMls7Qgj4yPsflPYVaek3mxw+ep+o
1MOyU8bHbRqvuUNkRioBzBtPyW0sEsZerOegkhefsflcQvfiLgtRJ6xULEkUoaV7mcUoanj0rJt/
blB3MY61igENdX6A4igrDljaXHwt4ttGKrKc5qTrpGLlkJmY6dpL6XE8XjDrRT+M72JZb07J+OaO
eYEbYj+28fHla9t3qFlZDuLulTz+ptSIT5N74nI7ai2EmAZuNje/mJbxL/uhWpQbHW2x93PgXpZa
dCN4wkyr8hApZdEdC9oFkyhVOt0LqqqM+sgvUxvaDboRyXg3k7pV7sqPWTTL51rU2wstoKk27Tqw
y+oYc1D/q4RxhaI2T1g0EixAgDNk3ye04Wf28xDbVQI3rhZq1/Inak6EmRIgssRbaTeic5xj5Mh6
Ut+OQYnRTwnr+Pvcn5VLawGtQA+hPxESzQW5GjaTLXZKh2YS+nXA1bbvxy+Kb/vEmFjUSCArOBQs
dNzmuqtt05CbVpw52IAuG4Aa5CjOq//EtqEqk/voB2DBMTfbHGiXfT69sGhmGkyk3Vr//s3WVCPF
vkHZj2eCzX9GWTVzMWme2g/2K7PKkF1UM5WqaPzCkrcGsHbxSVFRIbrzlSok+QVBlzcuW6mvzEA+
17vJhLBWtAimoADpa5AfHadMeeTpd1yOg/xz5GrCLYgoHitqUszzlLECjfASD+im4CItXoAdKWyC
6BaASc7vomWDFBSRsI+muLArG3wex0EfrkwpjmkdkmmgFpNSKhVRuMZp6UzYbI8cj14ss/nOoGVT
yY3Qkqlt84mu7K96U+9ie3tJYJoYzWs7I4jjJtiTDNnKeYKaRsLaYyBVPGaefXuL8s8ndDQHglHl
GRbhNMocADa5UyZ5RQFf0dipiPkLuGlwB70vtjYE6jvxH+Yy3ynrngqKWrMwOgZVA0yMAOPOPg7Z
Zw+Om/r/MSqPxjx4rhRKrlSmi4LHFwINaqW04NVaglHG+tXn8cV61EghQBb7EdSFMQ1V9Q4GUe6F
t7AXIpULsrsf6zhHv7vn2zgR5iPVBa7KSFwKjqraWckJWXqZB56OzCIHSb2pL3LO7ogLeveKjgO6
Z9pdG98Z/H3CyGpCd7HyaLGKc/0eUFETMtNqyXEwb2sgO0iVBWIYL12eNCM37nnCTRC2TnhSOmsS
6fHe/ykL4NOmbUt/8ULnJPFZ/Zdt+pcSgvmYHCD3zUldWi5OuvHFOL99up+En3waCcWFn+5EqMDz
TIL9epXE5TeAid+DMqEdCbnXVgUnfMiKM+QdJFs4mLCfEuslFiafvrD9Koq70d1RDL5NrKzEqZdd
e/7o8AhFljxlAv8wGdkQyqrK8YdE0o8A1meQcBzfpNe+nO3xp5noZ3uvcLWHwoAUlXlRJLrerSBK
Um46Nq/1WTCmOSVM7tp7oQJ0Wk3P3SfXW9toap1etbNQ22EWgB17c8wqJTLRQOsniwARE9+8ewAs
1izhDPSwLPP0D2x5hf2TJ42V1moLcVQVjlprIvEtWiVLVgz3wXVIYnVyo3x8D+zSejbsvLk3CLoa
vujY/Kq7xVhMYtJMijDF49Zah3GP0KkwvPa0pQt/fAPdIIw1h39IqqSTGveL6Y5GU+tx0rdm6+bO
ZaaJFPOFhfh9CoLrob4XdRmLJC3AdgVb7yk2V2fxPswXeGth86219p4Exp7gceOKNyAccXdhRfXr
QKqJ5jwKWwYD9t4p3tONKC7c/HwRM0c8wM+Ry+/9lvfoSOmJrKFDGh3mAi80Aq2xy0rjlqFWM07f
BVUkRelu+Pz8sAEm1fkK7p+5QV1wnVLxFEaPWGXkgItDNOAAK1gQdJKOmUjL5tQJgOMla8bduvBU
7YQDfkGJZ/YDtWv7muUvSgcofxCdYHB4mYGb98+DKkv4DLKAwATt9F5p94sVxvyBCqjW2OsMlSWk
+m06BCLdwRXRJMujLKuhVvpiovPDoTqxBB30M+1gFhMmnlRAgkl9coUJlzv7453BSeXlpNPLvVU/
lH9bhhP3ItnXZtXEa8zNq3fewfOmQaW96IpYM9L7/SpsHHbh2ZHDhH4HCwuRKdy5d0xDS6J39VfZ
wiSjWH0ppVSzzAGdk9/ucjIE4BSy5ld9IIy3CYCzt1U8BSKQ3T/QtsaS2F3L3c/Xw4iOffc2vcmJ
5JPsbJxs1Sqgg19ZBiSUWGywMeUpr44A0PE4fOAgnWxZ0S3oOwgfkKRw2fydHEjNq0lM2eBd68kJ
7uLCwUPbRaTi5bL6alyz2qr4qFR2aIikvU94we5fwGRndpCn1RQkGir3mP2jQnKNS2ys3RM63ELk
xMCOxXHNn0agLh3+VWihZcNL8wKnWuZxNv+SNg/PzXH3KgGWJO8wldJoP7WumoH2i4gNg4ue8FUi
kwxI2HZ0eL/H5/Fxr63g6evVINCpIDY8NBg9fJEOgPmzEOwav9G8hR1PX8nGxAOfcyH2rP++tWYk
FSlaAnqxwo1HKW6GLjJfPB5rhE0RqiuSZgcY2Hcl6i+dHtDs7SF22ixNZqBS1E3ZiolezIMqd5Gk
TbqyVENrTB245uzJHUsIX1I6mH6Tux6J/H6dFybu4YAymQNxAiMyRSzHQOgAoggtRm6Onuiv6o2u
5y8BE4M4MYP4CHVoQytuws4pcBXYC+4GHJHZGkiKdFMjKDKd7jC8qUc6wJ7G33ZHSrS4ZadCfSnm
Mlj18MAzSaT4Y3yjSlv2V4M0zZjE+MEKfCjlQ2s9dfKjWCEha2nlD1HAZuIqa9s95Grr4SB/43iV
lM5mnr7X9tmcTxsUXDmEgSs94gJR/M2f2rr8TuoWUjuMjbc6GW2ft/99Ef9ygVNRZ46Rk1ZczXRq
XC0xduovQn8NVlrdSoird5oZdwp8N+LxvR4eYW/c5Y6RSKI4EhSKYx+amQGI5CXVOki97M8KRVXT
BfInD1qSNPmGoBBDWd7NZp11gRUiyX9dacFAM8lH9FS6hmdFKjdrmaN8jerlvJgXtl7Ai4q5I8sv
qTTkVaZNU2h+vP9O2Ll2gTJiuYcKYW/Ejk6IKnsw2u9Lwqq4W+QyQ41scPAQfN+AxmC6+9Yy6a/l
JHV0nfGEc3fBvWA49dNRtQqFbDKE8jLvLqvzHxfS4Q9WkwY7e54o3V8AZGPX1NWpLdoDuSibzeFJ
SzecYT684KEyDr0PlnxgKYiROla1MO496/UEHFH/2eBGmGl31muaUd5OIecXH5zIU78uK9SU9YBu
TLuJaHNuHh/HjXXEX+nzzMZS2KdrGGu1zBxW6BHFIZb/x3Xi1fRnKiduPgiZvENQm7jqfHxrdTxC
ZgDNex8XQnhm/0dvY2RpMn6c5FPN49cbNRv+hLS0BQfhWE06vRfWFVFlaQhM2SbvRJKnXgFk8miz
X8l1w1usYPYlGjnZ4ioDCTNDGrHK2qt6VDJXzbwLpctyPpLRoQlo9Eg6rPC55hh7UdfsojGGrIwj
wVWWaZdpnSW4/q2zd/DjH8jkDq0VcsBtom122cVGphgpjj6yEVWUpxhkI03r2nbrNJGy6yXIHWTS
kYbv54BYnnp9mWOMyedH0CkdIUzI1HK252rXu4Cb2hl0fl0dfAGEOuwK99SXZUuBv1iaUtMlH+TO
WbEkwN5epEuU/5UhLrOHXrKMAUW9/gyOUk46XC2zBeTXFZrcRvbk3zsANhmqqsy8IV+gfbh3Ym20
F/E8BKZW2Pjnz/BEoX6/CtCRr//6QzHkTFyRCApk+N47I3nv2KvLCc8VAB0EX09UZrBzHHDFB+6F
BqEOj4JjiHBsTAVsWmVu2bfxpr2TMrScGrjWpeDZlfFOZi2+O8ZssBcPduRNpUYKEPFMopzlWUOE
77gZtKyrqzh+ILFv8vtrREk5RqlWjuS7DT1ZfXZmuZ4qoQFM72oKw33UwEionNG1+yIRSYonc9KB
qTxtpgGFbWURBL/fJ5cHtW9Ni2pb/qb6zB9aTJ94qEElw5Ltvl8aqeU3+qsYe+4flnEDRJ6OWtWE
Dw9RdHxk62GbmCKq6Qa9BHl/EVN460AZKk0rohP21KSAO0KWolE4euzVAJg/JGzdhSBGtRzV0unP
7InrwuFDqxOvyFzXOkeqQTMx+WKF1xdtt34CTnVsidOsy/kzu5aKbaBwIgpm5aq5PPgxZimN+9RQ
tf10dJE2VgdLiK2KhHpUuwQaHVYRHjnjtpFnY5gkLcL6LbkVXDdaLbn9RGUPUpj8gybr0besJDyM
V8cyOf5CTB+yKYo8Sx7BKQ+W8BlNPTX2Ia9GgVfkc5qm32cH170HFJDwrnBjqAQD3Ao6604+rene
n/LDguV6OmLC6bE/1zkeBsiHa1Lv1wl2O1FSDpSglCSjrnoASQO55aIcGDSa0bfb7vBXTY5eWAaQ
d20XanEP6Im/icoIRLsmR0u0MaaJXiv1CBvM5+RscJA/OxsPLAGxUe/ACAy+Z0oO59D2gsfUQFGk
GrSWV1k3gl0P8LeK6YwHvmZhlCACuoDnjrYFrvwU2rfG1o49O4xuDoltsGPaeM8gfK3enkZkgl7B
unb7vHgoFmdQCISpd/4+y6zd46FCO+SexgPMCH61a/5xPiXIOLG4082hWFj4becDK1bqD3RJ31uq
i/rqESXGgQ2FaidSTxRLum4axYami5+BJCIrtJb7aM1BHCdo3iTLn6F25FJLhbfiAHix8b+wuri4
S4NQyI28zBpyTrc9lOUqZ0yZ5WcmY8L3IN3W5sEO9IS/q79GAZTxGQcZZHPwrnmG6qY+NW7kDfOl
qkQsLCwgQnJIIoGvylMm8zzlEhBU3DxcVeBKX0wRY4+LgXI4tSc79lQRVtwz5jzkUnrUwiUzH77a
mApGf0fgiheuHMx3gRDaxY8a9DIYbtH+udS4Nxv93cWobGftw0701UgrpmUxnDFUHxzb9ixUllBT
n3VD92j7IOzcwavn2Y2XPrg9nGChi51zNLldDRRXIcXfflIgDw/7oigUpGByN//Hj7CqgiI/kZF+
3E1VAa2ZFIKkpJEu+JNFpClVRugt5GA6PsCh6OiBRcAi1R74vIPBVQeplV5td1lVDf/7cM0pTd25
L3SV9KtAL9/S19Ui5d//W2wqP6w4U5Mv/ifL/FpJIuSW05IVlpJjMCIvLgkonyVIzK7qW/HF4x8L
ERPWv3JlW1WryF9AoBCMRsBy/zGGr2gYQqY0BwCI1kadzHWYOiHRWAGwm6KJYP1royOEf60SMZjo
h4qcrLEMY62wcAXqDwew5FFSUAXc8pRHLAcmDDZecxUuyEQnG+mdniV2w7iHTyGQOOHp1eEOvFEl
rnNivIv601p0UYhf30mf01FUrA0vFQmmbJFXVexjJ89hUzJYUMxg2Qzp35/3Xk+gIwQuT8Vo11DW
5U541dhr1jWVT4r8YmYdsiySaA9RUZiTFWQri1BG1YC9su16EVCnNtP84+uzHlmzmnQW5wZR72CP
Cu48/Fphtm8rsqiDjBhcubcS7oXTOW2xaPbEkFrLUy7aSgPeJONV0VX32kA1s9/tOfAjSb3eYlJS
tZDp5+2wbwHW8xESYj/Zz7jypA5PKBl7LV4cwNaIvQYMcxrtoL2m39zvx6Jz/ALeWb6Lr9mJdLQM
a+eORDyB2Qh5EIu+kvVKLV9E1xMFFgIx0cmjk55ccGXvQ0+JI7KzK+WMAOVaPDvec8liOh9xqL36
XFB3tSLah4iwyU9ZaceWMPjffV0qg/b62C+S2rAg7Wfw5stcrFtQ/HhbuvC/ktO1ReYOjXQL7CpS
jBd+gPLwFw+iu/vV6Fau7UObe5RlfrJuWEzNx4BPVj05BuicocDljS5pa2ni02+f4na/8WIu22N1
BpE63YpcBkcd9BLW6B8/z8UbLTm9A+uE0hkAqLYU5bo3EnthxZU0X41NBa1AKyCKdkll/hBcabXI
qgZjtxVSDwIoqRF1oG8Dh358EcD5ZyL8TAvCPrcXse5g0wUp7VAuFH+J4viouq0LV08SuvQaExiQ
kXKkkkmz/HSulFeqxdsAHWezwyzHn0NFHhQlsDaXoSn7aJBmh30UkQ3hNDuuvDosHWLE/Ei4AUfD
PZ/KU5zqS8zaaNO4+PtNmd0CYZDop2Up/rdZ2b8hWOJwVlYE2H8+EPUzvgcWbId0bFfG0rnRw8yF
bH1mCadMdq3nQ1c7sPuZaO/BkJzDX6qkz7KTTOmVyhyuCYDWQU0LirBDFd6uxmacAbLZWcTbmBMM
in9lRukSw0QYWyTcxMlDwKD1gWhnlCqayPDjI3h+sTHu+ukbNnctTPJArkYVZzjRO15wWNerXCBN
z0v2Vv9KOlaJp9SVFlmtJs3sDR+ddHSgKIpxI9lQfa46LbEdnTIL2U37g5i6usAS7mFVf8Vi2egI
xd6kaE9g3kuC1lui005g4duqOzdo0Sfo9FGjoPaDpWDwz5xd3ffnpTYVzE1Jonqg25ArugAzXuSg
cGKuUZ+yBQS9R358rdlY43hgYFPAYhfcXSQ48BeclZ6dLZO25lEjC4Z0DZBuJCyhOHEBAedq6Vt/
WIzrj3N2hIGNfgNn2RaRM06Z0leuBvuTIvtrGWpTJ+3OGpsZ9LVeXMQEELgEjO7ep90IGMLEcUl+
5eWGgG9V2dlP33yHtd+0YTYcN7WpY+uBGK4Qx/pWYMdAdF/1/BNn6VzXIYJ3wxEqHklQQXlZ/N1u
DdHuYm5+YRjymxBhXzIZ9cXGZu41E/t8L4oOpIDdForDwjEstj0rkOXdSezMkUUR1eaG7R4DoI84
FpahPj8BaDn33LPeQX+0kw50/lCdkyu3tSAuLvhbnfeNqUy+z0yYsmyIGj5NaggGpFuctBp3XxBU
wKaw+Vjo1WdGeIz55PCaXLTST4GPkZkP5zGVKM7x0Yn+/2yE5XyoL0Om1o5/HSDBVC4ohNE+r9KN
aX6En936/ScXioRJu+hI2TZFDGg1N6Ljoq62y6fxvtsJqGKN1mHlW50i8S6opvmj87LlHrr56hF3
0tGtXtwWDv9ESkHBT5tPZJKJMY0dj5+DDgGwtKpkqINzqJN99pCua8lPGwy8swQ4c8jPx2RDkTxs
jrTBXglq50Qgf4zMRaeoeWC1YWU+vnH9VdmqdicUp6xvfAainOGwDNqS3QCK37t4Rg1h0mXbVX8L
utaGyHBGunw+09wCy+upWL0h8z+ItvAX4g9XM0yB+JSMvfOfWUtzgy+dX3UZ/1K2uE3s/1QBFRiH
oJsufrC0q8UZ90+7XwUBbrVSAfNRfaHY1omCsMcckrWBbDT6HZxhjo2xi/V8gcyNhrgYTOPkVb8E
+XrH3aPsyT6XLVBpu0io9ZBezfO2Pa1IjbJbpBFalrUZnFu9Lbxz0mW4QTISOMg4Nsed+osc+5ax
4GWMoSxYUMb5JqwHoOd23dhqZzeAuSk2gF2EAH7pZ/trwbJT5JDYGUKND199Zoj8DxQye3AxX4oZ
PilVOk+oG3XmiFEyekLKvVcq7cn4acYHDvUx7wCXH3sxEriOvtYrsfPdF/bXDEeCCAe84mXBo4nA
7XRuo3YhJ+ZXY2LGsHGlxwdCtYi+SUjVGZkMoSYR/t8OcEowCiMIilKwRrnmv9JZ/sg2c9rOrzV2
Wu1TTt3AdAMlOCpOZFmNCZlNhnkGYdJCnuKHeEr+I2y8gUnPQk0bPxiRDnjhJsT5YxzvEUTXujTb
7bW50u20uaUsse+3qIeCyOfxQ9vleytoK1y0GXVi805Bi8w+8KxtAEzSdSi31EEJsRsN7NgdA1s8
1CoNbKj02XYZ/7uvYMOsbNJGmsNxWb5936qn1vSWbJlj9BE07RXRH6e410+lFVkfxLTNOS/5j/Uq
H+i8UaRv4ayihahazBgmtZXsOg0W8TjzrGMLOXYLuCz8b7nQOFDJKaJjZ4Vda/9tpntvuB6ePh9+
wtKuW60PPfAD7TDXOuNVZ7OyyEXvQkWCqbepi+JpLHFYd19WuKmva7R2i6/3bzd/hR3obkaEhpHT
Sx8W4dy6Gr+R/9TaJGWROO0wfNSdjLTS9jegYkzrLqyKd3NXa5mzgFJZQsBh77lCw0ihmk/4gZPP
jPk0r5/t3zDB6n6tWyG2fI/2DYkr0byJweacfpM8o36H+IbHq4tSth0rSF5xky9oQanGwRuAQ2gf
oE4LaqrssNdzU0P32JctXzBI2cCVI+mMkPK7vK/ysVU2jojInoHfqzlhiwUu12uqFNo8OcgGvbgZ
nRPY2U5fELtFsD/riB4gOrRYdbLyovULXH+mwfP6ZObP9yyhWT97aLXthuIWgAfiLROtUBpFQq/1
Ux00+O3uqXzFvf91RIoQirBDGFZGkF8knZ+zzyVkND2b3Lb9SiMqqXum9OOXp8rsI6nvTTEmjyMZ
5D6KJVPf6xt/ISXrdfJ9RYL/iH0+VWbDw0JaeL3INTQ/3J3E4pRUNewDgxjNGlEkkxbDSL3fa1im
VUUo79/JrifgYMr6+UIm92QGfzserK0bUn8ukYSSPfV9PSivh2n6PtYi7jQat6okLihjE5PSXLvc
3wBrPssaEA0Gcl1IMaD4ndEg6YTsErb421kzGnrXwZP5B1ax3gS1agc+PbwACnD5U03kKCWxCHD4
mRYdenuQ2aawBBPeKTY+V331bfTj3V8OhhNzfyYvllrL4tc+m9XFd1v2dxXGqfVQTKK7tZxUPoaE
BpP/JkTN0vl9ocHIp57wpX1jms43MM2XOOkMBulF4iNxSMvF38ySOR84f//EFFXYciqC5jHWKHO6
TIyJoxdk/YlqFem93C+mkoVJZBsKjjTgUnfOI+ZJxyaTw0Hf5C/fJjoqXDDzvafdm6dKwYILYczR
mMfmaqnSowlxDDP6SDe1ya3U+q67ro8MLcpIs8JsNIsvs6D4kJKwGo+l3xrzS54xLzWX1loOHRwH
iPoKRgjjFVjnX4cjbaPgoxltcVcPtVNdm+4gKNA1KscPtlV4YRDCalVUQffzGWVqGlHOiVjStW2K
eRogJ7Hb3/uvVi0lJgH1RYnJuZSr3KEaZIRV46HcBxG4/bU8eOEYFwnuI5U8vaCCbxxJ5Q3mLqoo
lc/2Fb6clKgV0jXzrmX4fkfC2H2Nk6B/BTCzgI+AxoZc0+hwa8cZIjmSqskaK8lYRw71uwUuGc7z
VAj61mdMkN4cuO7BjWXpLTeoOLjZrLaWjydYyPHOwpM2HfGiqRZCi3nkp04WEeckGVU1Yvcu8tKk
uW8ryuCTnextbHOAsF6fpyGQ2OF6F3q/oyXignmSie0kU3byoui0kJSxKrU/SglYnep/G0ZT//Qi
YH8R89lluN3mUn9DW27KelEMWmw50q/2JTfV8ak9eMj9UIQ5Nr5H7SOHmSqdGJ3xEL+Q8qE8DD+E
bVz2YUR81mS+0798xaXR69/2+LH0zupNhI5HeRhfnPNqlzkgcHzGJsnhwWw8YhicxufXA/iVYsRm
C8gdzWHJ5m84xsl/tW0enibN/kLGaJv5yJfA6JXzNBaywxbEhMeURR34p2ZGqKNvtBOVc3e2cWGY
B+BekEOpOW+kxp1a7xMhaFgGx0nL3DyHp5EDyEmN0Ukmu+WPwJ5wzQZaLvbSMsayF8PTW/9ThtQc
fU1JD5dOvOyLq3YSpHtMweYtIAGDMEOUrbJDD7Z6K7GQjhqXAl4BTmN45MMWorsCY65VT12zqSFk
rzrnAeDnBvezswNoVWYoOj2kUysrrR3ssv1YpHI1qcaDVgWat0FS61kouauyvUNGapTxrLvTgDRO
v+A/6qO1MK1Jn9aOG1ZmmQan/37ScTJN16mTvC4Gw5Vfayq0SbWqYero2BbjRshXecOo4NaOOLhg
0NNlsQzTIhMwlmOaqbsanFOGP0M5EMUrfGfMsIeUW5yQLfhcn/oTZsdUGHOlr5m/qoWQis9RTPgt
mqm1GztTXfNe/dZYH/gsDIDxV79qM6zu3h1EPl3bVsNszwmWD0qe0bCKMoWdjUwc7zicKkbzt5HX
C7srM7caCr/OyZC1biLjERJwwPvSE2O+SO5/UATObcN/aktQi4F+Nh+oe9tpXQcoZNwmAZ7SXc95
KDxeE3+LOoMLG0evS1tzpH2DtUjme3xaiQoZJuqYfC2nwa+sHF1+3WMunICG0LeVKAf8NfrxbJ1G
wwIuSZUQFeHf0pntt3obFus8aTRH2yRT4aIRsdfeHAPA5hxCA6ayLPQKIZUk5/ANVRsPJSOGNp84
mrIF9SglzuU3Aq14G6e+6XCg41yQVQrIxU/efdcYS+dYPLiDM+UNEVAkMO6VxxBynzAS1J5KwEWb
sihS9cg/4wHNy4J/x9zMaOX5EFGzcjsqxxIEsGIxvycO7Oaduxt6RS2Dfa9/sJ3VXe6lkxaZ204S
1khbHS/vRYexM5ksbOwyEeK39oGudWuL9i+E+975Jlv/yFnbFZ96bF7Ja5TPt6Q0sJVZQwcskSlc
ev212Sk0djag1rZycuYkj/OJ2TOs3KuMVRTooR2woIIRDH0x0oKsJRVltCrJnSlufEwwhlBclang
r3BSRaMSUcYz7MSiaAPux1RqohiNP9OA35CQ/sbvDl+2+DVIzBN/AfdkzzpyIJfCnxeh+hnkc0tB
c8QG1pNzq89K0BDbemmM2nNCuxzqiHaAmlZe87Glec48feFuoHu5XI3o8ngaxWVQxNDxlwTKic8r
K6Ub0Z2wIBYfs40amEU7w6c60/iCsITeGsnRXhEKBjHkeGgeVKAXvVl2r4Xj5ZAKA0phWrL0ZRI5
7fQDyn2/rlxyNN1vcofufQ67LPu4qZZ0/3nb+mAUFVKvOiMZ6ZghsCKnU7Fm7Mr2/FPaGugHSxgH
9z2/2UzNt3Xm12BwCTQYC9cyJ763crqGlhjqKUN/puQaM9pMg+66JH+FBzuBHrd3qTdvt1dQqGlF
lOxTf5D2RLV9x1rIWr+yxFdXDbAxGK9cxXCo0DW9jIEwTQZ3AoshTvef6XYUNik+N0eWAxmrZvau
4pY1pQ00xUHFzB90jASAhtz1ILhX3dsNvDaEHrbv0FS/T1RIXLGr59wf2HLn08/Io6zUaj5QM/Lk
OPANZD9LbIyKDqnzmZVyp39/uB48NU1dMKjl8fHom4eajL9Su19O0O3of98uRiHbvenEvCyBWhfi
+L5/AFGZe5ixYyG7YmbOJh+YHWV+8G6cOHGfWZvMFJprPWK5F5/o5PFlf/cIqTakVO13fQNp/Aoe
ZMZTBejRM32uC5mRRPbuL8eW374zGgYerPBXqv5r4bfxZHdgxKVEVswqUyMWe4oovFuOpIE2m9l9
26BI+fy6BNiQaC9yIC9que35bBZa8RjAG+HMqjyyEAhmGQsVTO22RgfK3lWA2bBh5sqk7AfMN5+e
/voZwsV4ntMZfsgINAGLv9nBVTTpt4VXLrxQaGNDes+Lvcr8oG++hQVXATr3WezezOS9fJjiIFcG
VikPoNBaO3rlbQhf7phrHexinVm85mPx7L0OJLpOusS9cx/Wm61Y1ntYehqv/0EVuG7RmKPyguA/
cuxpNRl5O06l7guY3dn7NPZJeknL0DNqOfpKxP4D67Yiz0iDG4e59xOO1KQoI+3xfwJVKFR5lwQI
iSIY+t6v5L0sDdJ+6kngpLdEwQHsC3QgQiYWiScniJf7BcGRHdyLJ1yjmQaiLvnxnXjBz0vi+3bF
cbt697TvJrinfMA8PIcBkzk0acqv1lP2/jjn0EH8sWgbS7qfD6i4aZYKWBbFmf6JSAUghCEtCjWW
SfMXNby3Cod2GpcOJM0I1Y6/H07pVT8NruzOz7bF+qY2jVgKE9csX4TvYxkU2/iD7DX+8WFQ5YnK
SCqVTB+ZQB36e903nl7yLMEFfgwn0R4QLCGGlr75NDmAj3vyl5ZLpm4ehNRpkmPu6pp2iVIZhw7w
WSTR01XDGNAWjyk+jtZVwRsm4cgwU9yu+Uu5E/Z+3bWmZQCila2Xl7N/fnhwhISYzMgwKkb3OHQ8
yrr5UfrAB7upNzLBbVk564fo/aYnwu6sMXLO1rwlZDQeiNDAyVTd4JJRF/4NLOBL39l4qHdf4JTD
UfIiDpjDbs4ZdA1larnQAtlfRfrACdKkrEp3qCgNCM2Mbk0y9b2jlVyJ3AqTOdTvzQjcqsWkYaVG
1gxvGpgLNwTMChAx2J+K6e5t+KyrBxQvP4XtMedTRJcYrGadHdGSpxtOme153DFuPZJpxDg+JnIu
zXEFeyeIlPSVl4DeVIut1ND1ogzcnioYOCqSkPdfuEO/3mtv3UkkhgUcoG3drffTnjrD94uZWmBO
LOn0f2opD0t/GdkrWgmt51cxnNphiRRAXspI0p57lNet0Coo68mIvdhkz4fQNwpm1MzDw7jpWlt9
m/eFdJPIdE/VqN+kv0viO+pjm/wwlwag5WNYd/G9rO50SKakV9IABpkoVsrQuFOusw4ELfM+UY76
FqkhvK4J/vy48yqo4Wtl0FcLNOzTs0yJkxEqtuUSgVKWFYk5UVUAyeETAqXrqIIOtK1rhhMkc27N
IRjl4ffc3KtJ4LxmgX8xnu76MA7R4XTye1wl8IGaMUBjezSdAEo+qGHXMkbH8muqcXFw+erhB/3c
+Zg/AoqOc6ZFfAm5t7Z3PNaTLEH1crpgJJJ+1uvo1nCWbUGhZgj1fJvRwdgjQ/pGgbieo79WWUO/
GHMhX0HoYNoJ/SgIKik+dK9fHtnUvpGHelqzCNAlpGRWHrQ3J1tvJOrn5XNil6HdA7NVurFHPUQ3
udMCSi/6Kl+1vHz2XWHvAPcPTYwdrrfpmpcrPm8MAsXS+RGnoMsIt9yNsikWS/CAczgQsJS7rZSf
OdXAlI6HucFkdZf6/L3HhDKbhZDtkLPxvnw+PrC6AQ3MepQ391k2sQA7+db3aVPr6bq63tx6owIF
f9HBsHUlcmgW6Hgb9FzORXbIusWR/9t03qkO0stnflkt/vO/fhLxw1hUSX6rluYn3shD/ugr8TdM
PmYUvD03Z3xZDtu8Cv29jGAsLKnffk5JPm2xeF2qw32VBs/+N5VNT8EHw2i3MIrA86V5PCAs7oRX
oaTEARkC/20xzW2VVzkWhI9m7rHd2WEGiMUEnr1Jla8uxjg6jRKd6rrQ0Q865yFzipjv6SDuMM8V
B6AgkWFqlGv9OakfnZyAMpdeRHYE7XxCVoJhFCU/L5aVCM/Yyougtlpc8EZ/nqR6udpV4NWO54MZ
gERyEIaoVw7moCy8Y2T0jLLCRymiKEAkEKft3nN6yLMQQ7NX8f/6NfGbJW4sK6vv3nY0Yip1MFEE
Jxi7QyEOQUY6L0KJWDBnmMhBsOpGudQP5BeOnPQwb1irnik9W42lJWxyYTzpYGmM4p/4DJbM4nXq
RnjWWWjCD5fDuT3OoBE+rqxlpuE3W5+MRY222q2Ttfw9xTpfncjk18vcXyx3+Trj+HF0fJtmJDvS
S/CW6zgrH+SCmlumsvPXzK2SaE3c9GiUlrKr4r35l/xfo0XS1k4731fsAioOGg4qSctqa8vRJ8b2
IAVaVJJZVp37duitZEFKi60Ham5RFzr/136HIV6bm49fqmGcb+TTogrDJ/tPWIT25R1FvxuaxU/c
BSiw8Lf2yWdTkQ0ObkXHhGOaZ/yBtxhzK5/xWOOrgQuVKQNUwsRTd3BYJxrCSwd1djgje6wYpSRs
QvLhBqhJzBbL6euR1oMOu1O0RhjiNVvaQFKAHO7/VRe3oMaRO8FVHObx7/0Y3UQ1L6AWxen7BJp2
SJbqZuKhSJPSD5UkpiSkL+F1GVFp/ht8G6XY/ICP3D+wT2Te5TuL/WiES0a+iHoIYZSb7CSYjcHB
IXnrBi3k6vcgsou/Q6gvAL/yjOzBK9h7G018xF2H+6Fx98stki8Ku/qDNLAmEzJ+ClM46oTVukqm
YZvHs3HUVUeLtg46uB62y4Z6Ix/AQDtwytr1B2jex60YdUGP4AX/+3bcyDNjVkI+wnEyCA2eKgBF
5/y4WmLXV0v7bPoFH+/+f+mkx+1IdcB6zjaTkZA9kcRJyWqia+q4e81c5iohALFMljeAj1yZFg50
ZkYqpTFOkFWKL1YzraIPKShbrF6yZAYsPjWyFjrSqKOXQgpeu+tXpWsmrynNeYl/Q9ESWnxUuYkY
cEqiFR7BH9bIjIXeXj1iAnw2Xw7oPFCOg7PNTsNL5oEsBFmZ595IK54sxGHO+o5xbv2dUhViv5S9
jXfqF2YSV7jtzXjs/IYyHrXw7WWmI8voLmwr75PENS7CHB9IPcJ1HUkCVaLdAuz8RGryQATr9nK/
Nac2DfYb1TBPBjEPjYvCQvXaQb1Oy5PRgfThppMyAop8LhqNXycdosiCpgs/VCsjHuL1AOR9PAiL
WGuseH8w/YtFFYuUrmD3Sqie2EFoxZLzURJKFIDRUGrsIMhq8u6araIb5IsYUVt+BYFqr20d9hLa
gStBhbuFPSQO8IdLyG2hh3Qfhq1+k98uylTvtwEn/AbjWoSVrcz32oiNS0ZixWg21lwIQ8zSHqZU
qbcQfZLcsB9UP1LGbPPtb3ppOdP2M9iV7HluBd0K5RYDMpwnfJN8mWO8YdOWowj6hTmk6X8VDMt8
srFiT/D150KXtQENUx/YQD3zUEK4YpaMsD6eAXlWf6oBazGH6iQy+GutwFOHPlvqLZbfTZTmJNjt
8bc1H+BoSJWl2ngpv9/F2ctF/p2hEM8KzdfnCo0vXaxwSYGRhLW/+o+ow92utDyU9UC6++hTzTeX
nGZmpSphR3Vgnb1CR+NWnwhF14F79F1yUOZuErTQBTnhTgjDgOzaBYpHdnuYD0djSec2Z6526a9T
ZWFwv2ywipbs4CoUhGOOvSzwM1QTBQ3lGcdS86aDZTDfhL5nVnQvSL5XnSv6hxFcj5OKI9riSTh7
KZsJtGKU7mhYFmM3iBInjbCz/ECAAC+KicGBbY1ZG2Vg/WWVOhuKwCq76V9mGYLY5aaDoIpHoHen
EIWTBG2fR8f2ClFTk0dLMYQCU30DEOsrCMpSB7ieE3jdkRlbS3raLSn2RhMBDlHArOWReCsAMboe
8l+GiM78NqcPJioakKRmOzfch9GDuN62Q69bc5UtUmKWmKFyDHDlbjIFBlNZp2B8Hd2PBtpuCHlp
8pu03/e9rL3H74BVB8Z/YOQIBjxtlPE0M2DbVakyW5D09MSb+U1VFutESb0a4UvEZgPlDkvXGABJ
9iq7F5xD4NChAHC4QOIMHhy7qXH2Q/IAqTbelWpBS1fw1HB/UYsFD3v8MHFSdcjDs790juF2TuZa
X+UuT9oSBHI2MaSG3PV47CNMkIcHQrBcoVKXkRBjXySdEwyDLFDzlHXlnpZrtw6xhadYPrr+Rmpt
TZzT71cbbBKt3fvN+LOG0GTsg3H2C6gykrRKdRVRU/5VkaJf4vUiQK7wzvP+znBcAqaL6Qb+MZ+Z
rIp6r1Vj+HtyWMncmlNsqB0R01E7b5CxfBbwwYdRH8sytawIOJqSDMv908SyIblhxA8NL3MmLpie
eMaiYsR1IGBVi0dalwu1OxHD4O1qMycI5gYUh/gPgKzqntzvfglRtvbYzxNIfzN9a856rOwixFI1
epW2u6CvyQUEpgJrPtaWggAhVpCsamrQhm0Oz+/E3o1M4Igq5nyO25oUlN/JTmgRIlfefWd0xCn/
x9zkYFPzmK1YlYc/hxtgih3a7CoUYR7cS6fPyyyEwphrFeBB+ujgFqzmPd1LRP6xjpAXx4rhvLqF
nwV3RCCGypmnoPOwlpWi1zs0O27MR9WIUuXlENScT4zbrfEGVLD+P4GS/BkVJR1NwL0cgDaaITgR
xChuDH/40JYItUxXWqtTZNA+PBBQrpCgP0px1PFQRgu7/+Ga8+fxEvH9JlwFAh8HglSy8Q/0ny80
85gexV8FT50kM/J6pd+ivHz50HZnXVtxa50l3drySylk1yLtZipLgg0PN/Rx84e88lGD7Y9MM1JD
nDGl+Hbvc8wZEWjJUia9CAB0dqIoDx4UZA4gC+zshBmHgef8Nrbtjvjb4CQVG6rijrFyKsjU9yWj
vR1oCw5w6NC8XUym3iePoZS5lsaNCZooh6d/IiR3HxZdmClXSWEpZEIBDq7vcopxWyLKsvaX8Zq5
GbT1f1UVy9S6dioKZzJQnRW6MfBrX4isCQI+3PTyS4NCAAt6/eWuoL2PhEKRr0lNyEyBNNuwfB7J
Qw+da76QIG9GoaRgC5ETQk7VhE/850LdnHR7FwQLOO9Mnyq020qAqXdhk36eegooQsjY0GQ3oETh
vcAL3iQAOQk04gd5R5JfAre3DfSqWdSWOJ0xmJQQH3FDTVjqoUOk9NbGAdLwCBUB5BQOJthRs1yC
DSJxu3K+z0L+Up5LUDo3p200JlCuSCA8fzhx1OLGccD+t5GoV2o3WoXJBLSHKK/65x0eTimRKst0
htXawFi/ZRP1kRmy7zsQbIivlEMZyoH1likMytvGpM8+jPK2varCKwy5eUABlOSLUMlPg+NnbDd9
rtYhHe5FIcCpsp50GH/XT7hKj8wxqKstTFbjxZ3vfR/qGSgV+qJuE7elFgTuFA4CKoQq8dkFanZA
x9ti2zb9hoHJ67IMD1hrB0Ojjzn7/pzlgoK95ukyFjPiSuxS9Uw9ZWZsxx2ygF1iDYNFUyh1Xe2I
Zb2xb5JXry5b7YQYoSijiMxbbteG8mN6lrQ3EHikxcvGZnBUgTsz6OyU7+IMz7EsRKqd96iR/98M
NtMRW5lNsxrlTNOGHVvHcbtzyw/L1XuvpZudnDj0lST8YJwc6teS4vSNVxhJjzgqKJb2JYgwJEbs
uoM6HMWgSyO/DJBL6BQmD16M5ZeE9tiO8VYdHQMfeYjtA1CT3q1KOXvyVdi8Xn+Dj8AQe5/Pdy1/
4dRTQU+djjZwivxEGSVSHb4PrdrtRYRkEKQkz7RyzhFTS762rIq98uq6e/FpolGRY+5dL/fjic2C
0MRjR6UicL2Fgu2oMOk/QJIlVg/dsIhEbcoTBXFjOaqC43c9pMcIBImbGVKazO0P2QGQtS6ZhwqA
AN6VsxTkmQFhs7Hc0A1LRTeKeq5a/peyuEtXl8eZrY7BHqceF0xAsHkx1G7iIORV+w7DGpqW5oKU
Uothj/jyZjr7RZjFFEJRj00BWdPKo7lXJQYVknNg8NmbFDBN/JuRZX/zm57YKjVbUBmbSLuPKR+Z
Do6Wf1/0/NrE8peraITLWpdpQAnPMHAnjlB09ii0zBlFZn2buxZzHmkjj5rj8abXgn/trrXhFiuH
9DW96x1N6HK2CZNMD59yait86USpIsy/r2R6ytccGtxX/WaaRJkMQzvGcXiI7yXQL37DJianW14M
oTPTGQMEoYdVppbjldM86OiS/0oxKxSp7rm5RbyKV+s0Y5pcxNk14B8ZUK4sR+FwFUIA0KTXKnmS
KCWnxtlga/dGlrD/Ce721jpVzzjOGNWs2RHM51LomdKcde2GGF2f496vElRy9YBim9RN9p/42mD/
aQht6exAs83vhjpSmhHOGXFDZ+Mz/CoAOLr0DtZ44+G5p4Hu6f26oKrXjg/LqnQSFIAYtl0aywjI
4USU2fWKw1l9ZX+xgK1V7AupdRD6aFIyib4/GVIKnusfz4zmXEKdIb13plohas/gFTSod+hi8wzu
JrtvkKEbdh0DLvXuBwF6bXR6MwFjq/eMuqxGp4SJARMDfWhrYPzl1dgiQ36q8MEMs2cqQWspF/SF
qY1ybPv0hDiB5YcjFIZPOI6OXimymJbul1Pv7fDT+754r9CMnmJYxEnn/3dY0aWV0YsxnduUNAWU
kYcDctSbJPD92bhs6bqnOEng/j71k7Ed1h29R1E5+kYDTIKAfG0NW+58q2nR1cbP2CJgxqKKGKcM
GUwgNZ7QTq/GPrSNxWBEnSG/FqrIJjpPAlY4r1IueVSJulJzWbBThFwXrpAgxWGOVGApXt7v7vwl
dugfKrHfwrtn0+uoepu/jWPFy1FnMVoOgF/eG/JDvM8zkVcE/wy3IOlPeMZsaYcFWMwh5d96keso
NGozC+W0HBuLiHgh2Wkqms5o29S7XfCpF3G4yCQjtvNN5/+KVj74NMcSsd5/pXbMj67OBPkzoqgx
Nj4YWLdS/1muwW4QPUDpaOqnkfFH+3qIIijWMjxFdSSXewMPY4JiX4puDXkJhLyvuI3ItLoyg9Jc
vMTgAm/J+G4uq4AAD2ByKp200OhSX1FAuuvPoBvObaFbAjblPXli8VKPztIcl5Mx8Ngp7oBUyiBM
IszWv64QyeAWXtvjCn9Aslfr6sGrX/O7iQwNaeZf50lr9IVbR9LHZ2MmHgrDLfRUP9EbYx7zMnRb
pJGuwzDp2QnjjqjadGJgWqh7tXkRfEq7DaHI2nuuGs8729XKpxSHPNT2aNaTo8KyOpBE1knWK83K
6Rqh/sp730a3SOXs8IC4j3DQ4lkfS2t/y1BJh0PKZbq5ZTKjX0ZA4TGfvveX6XMYC5MAHyAPoWeE
CqRkp+4EBIsyZjZMWJ+Mk6du73XGUNznBEr+3NRA33ehl8I9a+bcN3Og83h5D++lj+qcTQwSp036
HWSucEwHJSHKCuKk9C7MkPXXv7AKyDQnWbZB1KO763EQNHU5U5kpExGnLNFK2ahH4/M2BT5o9TfW
1CchSKI1J6raQ1wjtLxub81uRlU2luEMDgWdxWntjPP9sfunEgoS4NfVipSQ+SuW4DV9MoJCTdE8
/vZoLznIPp3l+gBkM+L6W+1gQ+6GeXuUaP1MVF2loBzO/sAaAN2UZJHbSe+OLfim5MV3TMHyWg4T
6hfUjsl42qnYyVTK8bM7rQ5hiv8XbPQtmzi9FIQ7VcshCa2/nJd0h8mquPy1IQI38mOZ2L4ZvKxN
6UHfamEhiuOTuLX7jUpPqMRf7hMlK4qAEnOuWuMy4/tiR9Ey5YEH3xjfRGwpQc2FaOo4uzx3LcTi
15DZaKGZhVc2/0llTAHQnEwAYq6jNqDtGYneyg5ekvwqSyc/W56LjSM0sCs8L46F4xZZexYlZxPU
K+LSiJYMtBusDQ9qQP6FhaN3JMCPX6nqKci2idec8IXQCCizyKUCOi8PaHmFFygk6EnDHiFKJbzQ
mgdq0P33827ShVfFn95kuAt8qWEiDl7xwAAzdZBswgAWa6qM1SDTxFNMvStEw4uJLjmfmkNLzC8+
qZI/rR0a2eomAbHnHRc0ehlQD6It0X+GEKGMlQox5KNna/iE5J4Bge24blW4JteSUM0ozFoJFa7F
eIeXoNhoNzF4431Fw6j/XdWtlnVNuAQZEXfXfj9aHBvQjYf4Crtb7NBylotjnLUzUPfD6/XFK6Vk
NDMZObMT24J6WFKq4pXkax7Q1FrWDXVsARC1MiuEkdCXTrnduYTAYYYDvjCsObEIqUtJy8b49xu/
QjQsqredSJpcCMjMb7zKfTxHh10+IVEsb6ocwB12bqmNDQjo23ctRTfb6zQLZGdVaLS3xk/jAMKS
AFPZUH8WiqSYb03Df+kL6vwdmwAIHucH6HJZ+hwqXANHUW06Okq/IWHfg5NPNDiRt2ZhN344MF0m
CrGVP9B3+FFtncGxiKPXt6cUFdBsSmyjCsQxMFhBSSGWeEZKmQBHYyZb9Kbbsh4/SumF6jas2fDG
diaer3FD94JrbIIxe9YNsIaeLVtDkGZvOoQKtD+c+Bj4yGZ40g+Qz3kP5YUrqPtdHrnLRLQa1mHB
6s9/xHCQPE5sAYvcdMzCfLUXP/wy/UFYNoeEo7kIXpodz+p7ZgLkxrm6V7jXqzF6lACAt/pHY6XD
u47HueR+3xve1MqK/MImMBoFV+u7tBwyinOaU8p4nYkGcFEe9u5CAF/U0/mbUCVqM9iE7Crdsg5W
KAsfH1J5EbuDLw+pbpbu7hryJSLQk9sJAXHQRMkW9w6Li3Q4GN2v7KkYiBHMbkaWycZUzAg5dr5p
UmVHcefrVqwWElghU38R6DE0MdG0pcpLQADeWm9eJRaGSGKpN8vBUrO2FRurqCdamwD+Qn+Qxseg
E9L5B8XPtfA9H/xDWLrW2D3zMmsw5ThQ1wCffTSnQwbq0cLuZMb1837fSkM5Rp9iCYC7w5ku9io+
5yG7sfIpAxf5aubQlJeHK8fxVcwIwiKy9/gAwlIOX+x0GPkas7Anj8eAS/VRczHpg302ybOh0IBv
/j7GY7JocrIrurd4GD3YJuwDl0Zuo8Wf+UGuWRvRf3Cf4S6dOGq6r+lw4MGXOmdQvFT6F6cb9EI3
HrRLfomvwlFqKCURziZt5GrEM0h6A8NQZzikeAn0ZBq3S69U6COvzNY2BEyTjYzwvCXWQoGAqqNy
Or+Lwod6jgWYNGAeTM98YuWJQFY7g/MTD3Y2C/rzJ3jNDYKawsdxlNmcrBYC/ielKDYNIdC9K90U
Utw3AvhUmxVjWVWsz8r1HPfYxRVRfvIv2kcHbDbteTH2eTRZzfAiGcFE/J++IXTPGkgQKZGw++zs
CQHHv5mKyzDC8TqYHcuHYYszcA0HIxleJx/Ble3aFcl8YUYEGxUwmFI/kuEsAdUpj5prlD+3fB2y
+Uw/lLtvyvB5bez5Q5FenjFaKgyQVt4Q6AaGjFsbKrofVkGzusloIFFY0FqCzEu83MORxZ9MN0xi
mGFAXEWdxpjNnydbkZoeHzi4ugK8o1DxxrIHOroglemVutjqC92eSAiIPhD85ETQ1jccNa0sa1t5
SzKFKCRtSBNo6YBUezuw1N0SmoWVLsliUU7nHyRMz1JLEYC9+jKXqXvMUj3vmm+Lifd5WbCH/43g
ys3zvgUk7OxmCyZYNp+nIRgd3pRbHhy/1SPb65Pp1YGXoVRya7f5/TqNgVeqEv0VTasG+G16IeHL
SqdYCBJnyIYdvzV4Ttj1espZadL4nScXjitsRewXveagwBUwuntZ6A73tqlNa4D1TEWZAM8dYdYA
+TwiXXoJWrfWBiuiMdvU7A2cFTnZk36TjxbV9PGrHR8WXzf39XFp5esvAdnwvtV7QUGBl7opE8XP
Lqcp0Nlv7K3nkVqkY6xiM28q6ZT3qEONAVIEAORexYETcaQXUSPnNCZhMg89DdEquHxu211WW5pb
Z/wOZU5nT8x6hg/VkAlUreMeZRvFL3AORXUtC1YFpfVsqLDbeKPYT5mrqHOvKHVzS8qXiAXPlFnT
tHXA0kR4W+4ylrloaZVVWGPgqnGMmWaBIJVFR8h/eUYXlgInPMQm1qkNIv4AydKXzJcjqpqJN4sO
TD7zC/b+uJ5xTqW7bU579rNyuorNDGq6obWqb1dc85aDT/xLakrrNdlqCuGJiGYUxbNUJz5T1dHg
GvqSvHXjVBCvW7D1yV14pE2m7FOwt6ibNaxNQ+6/WPufBlIyRGJxm/uqCPIM6TvWKiLdACHmDYKa
UU3j0KFEdNTEmtdGtb9xQ8P4iQaBvGeg/3eiCQF8sD+bZDIBOilVgz01VeuBB3fEemZuKZzOlJX4
wfZukmCB3mvMr/XOgdc8MTXOfTt4RZJIUmP4crRyNRjqAoFJJmF1Zp9VVfzd1ugvdc//qQWr9l+9
RTUd8fntPhSvw239znVvJkcAtdrD6G2SbY29z1KghGGc3ojv9j1yj2b2zTBvCD/dq4Sn2IQxZvcg
BuzKrRLghPlLhHZde1/pAMbvCWyfdWzj3f7fIQECjR7rX1VVKx1d0w02uOp4byw2nf23RvO2SPOs
UNsR9lyDy859N/1fXplh9m6/9VmmTjO8yQjqNDecLuIAOhR8AVa6VlqvupqPsOBTB6IBMazguggE
pIEPXLruItgq91mNqY38biTsS5k/YYjQBQTOIQMcDLE0SFj5L9GbooKHV0fQp/Hjuy//vI9FGZCz
2yjSooUYnO7ALuVYzG1LaxDM/OAsiKlvDWWw9IgMPOM5KUuCiR2xNnPqEqu4JHkCNHsAugsLQ8Be
hf2rW8VmgFY7Qeg4mD+zn2s/v51MFuciviSFLAnEAGzjP5ON7WmlSaq+WrccCvStZ4ZPhcsoeBfd
FvEvIT08sS9llTPg4vDyTWhwm9t2ifFJI/RL9Sik1Pp909c2w2J2A2s2PsGzLjSfvgLIhTNqklot
ID7WeNnXc7eVNJ1wngsCqr+N7LtV0zgbVmk/3PVU66kOU2m5sao3fZ9lMDtRzmN6kybWjncn0TJL
gcIAzXUJWI6rNwyLF7/K8VYWsfddKBHsLi83vYWq3sHz9fXatoqf3wkV30C2JBQEqPXFviwkOZqx
OQMLpcsehP7EVZo3Dd1biVqreQYehBr8Pab1sVdqG4e5Yw96Axl5TIyoG5YOHI/4WqOVjC/EN6VK
3G4yKB7y64YnqMWOhV0felj/s6adDGQv1CCKlI/Y97KoKMSNsYSOPpNihEUSiVXwQyb4Qcu+oDxs
4oe/Sg6fi9phQ4K0cI2+0F0tlbeSrrRdJmiyCYpY9zNaSLiKyqkGKFJieiPykgP4knPar018tWwE
zWlRN6cZ/yKHdEU7TTyP4FMywhR+SbunoKylurKrw0I0l2AyYwWHRDtZqgaLiRGe4UqWBJcsoW5U
hazE37as9HOe9u1nTvayYqVZHinOy30CTUdx+sdVztTMRFbUh+Qs4xezMu3USa8vGHGEyG4qNmB6
D45WrU4bgTofQayKAsLEOKLkRo4klWz3rq0gaFGNKxzdkoSHgaLIjOvd2FEgH3eU7o/wP3KRyOTH
0DKiV0v6UNPg2Odq5msCIORluyfllRVpyRijbk0/+wA7MShmOY+7Be4+KvMY+kCwS4qDd0COhRbl
i/cTPCQTQeXvZBCfSF6Qi9jsWmXYrXq7ADfy230THbetpOeRWooMNK97Tz373TUK/8keQHMVC0hK
EyUOMLH6bJ4UklSoVn0x0+0ncpOjLKCt4aoOyGV+spVBVRKfpSrTzGN1GQBhQ9xCLsOMorREnHrB
P/18mwWpLkCQdRrPizQinCFYYHfkzcnDY5uSTke1MPJK5R40DRe+g3vjcsncgC6a/49ERu0v1HCe
2paPU2tU2qhtYH8v9KXypWusT/ZNmQOkab6q3cwUvIJNySQy/QtAaIk+/VvHJLUPsZcRh6WiFRd9
x6L874E4/ZMgl1bl6kc4aoTeMSYYZlzC8Cia4GwRqI91dz3S/8npGWO+DekQYFdeoD7fY3ThKKdp
MNhVtiOxK2KOY1ZWDbTuUZkSyqMxb+AEUGG201q7YFRT6jN0i5AcvqRE+Hl1G4x/nnjja2JeZRro
qiRdqZK2AEM0zhwWt+EiG+s87vZVfmwWbx+n5+Os0NjiqBCF3WKfPfzMIE2xu65KbY2ZrRr41rcy
ucMBNVW7GmQtVv/DUGfkIeiKCcwqHxd8uBmPDExjY5kR7y9ds+JfOdXDEx9apXi9UzzZWwqn1t0b
eKZIRVHJA50K9MNz8PxRE479PcsZpMkT/2AVyynJSYyslsndGDCuvCkIMj45+oyMn179I7aoFTeW
+Wsp/bi6tYGqb5lSzKlPP4paEj5g3Jh+72h43qJK+S8Q1Ki5Ebqrx0SYN/jry8ll5tDJLk5AKcB5
s6cJrZ40QEnBGGs0SrZg/L+BYxJEK8Ol6d4FDP9zf9/P9fas8goZK0p/gudoJ/j26/68zGhFJJy2
UuD5gP3BIdyW9KH7GngYx3BOpf2IDq8C19FV5MLlsZ+GJc1EkbkmorMCuidkqKZAaTB175v8AK3t
Xrftpyl/ATRJE7PiwMD3Ub8PbWOE0wNjGPYse/7Y0e3cs6eag3BRmGtKf9WTllzfC6w9nZ2W1o35
KYoLnyn9Zs+myPfaqBaW1qfhJeNRqfF6idoqh+eUTxgwrpXJYMG2VGZRBLaGAZwruNIZ66RNUzkm
18R444RAbZx2YchsEyCU+YLvaSHA6C2glEsZ3jUITBJ/sxHOKZua7OqdjMfXZCCqrZPXPNV3Lraz
ne2EjtFG6q+lgAhdkNdZAqEPvxHiKuOyoHYHvN0XCl4t/ZmsY2jxm8OLFqBzTZdqv3l1Dj9Mos/J
5tWzQTvHi01vwDwGlOIt21wOcNOFS+RfGUj/kcipk7aXjOkFrxzplENVPpOQCToTwIUNM7jiW8RO
0SJMJDOXZ4ZHZGrcTxGWX9OE5554ImRK59EReXh9ZajlbcQOoXp+ET1lp2Jp2Hmw6tq/wlzx1ETN
Eso/GqNWtYsWiaLi/r807y2voMEJn2PyU1wRwzLPENcTLadYEOlGn7ImHeKDpLCM0VltMrELWjcr
2Zquu5PHifD8zyA0VUV8+WBIzNUno0qwpmXsu0YuBgnoEW3eQ0k2m6xyA3TUeIyf5rRM8icIiQYE
sQ+UYP+PzL1XG9xUASHOMYFAwzks22ApQ1xpXyKUii3EECefMosrLSLhb97urtPlx2dFcRrzOmp+
H1+te3WW3sOgSwSo4Mcy9PBrIFSzHmdSOJPBY4JYQyJYMhKQdRIN7sWocR5ukMWC+IWtDZQCcP79
jBS2yoaAl25JViPizpGe1ittxCS70lRTXApss44hEL0XXvTHNF/uKTZwa1ec1mbwG6d+B9BALQEz
qZeIPv4QHuhZIMyDNrOoZwXp8pQiOQqDfbL8gowQayf9nKfKyrxgg6P3LAYZx8ALz5t4LNWJ9lIx
NWyYzFSM2JXaS6qJaCgJif1b1WpFCKYeLS1+t5TPrM4Yqkw+cFeYcbEaqlPpgMidLhVMna659+3F
D7AYtDszpxYv1LAZtxLqkt2VpA7ysIKBkhbDJ650+lsMYV2YSnuNV/gEwcAV8XyG0SBUmCBJuEXt
wioACy/nS+9pB+8JpsuUrUmzOLwtV1W0mZHYZWyUGbADemNAQvl7dg3KD7o8hicGrsPEsrvKwQn7
Lz39U/CAqY2aGXmHnNuoRusY2bkgFVF0hDfydd0YEAdkcphaqVoWl4LtyGVmJQo3hzwGG3qV8maW
7/5VIb3rh5nYMd1FBtVRhZT3B+jk8yP/IoIM21K0FwkOCOZWoNrGBljIyo92CV0C8kwkXaRnY6wS
LFsIsiT7Yau2EMxKw/0Cd3xdVNeTWiOb0g3+fBsDU6N/gBadnoz1/NptA3KF3KuWjojby6FJ3MdQ
R8c8nDWxcTIOLvqX3TS8Su0Kr1EcSUQqKY8Cyig4QuXbv4kMa74diFAaSCY+AwBvsR1jY8AutTDX
x2mdd4wvA5lbrL1gOToKReV2Y9DTs9JETCoyLVw3jtRot/zGGKAeUhzDlbfz0KxAx8UxPO7uQqQr
yxIYdg+8gUUJuZEybBQujAJh5OsY8+AzNmFPzOWuIPViXqnwdrBEcgTUHN8IcruajWbAvmfJ3FRv
QQIft9Ltborfzy7ntMJX2odO6rmSoccuYcgeUqFBCmkDI2Sy3zW/hSTw/K7GCPwMGweREA//WmDP
pGMtyS9MmVKqLy/ThznMGiXLyqQ1fN2w/XHOz/ZkDkC1cniImmTeYezevEcVSPKrZ0l8WJ383hiN
ciBHX0L8dU4P5nKrvVkXGKMBnCz7f0O2efdRo3Lei3E2hfLL1dDeDdKDCD3chsKwUwF8HQsElrPj
wXndrSUGPryJRZslGj89wNpkOQXMiOYoRMhnhZw9CBWVcAWQy1bURMJKtRITrVufHb0piH6FH+3I
mz43N/UT7WO9rRD5RSfnCmGZRFo4JCjwnrmZgh+WawwlUPolcb9NQNPVIfrR1eNlA1CHyADu7cYN
Riyta9ArD/WQDCY95iUcCSBtsHSbreNjKtY8890QoGdzTetmEfKfPFfDWDugXwWYfQW3DUwxVQpY
ZnBDQLY3yEtmdd1Tcm0qp1Lu3MAl+jcUFEJnpEQwqch3jElFilHEzyG7oR5HPeAq4f1Jg6TXxQbi
bZ1PGqrSDDLPTNF312r9PBjfBbQvaNeJKoghO3FbBxrSVPCW9//kzqY2po9ekAlcvBQ6LLKxta2q
s8qhjyQwpWYRa/hEPsiX18mCwBfxS3W2E8T0cadf72w1Uh04LABlPgHQENfEewpdH7mQHeiHFIIT
h5v9vbprG+kSrdeJae1z/XegTwtJBj87L9fOrAP7KP3urJU7nwc17CuZcXCfkg/NiFe4XC/sBLbm
y70ZxRPXP4BZju0nNKzf6aGTwYcy9R6D+yJTlew/eqClDWdZi//ZC5WOy7BqJZ5xjU4TsA4+FnS+
p2/Ew8KuyQtpZ0TsfbywshfU1nsgPN34YlPTAeTlOQLa6WYDff+zZE0yf5I3yWkWb7v3iUMDKeec
7ByBmL1u+YGXmDCbxo2vNIR+P5N7FqKEkpOj0BA0QQswG7tfXs1ozAmVjxUAAmDTicZAAa5HyWR/
QvXEecOa8A5adwMqSpN4Lwob8ZC+C0v8+CGHsrcCdB3vFmPlgO/Bqk1jOCqPwJct701rOLxvEMvX
3DlA0r0Uc6uUn8ghYHBUYysoM9VFsqSQOugkp/tdnjD71i2dW0yVwfG/BiLhst/59oNWNhxL+eD8
PaYJb5YJxFVlaNSd++70iQfW0TbJfrwGjOT01Ut19ODdcNBiNyKIbJ+ZzAC8WEX6Hk7qSH/hQdof
2w4OvBPULM2TU9z1fsE6tddPz2XA5gZz76K9OvQ1+dxihlTczoDOm79rLQhkFAAcz4hxWnPeDvXD
MAPxZoAc2fIvLZQEK7XKJzL/x53wTBqvTnsnDd0wT46U1BnB2ABUaCEa5oJmQM7Rxekkc6YjZ4mP
h3N/hM3uQKVu5C5qsE9Mepu8OQ/nb7cm3zpkFZuQ9bLps6wm1r5YahLUDhT6OukYTXYuU040h83m
R3EPTLXIcFRKdHwt/OB9ahLph7Tv/9XQO+sjyOpqP9Bqu07637nMmtARppxhxyYmbvO6OhZl7RA1
fKq81vwn+HkGHbN14vTDXWf3Os/dCbLlasUsz18+mSR/Vqc8I0jh1BDmDKSLCNNIup+EC/aODLvn
IDGmhu2xcgjrewpTwIHBJQKX4fFLSmw/zZUu5u5pPw6EgX35PXQX/3FiMxLnwdmjO4YjJAlPxzAq
qNAhWV2Ryza4OLit2FP/sEzpjo8r3ujL8r7+s9zLNiVfvHy6X0yNH/3XdbJ5fEhjH8gmtdHrLuzC
kqDfzBId+tl7JrjEXacE5Z9etF+5X+YvreHMvG9++fLwmn3UNwQIiw0brlOMz9l9Rq55VwUJz6wH
mBnWqYOk4FMySWdUWVPPqOloUY0JVpsbxaYHdo14uf04+2xH0Jincuajug/w6+rx4bpnrBlKcCDY
fMPhgfxKyrbVh3EecrXA3sYbfOB5YwcowQLZ4SoKZbtGA0UDdqq9kERJCacdxYyfFKAoE8HimRpb
/UTqJjnack62wnCh+chBZavvllmTngrhug3YwU6vb6BgZ6H/WB5irwpfsEjDPFnTVhqn0xoMoa+p
Qwt8RUq1jfnaW7wnlTwR+Kp44ilWFV48T/OGM8OawTL1cwQCxhMak4LESpCCq6QktaYLDpHWl7ns
SjtGfuEtw4hz3OSK2VNxjqWjAwLG5N0diKdQ2VecH+d8p23RVG0JfC3LynfuTwvJ95yMFJ2jzeMB
Hy8Z+vDPjWLrbRDnW1GDWp15byv3X+CPspWDn4xd3F3bCiVVPX6ASD3NqRGtUkr6zYI9ioBvWgEr
j+szoOKYPLYFe8TTqpLsUgMw1DCEhSuVjRN1OptbTpWn3UXIaSix8zOoGGYbZV7NcXIoZTD/ZgQP
8EegH+VEeyZRNcQVVeA7V8NgDdCgAMYhJdwl+O6opCAXLHeucToua8/E/F6DSmB0bi07/sIurhaC
VDJ+A6pUc8UnWLyz35ruGaMtrNVYssNUqDLdQZzp4feTAtzwKV3UF+1SRLP5bNItBZrTMoilbWO0
4ahlF08jXHBlO70tSmojDJVre/ZefPXXfm+RnpR1xodUoMLqAkt5Coq176SLsXuNlFD4FhktF3zd
Sw3f+A6YNe5CAMZXZnJDvXdojI/jgRhB72/DovBRbRrGh8JyCfk46+x6vlBp/BDafisnl6PUPCxY
Dr5XxP+AjgbA65Az3zRTKYnVjRJiAMkWdUzBXR2fsiBudGn5MciXssoyQP7wiskX317deLdAI0uL
QKj/rmqcku7F0lD26oC9W22ac4EsIHwWYSYFYj/LcujGhjJM+M1YHI6uVClJC/rNBgrMTC0UH5FI
LaxOXUqWOxCXTDeLwt5mu9J+7vEvs/uuvdhjIOr5Wk29xvKLBahQXmONZO8xm9N1se2aYy9xkKrg
SS+/SBQnFOtlIbBz1ryh/Q+lAP/oJSdDYAazOzMYfgqIssrwjI4k0hdki6z3GJUqrZAQfZmUKbG8
A5BdGRzeBcudkFrY0xOcA7qAEYX+rh8VQDBgE4vb4aB8HKDAww5zxAeAuVd3/mArxVbba5skqQiG
+N/GdV1S98PpFvEARzoiWCv6oPHwIHTkrbwLz97PDWTRzSyhsOTmXSvaWuZNRQJQnKgQRHO39nWW
wIOr7MfTYnDigXB5fvvdC1/zG5Wj1nPzeEJEu0Y4NkVGR/XTFhSgziqI6BGitCv6CruYl2jqX97/
9XGZjb8RBh3L3xVgdypB3t6iVXYKqJ2Al0yXEelt2O7gI9iK1W0iOaDYDjxXIjH4WQLRZHhS4IHZ
c3PG9tC2p0berfgdXmJjgeDTv7dbdCtZThVh9tUfxJXuIhi0hoibVUenaIHVnLbrmR4uyo/yAf5x
VfUhoMo6//wjACjvci48udXjEvMEG3Sl44CTHBquQa5H//NbkSvI+2lGmAtiJSYrD2sYaKeUarDB
q1CbiT+60hV+BHnq16oFqpcklRgFwPvIQe/rZssS0QjW6JVuhJIOqD9vPe1O8CujK7RsdQwWGfX2
+YZRh2+b4SZ7BzlDLOTB9XKAFiYVbB12chGUiFLRiPEXyJ1I1epmxOniivnoXq6tDX6OZvnEtCpD
SmaH8zScKg0MycfivqyErjB3gSFeU19vRO02gwmdOSr1ODUBivfieg9YMzQxMxNFiLuqbKIU4169
9VlmAVcHhafY29m9A8MxdpRodWiTbB3580Xi21pmnB23JeZcuX5b1E2+yZmzTTpMwuhnAIA0/raF
fo3In4kOssHpt79zycxjT5VA/ftJWk5nT/ZWPt9l+jz6I0lmTuua8jRo6S8ktSTOfIu/P9SrGjKx
f9N6NshTxh1dy1fZOfpoPOOI6AjC8pZ1QcROlUJ2sBtVamUJjCYljblQI1Xmz83+0Be8e+1Vqkvq
2EVvRHJmNIOHx7OlRZNP9QRt4ekpn8c5l5Ud3EungGPxpNqWGBVfaZg6BDmxKmBE2Qe7uk8DGjVa
cyFAmDciSFrgwhLykvg1kwBpPLBGzvvulRTtg6482W4b0V9JBKoUiymq5bSrSDYHqdhOFpXEil9G
7k/vsyhQWAR2sBd7oRtMthWQ21xXhJOuVUl82muLIJ4ncLPB4z4fx1aU4R4Wi0UVcczh433JXpTM
Ka3upeBEIWOd6EHgr5dN7wJVFbyX6o4fRw44ncmz+6En6/gt3aqLNb/yuxbhh8opil1XomnO17pf
igXlCy9/+dH9pjvGCZJ7adMjNqXyfZ/wjtFmT7YC4j1Z0aYSUO5ZGwdBGKT8OjjieeFl5usLwYJx
Lbdkmb1U9OFPFCP25kY0XMlF5whK3SyH83eZxsS1d67O+AxkHkwyT7g9deSC9M8a6SVS4+xWsdU+
5zqvop8ei2+fFaiMxL7KsJHbrCE2tl1jlwTMAMMokfW208zT8SBnYWVhz8J4/3y8HgV+8c+kS33H
qs/Y0Oas5qoVNYrAJH3DLmUhBLZdOQHjLPnVghagPRoUGgUUw/3I/ALPu+kcnxDfPV3JW6PCSx6g
lxUd8i1/B9A4+gJGjIwEPURR878VeuEtN0+VrpPQl7a8dfvrLQwE+90YDvURHaoZGvyjBH62LXY4
HVd0wFrYe63ITapHDtbC8bIJEpHQbLX/JNkQOLS3YjBOU1nb0IduNt1I3ZLnqnkVaZ7G6LGICn6K
bvUOmpI5Kh4WKplFkVcRA4g2X0dQynzcAq/B0KRXbyrjlBhl1TSs5WAHI+CIebGMXIo2Qwd/nXap
1Y+q74RzAuWOje9h1Yp7mIbJYsa30vIWvXtlTdWSnPvCv+/vTed+moXuzTLbA3kqqjXBvPchX9Nn
oiEVA/GCMG7gczhpLF1smRWjTG8LXPeutbOfdGe78sGWusir+156e/2MnKtsCIokDOhDAzEXHH3K
T8lHDPgV/TZzAMsnKe0HYTwKbl9mTutMFX30Glx0I67R8ySj/WeifZnPra0tEWe/4Q/WOPsQOt01
M0x5hha8fso+lYtVeD7PG0NqWm3pyVF+qoJ1JEuW7s1ryzNHaTNuB5QjhU2drDaU9+nS/1QZlb94
9oVSsPgQywrfa5QxOJ6XYqWQrg4GMTa7vqCh2aftTv5irWa7BQJDTw3BMKzqVNtZuyP7hRLXXhej
4MM48HDo893obVIpKpPEAaVsRNKJOAhM8kPfUQp5XJpNxYbfn0AchojJrhLIbaVoP3/dC3BTICaf
rkTRHjNjWAKJ0TjTIG//TEWajL8tgDPCA/CW17yvQJGhWifsC4I+KAOYbqafmplDrRwCHpyQ7bcn
+hadaBoczp6mB9hIycSvYN/oBuDQTeuh/1WVNypIMeV0Cvlb39aqcjtx+5/3+yGd0JFZn0bWJC7B
aXo3S7j7acnSAhpPxGoJi7Y4SN+I/FVbFLnMvJSlXfW8tnBOjdOlYn37zdQUkGjrMk89zPz9KuXG
VIrPd2vNjFdJkskGYknq267jFoOeoU1xdA8BAxL6AiNVIrLrRFEe0Wg7WqSXrR3SldxBuY/l61BS
HM9HJ6v40J9ACzdE14RKblQeew4GTl6d+80lT+SbV3SfEGmDHsbE/Gwk9CKXVoXuXHxW8XAzJxwT
M0HX4FsRqLQPVAjqBzXOagCv/pbAuBUWI7qzTzZzFv7kEDdUASsHj84jo/nYLW/j3eCrRPm1Dz3T
h2ivRPDXd1fZOlnwMz/IGv1Ib9t6sU4yDk3IOko+2oczMSVEpk80daFPlOkWKGZOr/iABa4lZQpQ
psWSBboVsCYFS9D/huHRnEeIil3etpPbSlhp+mDQ0op2DiCqr1uQzWWvd5t2JsVv5yjUJeN+MuD5
6f6JKU6rqJ8tNk6LY5Yamly2oowwosiu0nwd/V24znKSEcZeoIm72xisXsR5BtwgsC4fqKwml+A6
LCD5ZFusNYCasOoQHWDAO6tVOAVpe7hz5AIC0Y6Z2uM4tTG+tD4Gm8aiELgD88/L/iNMZrIUgdHh
xmWJD7MgTb99WTeQhN5CjSLYBYA88uc7iSzrE+kJ86lJon/XVjDHWVTIp3T+CQcY+OYfNOiQ6S9i
DmxsdgGYxA2DckkhDBFyL6MNAv5RuR7DcW1SXlJ3Plb+Fnr71L0uWaQdpAcGaHm/KGVL16pidXBF
Fg5vgaOmXzhsRN+xJUqqdP0D4zQHbraFaW/gMMrvvdVCo8zgJIlgs7sAwwSg4itsjwuI1PQcbayn
QWDBFseATAbYPCHBHUVm2ILD6WhSfyn7zT8N/zkDtz9Cm6L6C5CsIz88q9erWQz1/IYvuieQGOkt
ScqjdHnsJ55ELf+FmVfM1YyjFDa0xUUWDihK/8uILQuDtC0lLUqTCIVyGBeFbOV0y10gU25/ZXpZ
5/bLER0HjAerb84pOqQItq0P3jfzqt9thpnsz6EKsx9GCBMOOIqZZvgfzEsLwzRo3gJ6HuxXAu6R
r2ItUlo+fjmUSh9Dla8bSsGK9RuU3AQW7OUeeJoBYgs5lCtdSolgtvROCMRZ3XkhWQBbZBSLdEI1
QoGa4MxiZbmBK5r6JraT0PKjjkMmkxoGnV1ibO2ki3sN9BSUZByjbimevmsk+MIsLiFjm0TNolui
EuVoAqQRc40AZ7MivNGP3VRtseUkfvhJt9CZ59dx0HVb0ooneYm2/GlZxcgkN1Cd3cuESiq0AUP4
NuJKWrEjIZop08fj/Wulea/NDTjXBSd6PihVrHj37cQPrrLinm8wnQLmTw2/+cS6p6Ymv6Izs3ls
/NW60TblEHj2q6+cCmQDWlXqfEQW/viwdXPAeOHnWBlRdf7Hz/cs1t+1zcj33TnIaGrtLplOfD7T
bPfp8gAoYvMGJ5u4iw5mR7RxfSXp8QRPfRv+Xen0ot+d99HR4vJF4V5cHoCEVIsKjasNIhTwxm7q
ap1YixsBpBVWWZ55ur3WNfnQv2QhVuaukdidlXydx3JgzJrq0fB4+hnedA81Z8B9z3fr+HM/8gyw
IHzFmBAAOor7NvOcWLmS8/wfJrZJA8y0rD4PDmJyn1SU5/QyB9yPOuAQAmpVElHSjakbnh1stl9/
j8TkbyBoFSARg88bckDfLA/MNs46WOdM4cEQ3+Uyg0nKbvxsECokrj+HXfs4K79dTIuBC7KO+QN+
RBTCm1ZERr5ePyhbFQw5MDyp7z+22CmSKrDDa1ROsXGkF3asXcSjUVkK70BOid7Vu71+fyv487W8
KXeZnQSooYKdBEJTtUtJktNK43dctb4KQpepkIKlR4dsa/LbTwmCBpFDYEqvXBxcxX/AklEK7ngO
MfNjUdXufOMrWw6wfFPHhcMQ1PVgW6GPk28v94THff1GW7GvjTM5UqoSk1wBRB4IFMKuyCMnicvT
tsh+Vg+qrLk7eOet2aFEO2ZOFHQRjgdrVgAQZIbMSTRD8EG1Fwa+T7upoFz3G/bZJS9/7YaFALGB
tVC9ysY+6dv/9MuXkbZe+qwDiUjFBK4kkfhvBqnEtgzzcznZCCVvtQ/OwNstv2hktPW8FM9m6fxA
HGb8M1fP3js5pFS5YZno3G5pASNrsdStitTQ0eW/jdJiNRvtQzF27Rml9Ar35WOUXkbdLpYgG8yf
YOgCwgg8vTAJJRERX32yCFWPvQy8FmhFSJGxPAlmlhhWGM5545JcMdxlzHN3oP17ujeBzrBJeLxT
OBSAmNheN9Wwez5VMKHMQW9FtSg5W8fj+LayFjP7Cenr0p6RmOFb13oaq1ShHck+Fa+/m3dMP9l+
IZkdI3D/uHV70I2Lb//bTrpNr5PtPCoQY9QBgW+JlAdoD6H1hmUezLsBL/Cj52rV7PUiYR52x7PM
hzQSlxFTuenmhc+WsSj4NNH/VHOQx17Ehe3f6jYhW2wtKcC1wbxZnv1suDYaGsEJgk3+8XJLYJm4
UpBPxiDQNuyv7ldZALTnJoVtqAR4r3u6gHrdKKNsXeheIaJwHtWtZyBWZtkQKBTXwvdekxmQfcKJ
78bSQgseJMcyBU5sA4UXrd1G3u/heDSTap5GO3JyELqq+5r/cGC4kEsHJSMOs0YynV3nttfxWXSF
Pjg5fv1DAvQWLg/uMR7iXOM8Ms2lAZSbBkAlMUzceMUbbzxHoU0tFkDEEFxOZQdIEfLTU5TrnTei
1mZTMYEanqvt/pk3JDgqvE4+jm87R9hZN3lwRK5RJ++5zUfakYYcRkno/qT33+FjPthQk5kDSd/y
vb4yNjTxSBj+zGXMhCzGvBOTtddGDpyzdfH19Plz4ZFDdqzCtsVCTwUSVScQE4oWg1MYHcNiK2nJ
zbUJqHjkJ43FdGMsP5pKHqNbag+7JN8v4o/unFtb2w/ZX/SkbH1Wrlp1aGnaPjhCb/8kdoJIyDlz
w/CIRAfGHEJg/9RUzP2iaDZwgHWh5hDUkiK/SYGqikjSSk2+rDA9hMH3W1oEuopxnRAkJE+hQz2t
6zzIR93aJoG60XfmeFg99XfFL5J+0jl4DxhbQw4f4HOsK3RvVzr5B3IGNaj+rgLzDAiP39uYFfLv
pIgDWGP1RyN4j8iEZi7WZAmkhhvyA88kNzNeebaCxC8RrQV8EiZXT7HiXktNLxJLG2JlL4iNryXl
PnLmcNhIsuuCv4lAd44Q2/r7ADNOexsBoPMdR4C9OHiM4riKPpkH8oeKErn0fPwSZNuZyh8wB/kF
7YclrnqSU7I28bw/cqVqG0gCK4GI9J1ahzv7P5fxjaEptBirwBvVpGmX3KhcI/TBT8NOv61jdvQP
VG5Foe/ZvtMeVRpf5c5NBdUv/9zBNLnp8jcoFw2cdL23KEVCFqYkB1qkSuIN+2pST4QJExlrgCSP
s6FXNVmbeEXlFLIgEgz1cK+N1JFlrm96J5+3jIhkgh0ZjZPKrzhPuBGMwtK9z+3rxkfgtmyYVXw+
fIk++nfCv7X3hUOBsWrzQrN5Z3Q+LszTVnoTTemeYnzx83Sey3eZODAIICJpGzABqvek+2TXDS54
EMarbxHAF+c+HW81EMIlR13KRztbrw4wLECpls6+iU6b0AqrWHPWCfu8A1pWcw0UnbXBAILR6FRa
JIilpq/DAEAt3AA4+VVFZHifaNfB/Z7nBWUENvQfSso4djSRlpfZE6cDpqmCXm/il9O6rGghsFdR
gyqgOHuXAtfyxWxUCXu5svyzJxjntaNcyi6ktOAcIyQVEl4EwTcgA/WPTT6PZ7VG3V/yBF/Br1dJ
xwGRRaKHYNFfyl/KeStypE350SXyh0Ic+EZlP/hLTxUtnEThewjk08jTXU2nqe9H5dR71YcqfRCS
zrHNqHE9vO++2dpr7g7+a80+CY4R110/QOwX0RiA3Xy7KJYC12zowhxyVQYbcrScY7O3NEVhUTSP
TaAdR5/TWJrhXMt+88YtvpgblnpgQo0TXcLgzc9t5YjupbtXPGHp2h85rnnRCOzBXa2mx5h8HfmB
KIpcZ2cZo7jYQn+pyjwSBH1z4qSocUoEDwZDWD8yvhpfZmsSvIAy8YEHmJnFtBK1BMST9QwlRxmD
xZgio3UJoEpKmmmC4L+jPtpi9DICK4B0uhQBTggxUk47So8nYZnQW6NTr3tcP6w600ZkiyMg3E6O
MHp1JqKeweNLAfU7u+ET1wDthsIKupAoLFevnou5GJImPumJdo8poIvxGNN+PTgHKIy5SpgeVt3Y
qHNJfzW8K4HvEavKOF46WIJQuFrN1Zox+Cw5Nw9bsw1MxnXdq65yXiMef5t13+jGNR/dch7XSbiq
z7xX2+2LJcmTXBGRGMn7mHtkGaiewvnZAnQ05YqEjdoXCkmEdQsEuuj78t5k+D5yG3dkDLzoGKbL
a0ufy5Tsd/6+LmG2RFKs2carCLQi/0JtrqXLyCjP+8voq09Hvo5Jz4Kx7C7Bvbz1z3hp1x0KvAyn
881VjoSjRhWrM0fTFVGoDPsBxKas8OTBu4QbF0HAUEImzWgIIik1ms4UZmk/LdoJspN/hdn0kpBn
RNdDhjQSDuahXOs4s+qrJEembyAXtZOtbbVnkG4v+vdE8GdOd2Hb7DfRlJXGqmdLQCsJbGvsbGlq
nQkw0YRhXgS/INs19bQ/D8l40KTYf6xo6QtjfDzrkfQkXqdwvSHdxANQdD+L3Ze7DZFH98Plmxf8
nzy/Sz81BVlgNT5s3lVaarkJtFy2n6jHWEnxluYMlA9Spo9ildQ/2tdzZt/kUn1wtd6gyuoMiTJn
XlMx7jvUFZFOSVQUrwoqnJagnpg9bZIoajD101ryrXFRnwWG5n56HA9k2n2EWW3cblZghbj+OQ3h
9Kf0J+5hkGlksgMFeSGVkP1Oz2K1x3yvaoWemjmSZxRgmr2bbUv4vp265BnJEggj95I2jFpq6jud
IncQNhDjEpo+DvR8uHupdM3og5mvrEE1m+DtEueGRpvZj4a9L9BPfLgPsAcCJcCyxKpfo0b7rO52
BiySvnnbVP9QY/liIqu0KZ5tIhdxgodlJXkHR0xNjU1UEP7DfVEHFvv8WP2dIo6IvYY+j61//pxP
VPzZjMfhvtqEPxTHvZrGBgfHliKFOUGbQfBZjrOpAPkkczyno8xHryUz50USHGG06yDnJzi2uYbo
+q1nlKgV8xMm+oZcKd1remWyZ9KcBx0nBjLs5cNXAwvVHnfTqxqoZKXib2n1jDs8GTogFypg2iuv
kDmA+76hmR5pz1n423lQk0YTt4sn/IfW9oT1GFmJTmFpVypNj4t+SUI7wtrvcTz2j8UZFW2xSF0l
k3ztPSjNsfcF6JoS0YvBvbhgPM34xvM28uckaHhEkqf5T8sfsSmYYd5lcZ712lROst8F4IWgRB3e
cOEEo9QAakEbGBWc2yQEfnHf7ihJ2Oybx51BZAnuo3g9E9XOE1XUZN3hvuuvYU8PpXMA0LNW5GXX
DNSAY2gnJUBc8x9QEMvXkdcSI+l5nxGlMntOcc6RvkAwUX7kTuT3Yvi7KPrCAUaEuAucy1A1FmeM
pULxuVsxZUoM9O7IWIjp6/jG0hdFrLaGBqDmJyVcwnWc7IUdxlaQwiCv7SrtRoqloKVlgfFcnSNA
Esnav7xqKfuIJZYws7FLcTjZ6Hk7bhBO1ulVoFEokcUd2AqGnsnq+31HYKRf5j3mWfNVFM3J6EdJ
tHlS54jkvUQQInx80/7PwpWVV8u2dY0VvjDfcX8JmWYpbczujMGLmjaIhjxF0CzLTOmDGTK4UHdn
wkn1mXD2U9Gd2LhdmfrZMUwRRWuiDlfdzwy9IvkqJ7LPskiB15LymN89gCl65PS20lGvFY4QzGUf
uCkDtbT5OxBeCXCWvyb6UfgQBGnaOqOxUZ+FhBjBi4n8i8JnuwMRK5dj2C1+LvsgX5gtSJtml0uy
17I/akXMJjYgyFZOlvWg59L/RmlJkQ13tChfvN+flDUFDqEHb+QVidcs012Swu4XGr4fOwMH8gIg
yIHfx5SNYMfXi3iULV/dTFHdYAl8TUy0Htiba4cs/UDF6UhqbEhj9g2ZGAzA+qVvZc+k5Yx64Ahf
gqkAG60i4jXBqyWP2rHJZFU/9DTTZ5R2KiESbchFst73MixX3jGcWu1MIAtUG7GKJm/9mBrmuBUg
pxy6GM130IZi9G8sAhOHNgpkALzOdvIshx703kKcThZCn1wFy4GcwxCsgj6lrPSaiMHf/cNJDKsW
58gTxsAVjnW0bF3rjPaVshCvqxOwgxzNRQpVvUuavZibFqSYrFkO1WskXb05K2zSzqIGYPoREn8o
y50h7+jBX9b2yFXiOAYRc/r1V8p90Jp9Bi+eDgfuaWNMGCZwgL7dYlY8BKG9uoRWO8tzC4pvsOur
Mpyz1jFq6GjC1o66RueJSz8ak6yv+ZHBDvklR1XwGswkn5HAefFfVTeUK5TOclnHnhrhZJYkbrDX
IlRtwpghmc6psxFU24A0DluZ39LPvbqWz+bim4SKbZUVfUGKU3M2oDEmqilMopnitq7LCyZxoGBZ
w/m/FKlBZMQz0zSrMc+8trch7NaU3Eg8Jc4rPVC5Nf9b1xBQ0AaDeg8Hveh1OhEk9w1UzoR5uqfy
H+KnO5fA/giU9/KRuimcZb6AIoTBgBSutcjwmd6RuaKe2Yja5jzM/W5wrjQNCL0OuI+Y2HJ/rbGr
8BOP32K/refqhFAYr1qYaqxrrptdSOwqBWrQ5K6gTZmPIE2bR3hzhfb49C0mPABb0FSOOKKnTgby
fp8AzWFbd5J8A6kGlbNgsSLYxwzP5EqozZ6OejQaCijMAb/fN/k0ogqrljoR7lC7BTMv2dGafWi7
sDSk1V4YqdiQXRDUyhePXxJJL/Jyuz64B7x1fZ+3vGwkcvmn2o7oXqmrm6Pf2ZLIwLKdS8RHc5WK
MPAtoo2sPONyTsgl86yq+8AXOCju9JbkJf1Y3fT+ZzHUvEIGNBkOG7amvGt1kqEz+4gxkP6Nehv/
1ieyVP5CfBllexwCBXWnWNooebpbwxEk4Xt1HLTx3rSG4GAf98QcprEUJVQ1tt58HAgzlp7E8prn
lUswKbx09OBTqDyIuuMChAaqQcdNnmwUpG9znsB9+mkmouFZY/l96dcl4L6+pzZTq5UZI4yKtgUY
Cj8K1xYAG3qbWyUMMgUr+fJdO9+J9sJHAaJvC/yXRlz/04NIm1i7nUdeYEmd7Hh6Jz8x8cpDRa3E
8RXSCl8vfy9N9KlUYfb8JSMBDnPIYBbpHUItNJ9oK9HkTsRKnmffGjFNj187UfaAnX1WFtUhtXTJ
Uq/lQ6nctbMaeQbFs32jkDd8DSjkunI28fhzB68Qvy1VfrFKep1mBioucb1pbd7Gt/0pOdcJyY1U
EMfc9L5g6I7MrMe32x8AESFXvJieTVr7lk7Ljr/JOjeCEZpyxYHFfPxQ1AcDVP/ZRY9qcjg4PRJy
81uo43GYcKZjBvKpW6YiR7IIQcSY8QXQq+ZUy4oAu0AN6vmV0Cc7wcoFiZ/J3Ci42tzjziw96qiC
qhyFnPZToJ3UErRApb0zrPoD8F0YON+KzDYsAGr00joQa+J5FB16OkqeziWUTXjs4BfudB6Mf9qT
RGtgLOJ4sYyoPFXxejvkMEJPn5eC0wsyleAs2GYRMYD4Aq8CL5fBp7sU2SbsR5jhPuPLebE3MyhR
wLoliCbp6S8bFM1ZgXEJeM+JaDGny+291OAp8LsdWYNPYtufA9YRmNv02/MxMDiSrS9oENSt/D/5
AMf4VadaXXO+n7HEc7RgpzV5dpwUjGenoXL4LBUlt/mKjelge71NbS1ez7GxVT++EYCdIx+PnXpR
9vWG89E7JOfP3kITK2o7FjvRGLy1RXoMEs0Z+NWOkofLuFi0SXOY/F+wuSukXHX/IVq7l64XP7K2
NNPLOKmDyyXqWTLVafLDjdbuRkAGVzDzedjBswdAuOox1SzWCEazp5eLJoALCpTUczBwxMjh7uZv
eBdhEr3HT/WBDqW4xsGyU7iocwek2Fm9oFnvlB21H1CIGAbDZIFws2st/BjlrMB28/uRwts8bvbe
KGBeaTe4hrorvIHMOGpYcMCnxpxP/gcVM18043dDzcuqVe3mbkWKHtivYkcBUNeTTS3fc0eJrZbf
uawyCgIyesEip6oBPZoUB4MojPn2Dl1QXvCyq7ptexJd7NIPRg1sYZE/70sCFgl9DG+R/uFkK2MH
boWQyw+as2UFvy3r/cUQVJseJnVETF0l2dI/Mm1mRDyy3lv5WAllfJOyuyj3E33MXA++QR8/OwMW
eDFLxzyHDnVQYxAJOfeqKEGB/cfWRKRx7MJDLxNoaINqlkZ0LaCPyWst3vNTtu4zFlAehXIdgfnU
xc4rTNjf2oLkxmwWiH5WHzf2qTqENQeIRSV3ipKs2N6b3jVIIjpoi8VS2rSx1gD6iil6AXzSQIw5
dOBXjsxIVibGdt8Gk/LB2AYTFqgPQnXhJKqnKVX/yc1++d4VALi29YrEXHKZLagGiNJEKr3YyR3Z
sZNKhd1uwJwIPFjah8S2c1BwoPD7FhXgQpS2ZoyyGijug22HHhGJ9Dy380RnviwsVsymhx7n6g0o
mth2l/Z2jJC/iKH6DByoBzrFWR4UzmA0atzoD/yfMuStXzVy9wfftycaARnhrZD2z4McKx88priM
Vidp3ZEFrFa/tRE68M7GU3660mctz+2cxyD+q8Wq4BJPbH0Vuuu6vynkE/cQam8XfwaJJyjJBMLz
hezHndLtkWmsgqXT8ChwftRspprukw44uNNT9IrM/QL64hwUe+43R8LcSAIejIShQS+iyfwav26G
ouLHKENU+ziA6LGLs0YQTAp/YLwEae0wW0qCzH+iU4GZE/NZtBaretEpgYXyk8hmBow/KpLXXVfg
lcGQb+vklwKhEKQFxtPa8ypNLjgQOw9XalDOohta2wCs05oMmVhnvSzSL2qtzdcTEri0IxlVioBp
3TdxnrFtAcS/GWMkIXE1Se2E/Emd/UHyKJCn5lLtj0+bY5atGZhxBLKO/C1iat8tvE0zrMkWsxPt
XRx7UpqNNwZpJdVfhjoZNmUoFG/NZM9eZ8JJ26QnjkNV9uy9FTo3E874XWAD+MxrAuBVhXsktn2F
hHWR4AJwh+BJVwY1niK1Y3T4nNGrxrmuGi7xFAKEW4lN2/ojOfpMv7GB1YIzczRlchTj6s+xDcZ1
zbME+M8Im5On95BpnW9mxt6Ysx0WO5e/vb7PQnH/aqkXHfNhZJlNbjVOD/Fpgm+h+XXi4q4MrfnB
++lE26ThzHQdWO60GtWrcKKo5+9oE3frCCbam/vrhGc5F/mbWNj9gIvl/GyM8oNrpt6viDZxeafq
WbQJLprLfNJlzMxxqc28SBr9sJFaHKAd2MQSYHGJK9uWOEBmNRgDvf963L3WI679RoyrxFLXN0HK
saXYIIiAidtaFJ4j+6pP9SDmLQsaGrGSECy0X4H/jERxRV49QqEA18AgffP6jO9CXW7iuts229pc
0dxD1UM+jRnP1oi92lNO1G4cSuiQnp7qAN7RmwnHS3MdIJD3ugGu2I8WzVifOUBwXuS+mxUVXQcY
N4A3xyIOnOTMTM6ldKtfkY9/nC1pqSCKSuk6Of7Tj/Jwn1r418OxEg4UvBmlowB1E6okUB2hGnYE
RhW6GWg/mjj7k8AqZW1haYVtGvMG8r2hm0Zl3lWUy9ayduxsMTAZ1B/QkQWc0LbR8BuIpxucCIVP
RnJ81ER7WGv58PFKLZhrzi3MD6NG8cuE1zticeatzPapyT3LQR1E2QI998OsE2QWXjJi9qblzErZ
+WpNJ6szmxI17AyB/BZ4eHlVmwbUvCyimXOFXrSL+/BveaJ6CzvdLzxB5Rjqcxb0ZZl0EU4MaBpl
7ykQjlPzglphSWYpEaB8jK6GqyzYi9Fgnvzz4bH6xflHBadqB64ftdtSU9DhDvHyxfNPo2mv/QQs
EZoba51d+xi/qAKgG3acOvD7P04CcITeqqns0L4siol2PIQU09ZcwGBdnuokE71HKw8If0/5jUw2
SHsCFyAGPfMYmA6z9CjlfaGmzwmOIN8y2IAMB1MoiJhMGS5DGQZeB8QMAK7SER0iNvK3Jb2c7V4j
53smMtZyn2VBqe7SZIzpBTJ6g+QzqwvEEQwzP3gvVXxZbijVzr2u6yz8Vxs5NVXR8O/38UN0pdk6
L6KHC4z+Lybaf6ybJVP3oQUjZMEpExpG5YGEC/Eya6hYKd9+GAIJjxAQiPecnhJGI9i43yaUIlqf
nyis4sUmVsP1cH34Ea73qEjgY7RsDiUes2ceW9DaR5pduedxqTU3zbGJFYNNRhg1TirhQly+BCoH
eGVBvJknmQcU6PMfhCE8nCoDzHHgu+UMkCF1VAaaoGEj3YGtC44unij+0jK/nMXQIvazHJsJC/7S
DOgg/Nn7U8yVMTzzNi1V4HK1f8slaVHgm6DeOveEobA4d8vMmzU81o+JQKepWq9hr4dZ0aMaft2Y
y93ExPPd+EGl6ISLMk0VJbhSoDrt0FThqcD5u0Dpws3j+Kg+HIC7FPJE/AKEuBHA67u43LDCWOcA
CTU4bMFgAqSNVOezVJzYAyDcBj7D1FB0aM99ad0tODPi89id/lLbeOUiB4TY1UaLxNlK2DCCvKb9
odB0PmGjsXOasZ3cQE5huPbgnbNX3oYHmvHgjdZJaLoZoptSe9KhLbAz90h/bR3UZTgN7TAr050c
I4HM44Pa3zLx5s6Jho50EUO2r08mn6+qClNjBVKGLTPEKIxvL2mtRdGGWT1rVgBM9Qxi07MMaFJa
XlSm/CugsafzZwRLfXTANkH3Oqile3pJ66MksKonX/rdg3JAnwKmtgGcPr6NMfnaP53Xk+qnvUKI
gUVjYngpEInxO6rD9ajr+uk8ww93T800EnAM7gvblEXPch5/qX3c2j6uYnq9m4gMXTlXxIXdQ3vT
8ENfnXQmdYfAnVtYemREk38IHjpK7vSjY5dLEnfh9pFM13moPzr4PGkd7y7JUPnTDBc7PbYVIkEV
xp8sKxsn9q9aRZQwdZrXL+bF088mo5Vey3K1csnlLOSvwyOiLF4cdEw64JNFfKsCQsb5lsED3D3x
N35z9ypxwfGEoBDz5ex4HedSjnLK5cFWEgHvtM1Qjg8TMgK7eG5S2uL3Fjxy/0mzVb8lGcf+cnAL
LuLdvgrE4NgHxiK3kjaPZewwi90bBujk97c8emh+EgeQgxxu2EiH971RQwDVeOT8wS+JNS8IZn7m
O2U3dQhUDDahhRcX/OJGzk5oYLd7WLDEhuioLYV/YPEUtPm0t9QPjMppLaQzdLiYyp7xYmKaXK1i
93O8mi0DOmsZwcjshDTneVffDQkVfA5rOCQANVedgLJ1hG110wiAorH2jZ/d7dTujI+tqVp9gfW5
FvHhgYtZW6+8uShNrXryQOfuP4TNrAhr0EBT5fe8nQXZDYfAyhht1h4CYqrU+0tggXPc0yfPGAD3
gam38N2k8rNpgfum3Ka7Uufmz4ytF0xx7dqaRZIZo+JlybjVsF5h0y+pSlQcAs1gN06wQhMV9a56
uDH2vHnjmN1pn/4vwFjj6d5RtP2KsXj6/US1ks0UHB7wY3XLNctAqERpuOSbHWUIruHwR+5SdGDw
DO26L6HWU/ZANPStXK+lfTXTVxcAZr3HGZp+m2vodLOMNqQ7ub1PwN+YU6Kd06/rHAL1Q5Wr6rJa
uzGGwO9rqET1O1KmmWIJKoNpQYggKsw0OXLr8enQd7EvqXhngF+Zsj/chzdiUDORQwdPUHqnHW3A
rS9ZXoxtKsm7rWBjpfOn+OxW0Q6c+N0Nu8WlEfdTatfGqCx57zXZLb+uMd2+M7J4zPYIQyenyTHN
PO9TByZ7KzXzF7jGpnDs5dSm9d3eB5n21EKxdDvi0faRy44bEPdz2mEaiW9kQ31uG/EvmuLodudB
wBnjerRcX3zYKZsNhzh6orjYavakzWNAI6t1rC89B0tG2EHcDXN0E+MaoFHvaEgwnbOmd3qnh6+v
Px8bl2u76nDwlSQdjBL46Wo3vQDa/4O7ts7oMEy48/Xw55ZgA8ABG1cJM4GhHVqAhxGxv4zkwM9U
xbUGcbUEZ6NnyIYSXGCfURT9ltJBx2vgRcXFIYyQxdt3sfOGHFxpX1mcIZ0nvoaRzByhHqnk+5Rm
m0XaJ8w3RZ0t38hV+20e6+a/UHABK0M0fJ/m95BJ5PcShnt8AzdCUhDV5adfNZbDzMbTXB6mzF5T
cVzFL5T83uVNmD57Yn0X343vXGiemTWRaZzFrAVrSdHPgHxkq8eUE6jRKoeNzGoF0StTKnQ9DHF+
g1/or1/3Jbh2+FKL8rkNDq2y3Bi+2TnEdoTo4iogijs989WySolaC50ZT8MJnRy1e9NHOn+Ek05o
JJzzee42VKzfuwe6y/eigL2OT7bOeX6s3KJnwCRkQ9pC5u8aoI/i9JChII+BqWch7unn9KWjCMvU
JxeW8JcC9OVQpA7WLaWZRwYM/tSZJNnzVeFcWIMJD9YT+kqD0anGoYRs9xV00cwdRpeYO4zb42zw
SBb3ZTolLSyyVtHS5xv5fd/7nCiyeuiQeaXpOs/cUENX1bxk6sCDUSVjWFL/Xp/wMGT0b/kM9Dn+
LIg16u85kMnfw+/MFwFknjSktPVzpRbMwANXJnwM0aZ0Kyx9AlbUre2IyuovCRZnDZuNUS/Rtvmh
3N5+WF13o8DFWR8F0A8AbZhUJVHc1G9fxm39PSx1URzClZwz6roynk2BPdDnWWZLoHMT08pQr/Kd
BC+2zQZ5BsbOJeCiKJOMrbMESgzsMd0eCm4CvEhi54iF4mY2t6YzxxaOmEuQ6D2sgo32KTsjEPKz
KTD+U0IPIaVPuo6I6ALaa295AlRP3m5D+U+Ig2WyOPHcjCTuSqdKCdK0J3k4rmHZX+c0KodCXbkn
MVoXL0O+AI1C1jmcR8RIJPzMjnAiCAKusoXc2hygTfWiwdDZSZgQ9aCMMlgwE2d79nhWZYa5RR7n
lk9sH92Hwo/kqybPxo79manGf8g1aEk1PLl6CHVA4vDJXnS8v1wAkftf9KG01EiMf5OwDpRxmL63
I85wZxXJI5F2YARIKsLjWIP/nW1rnpGJVUr4yGtEWUKZGoy1UwWT5GV2P7UPBRBcsxE38AwR/R82
qHNWjyYZrn3smFF7gJHrU81C9SldqqhEKtgXk2TczNu5RWdacYxQ9Rmn1ngCVVuqx1ytczfyYGqN
84MOrhOu8BagSHjUU+iazHE3vBb0mXq1gp9P5mvpYIQzCSEIu3wQXwATB24RWWClnK6BniGi/5+C
EObskTpFcIq1axJEJztPpFoaT/pRRJkdZ5MKeLV/7h4OffMeEXGe1VBGQua4SGDVUwnARO5CyzhT
aBAgdl3PM10kxixRNoeD6Q2SkRf3sSsLb7kORGwgBopYjNteFI1k4jPtpcBMArASFsEGRWosLdnS
vYI33nYKCD7dnicMflEbtOiYmRIKJaftZTUvAnk10YTXqmYsdXktloM+xDYldcRuHJI3sYXtVqOA
1lvwlsa0Cw3pAnoUsIB31qExtWqmM4auvvcj0IQzgyBJJCgJqgeRut6yB4AHxNnEjYcjGWTj1za7
kOnyiSD3cp/+pI8K9J7YOouTGwGEns6/GkTBxbiFJ/EkMCa9208lH6w9hEeDg82ga7jKSyy+8Su3
JX5hWYzsxE2MWsY3GDKyYva4bCitoA7g6BNQAOkyK2yAvm6gahJQZ03HU2fuqZxFl8aFOsVh0ujM
dP4buXFZhRHtj2EbvrMcAbY1F2mtqX9FIHMIWO9Phf6WMMI23NQr3EZS+yG/5mZZCvHItxwMIZfP
xl5u212fS9i8audZTZ+Z7ehRtAdMZxkapbMnmYaZDb/FOIQApaJ4GzcNcFdC8RNc8911mR1Yxe74
Dd6k5NA7oXaqxetudfTy+aM1b9PLLRNRk6cdtG7JQtlPf3Nre5CY2UabH37UnxSW+FDler9fsed3
cA5XYWqhqOMqi2SS651ZyZN57Eh3tMa1+jQ8nQd0/ajL9rZs+4omCM2mwozPQnhW50MYqhhk4hyT
sOWwDDnjoPb+uydH34AiHJC3o3pw+GdvBXli+/UwFyuMSGWjRjMIc8pIx7QDkWPatN0DY9CWucqB
xUOr8geRcgW20C7JSrNaMlUqPpdnJaYyk5SrrXyjsqe/la9MvNPRCTnnHGDwO8a2R2tlJTU4rQyL
dW2TE+KuHJaMfGohAEiBvqdZS+ybWFzDqvD7Z630KGVBrVHqaFqhWyQN5XZKj0LQju//1we7cRV8
TdOVAWfrebbZHV14x4p2jtZ+bGvIe/0421Q4oAizk3viY7Lq+y/MYYVYSP8TZxDYWjj2oGjwk4hl
qO+3LbXFUKYhF6mM+kiL5WOJ31FdE5f/lPQi2PwtRPnAEDdi4cyEi45aJkUgz/T3SY1oscEmp+MA
yHRoKRbmmW6ZQJATe9r/Znlm9E1zq9x6ZrpD4+Zl9fIDnU7d4hnq7MtgMwnaWkqATpjM5bmlvIYj
t4EAponTNH8338g/d/V9O7JOkUQwObI8spRmO+3Z7gDp1OtgYgL5Ox5A9+b7yrdpi53wM2d5CQfG
GZxLuBGi3YRepNC9AYi9+7703m0+ou0tjvhH1EFF5FuhdvXA2DA9Gz0XrH5yed1Pw4/QxTyYieSI
fnID5tD8oiDr5opAXawbBPZjxbDbex0uMnmHKJvp01Pbd2k2FLV+GJuhq+drCYnobdjxBGjY3gXU
emmv+bTf7nyUZpRF7IJPMm/Xf1G4klHYdH0H6VL0T4sNKV3TQWx2QwfEmqvYRO5tSrsqHNXXt2Vn
Jn5evZgxE0MucONdmHdmg5sdxerip++sNxYhBcDKuVYjiv55872t7IdG+aZnxe1PeGlW008meZ1Y
3kCOyXWzH6HjfcZocL6I4UXN+0vOBxrrXsEO/CeAahUJE8GpWfVaSr8nDMIw02c8MnZRNgIKd7uj
0CrYTPX+KnoefsqA/ghopflQSD2RsKBm2Bub2mh3Nt79FfirSd/YrNz/MzzZH2TVgLiyaCmhJP0/
6GLYK4jKYVtetUbuioQPbGBkdeC+9cnPjLzvNL/82yM6Ry/mepnx05u+3OeQj4LbcqVfuNpRw1fM
vEX8V+jo9s7NOrY5UQXmOqzVg6UnByl0+qECZ5H8ZRtqmPw4nTFH3N13Uc60SHVNLT3aX28VRJVG
9XxpyWXlq3mXQ3C70vi5hTFH3P46SQpWE9lDjCncP5XkhJT+LpSoiAz/8QVZEzPsPP88r/xMZnvF
xNgedSbdw3mfedMupw4bXwpJKhyrgpl0wixahk1srwfupDAj4rTKXjKtdGoMsj7Yk7kq00jZCCyX
ARIsnJQQPn9zWdlXOo2H7NVW8Ch9xux0bavD244ZEH7Du/lx7nmKo7YRge3Lt0Er+BQ85KNxAiXP
1TpbDMUnyKcIiiIw0F0R3ujBPzvQZQzTOBsmu4cOyw7BKazojObGSz4RNzilrQTMAPM4EXQj6QsP
OAV+ScZvekjQSac3+xener56WNLY+jVjjM0XyAClox+Q9I+mEdkZcuoQS+vdql+Nk+AHCi8UB1xR
cWDiazQttnS5cHmKqUQyS7+6P/QNMVjlflWL/tkwtCEJr0zHRGP9xoWyywupP2vJi2Z6pYPZ4gHO
KlTABVMsqYoFdqBs+YKBwEXQOvBFViV/C5ECVm2MA3ODlkqm2EigmjX8SSElEp3JFw2JT/j+5CU7
s0SBavp3npVrTXEw+ANYeEd1cfTZOrUXC1CmPwL2MMVaIIYmlD15W2DRXxqu5vSql0FPrgG5EYYO
ApbnOWX8HVtoTMhlAsrnLlToRon18mo5qfdpnkwKDD4GU+02V9FzDteXKB03xclVW/EZNKEcQd9I
E5UtYQvTnYNMPEaYwx7HhpoJ0CkvAWGill24ttIGaxDYDycRwTIYQqAJj3BsIXdIZhnEc8nFBKtW
ej/rEH8XhxreuwwNPXXv85MLvVPmss9rLtNOy6pzgA5THnKWFzl+Tolmpmv4EMXj1I8s/gePzzJL
YqXWohH4p4jmmM6JuyjUbXbZR60eQgrYaC66sA29oBZtWFMCHDX3uJ+WMpj23nXC+fN1/GCyWpjB
Kf+DeZTsCM4XAHXRn5hHZWY51eAd1czx2VmyaKkYX5WMajWucQCz7PpTr+C5P04e0BMnyZJBdNu3
tmKo+x0d490uBGGg95A/EspRDTgbnze0sffl6yn9DmJdQBWnnYxi43WtIaMr1w6qPnazuCzxcK+V
/TnX9ceqLseJae7RA3nQJMUk290bIf//eBbWWYmTk8lHC6ZOmKA66pfo7NiUMKdLjwII7GbJ3F+F
UCFzrBoSXUxjmmjFo4qZcytMVG7INvQpaF5srv0TU3rQH3QjJVL7yo8xs6FNXCbWTGhglUH8YnO6
u9tLp23p8U7cfb9YP435IB/0U2D10Ch2Tu3J5VNh66v1N9XvnJrAJBwnaN3+0+Qh3t4B+4v6CRp7
OG2sV0UI6Zyar4qh8qRA/cDyg1/YCiL/hVUOLIzc7XUdYS2hPGf6N0eFa9Szvly5z2zwUm5Dl1o/
cZ6vo8/iefXS395Zli32HF6Mne4UuZyJ4ZVWkPscJGlBIk7gfxU5AiNakWs6IWSzC7Lbye+PWRTw
pTKzCVxBxYxVgzjJrcujyBorFYZxHPfx+ePkWKDdztKwm5NdAWy7zUs7J2D5eBzvyyZY738Yb5d5
VD2h3dJWSqADuMldgRtrdJ87QZ6oaScyGn1Ip+3Q7iKiJvJZR/YbDgzLseIPFnO0Ayez5PAqn8PN
Vi9OUq6Df0QT4+7QMF0DjhmQHFDUfrG44/PkqNLLXGsRX3tmawnOnVnZv1tKEJXfEhQ7mCR0nacA
Ag1vjZa1R7VyD8RAu2YlPNi/L0ePEFr+lPB61Cx45ivazATMvJmZvfdvyzDGC4b7KiwGzbX316Gs
Mfs3AtjvZYg5fiXUwi+7YqmyvHAsdqQZX85Oey0D8WTftKfj2Q6cNgsCTTYraoD2o8Pe2N3DY1lj
cCUh+AcRf21BpUI3Xn+KJPOZu437zB7ubjiAISUFJiDeD9ukpi1M1/l42VeJSA5X6aITMmuMTO6w
WsThk2g3+s4vYFMir4uxi2wXghXL1YFhlx1uCLOD2cEitD7hejYmhkHDETCv9/gXechmpTelN9f+
j9jk2Ha0W7/Nmtq/kbnXcUzRFkgQsiMJ3m4L0aPm+Mf9ZqR34aAwBG9tzy5+q88aJ/mIx9rlcz9x
7wQdVZKieA0LRTwDHttysevHk15gK1BVXsORhVx+oQpQgV92paphCXkqlGFE9akI2T7P8vbPIBen
8FcDkUo2u77UvFiYP+7HbmSmWilzsKrGWHWiWR3SOOq3hvnSjB31a703bEraWak4qkx6UKSyrHYO
NSrwi8tYQrtnTPgbSzM6n6yFCMNCvVTB4lqzS2MCybtnbbvylrCO5XyaHjb5GIksIU+Y78LjHtsh
yIS4gH36NG/IcFX4EkAtvYcMDSoRUeL4QpuAcvj29eHX+8uSx4yfTVRWSdpG8AXaTkyk6qr/U/s8
ix214snVC9Jv0zi8rAwyaWDv6eKFOKhK/CGk1CXLyL8NVdPrLxOVpk1pyFjEydN/9OXg+8g4vM5w
16/h1nxW8W1FO8f5m6cqtZlKWuDRgKFxgWaqHGMKuHpyIfJ/dTPBUhz2a/Lw44cJZNHl+IfdwYHn
agDlgB4s9rn05WmCmjeccFT2fVC8Z3hGsfBif/abIExGyy5yWlJJhO3O799rBWDCzbx0MMZjdnY5
Cdsj3qlSR28dMlS/0C+lCSeNY3LIJ7hOWcqIw9o+XkjQd2aMi+pNrK+buThogbTpz7ahyMlaU4xA
/Jc+e09aMXdXxpHr9Lii9QjTPzZdjWsQKgVLNfifvKjwoMyWjRa8cSDIY1VaYXhoPq/OqI8nBKoN
L4BAhTMhrQrYefrRpHwbKLvP5Z/VfR/st6SH0BqPSQEFUfjnQWSsewdV4Y+w7aVZkdZIi1nP9FVs
xbSAL1SlExnN+ECkytv3s0BvHo9QQgfghuWnm74jQBpVPNc4ghZ2ESa7Pu7Th2Gz4kxjbABYMBM9
PMsXXYAirPwjzSKFeqeRCTFtmpraYlYtMB5Pu1JY8534eg3yL6r4kigPW1qeJjUxSXimd7UnCgzP
Zf1BA8Kh4x3Xh34dGUKavfFdLD7xkV8JDSG44SIgaMB4bBSu6Bfcq7c7QLOSdBw2v3s//b+xA0v+
jrI69LLyWZbVPRSVVyppwdEY3A/UKG63jMu9PuB2wgjaBkKA5XXIsmK9Qt0pCz/uCpoaTSSJbbZT
kDUhlbapq/amZlZENkWf1oCJ8dIaE94W/KDKJgMbZ5uOZqdGpKmLY+slGL7Tk5/eRTwJPSa+xnBD
Q8x2hb5RcGtu46/B+3WO7v4XWo/FasWm8wdVPINZ8LA4oXdemXUgM3ZhfC599FpSL3MAzg2fV2rc
R8l0THuaTfZyrDetJrO1W846N02yvG34fKkb18lml3ZN1tTurjlEOYbYDier8IR9uzWG5hz4Q3hH
7ypRh+dz+EtayZvA5Y6q5IYoBpnABeWitK1cVGE/O8ahXUVKfx7SCUMKLpcL2bQkiNi63Nz5QVot
uHiUN9l7foRflyqICeuP5VyzhHOu0P72xZNRVzrFQe2rrBNKFIxyywHJMc8ve6GPllvWuyT1B9Ey
pn1CnMOFlTJOs7zpfzIiWNxUevKcUIMYBGkYAy/MXRRovoMBvBIZknqcwelnVLH61PDOo4mRCejW
mmhZxEG+pFFf1kA2hfYEDfd7yfrHoO5JWYDAylvU7rMQo1S1UiE1ssnZ4yFk9TBAbg4aeyZgfOIe
Otd1TWfb7W4vW3OTKzbKElHdi1+m6ajhlOrN0yOnCK3r2qvRX5j2naoQrLjbLxHy22qthAOmXbpV
Az7YOw9zHyXp5iiPoTDdVVPR91g/t7WZlNRc82sHAEMkMPnnQtQc/pgqw0qko4PRJIQS5Eytj5VV
x5NHEYr964geYBZhoZj6nsuuztVSAw27wc3JiMzDhMAVpRb06MfQELTqDo9PE390VEZKwLTdVHyO
xYIKh42DWWHW2SZwA8nBAbIXKE5cbUrqVKBjOPuWAWdqZC4H+6+WDp5gQLCgY/8HQoswaqbHHkm9
jBBQWYaJMm0qzZ0QAciXT75gd/SSddxPZKXKoSRVruBBaLwRHJgKvsw26hniTfnlHoMUKpQNY2Wc
yDuP0cgBy0cViVOiTtFRAhh+ijgBxdQKEk+XJF147vVBJHNk0UHe3lMPVfY/YMi6I7HI5XFguTIQ
0iygh5mwQr+0A8FDRWmj+5n5B+P/VgPoxyGvS0SbZYRSYaJnwm94CGatJpKZeXLXZ7NS+A9laIu8
7BSw2AAFiqq/pCWSYMXyq+xfcQfsC1bM2X/gHPp2+lUpOmcVtPLAhzVEfJWeB3kaax4qDTN3oBMw
OtRZqYJKEnXbrgq7nmizRjfe9Qwcj8IORqYDvOIw89D8DwW8a/Kedm83Q2TrdM4mQZ0TDgs5lA8w
zuhjDP5DIPapVNQ+yTPf0UDgzSsO+UC0AaDF0xeOoTPqeAOmgYFR4C7IajhqBOqPBTCk+VWOxKL1
E4oZb+zfE3fDvZmoZs/ifpKMxd+AdarUPah5kdR1AyH+5iLoN4ZLtn/E4n/OkbRl9vyb+GaYPFWQ
PtsYvOct8sfYPBDjdvBbKEpOWx7U9cURJoLcfVoSWa2TbJmfd5aCGSSNUTC/gcP73bGnPSQiyXkQ
HO6Q7KtrQMQ+uJhAdZ2zXYo+MEtIyUfvNsXCyPLf1gi0ueLQIuwfnMlO/r3N8BUtY/BrcfXKQ8B3
XaNH8Y8phbLFi3lDi6M5S7m4v1hNfycZg+jG4xfzyywrZawsLXRV6xbjUbmQXvMZBn7SKSg1Ybmz
qFYbtkV4rd+jaZUw9NkqiJHGgi/Pz2Q/LEGQifxzHQUaCaHn9YaSQnb2nqiW1ajTBnuIKgvivNew
ICKOjJXaWmBvP3ZF198vrT3xvExZWd/itP7aC+4/SHvfY5z7v7Ap8W5HKWo3WDL1y+C0f+MWgWU3
i6blunDxqCdgD+qo11li+bujUQBNrfrPyNfZeEDe9XP1VXFXQl/1tDBr0CS4Gr0BliJl22wPXatO
JFqn3DOnltqwJ6WUepqbDoqR2EesUWCwIEtjpP/4G5CnPA2WAwHwbeFnzxEj6ltiC22WennNnvk8
mBYUQeOfC7+qFuxDgFYrLtfsnQbPnsMjefC82SRSjPS2rMv7zSGPY1uiqlISCpXLaVESoK9+9axI
n0/OGTAFOOuxDdFyfwpxsdjaDBVlttE1d5iuPXpKYQrxP37lxTURS299yOYWmH4dk/ukEOFrKU0l
Ub1iYX6CxKAQhwX41wDgGuagIf5MbYgk2T9aocbWcnT/w4XZ55Fm1ui4zQ+o97UDRw0TnJszI2NM
uV4pOB1Uf6mPhUFuGYZHz6Us8N3p+DYdenTbMR7ewwSwOFz9UttT8XtBN9txJgDJUlnFIXfeNWhE
EMw/ivIEU+CHBh2nwcgRkT/PZ2fRTo4dQpKI0mTekpNfMWZ6xP5Zk9e88BtvyhLSBhl5Q+z2IBwJ
6C4mhUb67OC+xx/Nzq2uF4ijDyy/IEQ4FEBov7R09DdBVLach7vYAfTcHHD1D7aeuTmtvQVahVG+
xbFpvhTO+ZfEy1/qEPuFPVAT7yo+HXt23QEUlcWNQdpSuz1tSG70iLoZs5UFTY5KiNbucwUNqYpA
3R/U27lQFDzxGQl4pdzJBvzGiHaRgxJ0TgPpwYtPBsUNH/rBJcqJ9iryv0UZIwdkywN2woOAjv6n
IHENEkN4yuTK33dwE6mEgm3v5HFXLshCs4ZEsOtn0sBMIZE84MqnL6LLiMpO06fFPAQPrO4CvPTp
c8HRmHnx5nSdj0Nfmh3DdrBcYrdjXxeQIKl/Uzku9mt1XN1IlC6jBU1E0nNByq/vL6Th7psK5Wv9
Rw/v+yFUjdDEhNL8hd7mPSv2KfXYqZxMXs6Yhu0IIh8N494BS3txOnPjgPlyQlqjfFD46WkhxfaA
AItc5Z0bIGJYYnQc6XiD43iruihn8nl1M3bEwNtS9IrqxwdiLcyHEEo4+Oz6zFlOyTviKkzC/9zC
xLiLA1fim0jBI8keGC5y5954kMURynaa/1sckRCdbBlvVfAkMAGmlUHm+XQWb9Sr8z37zk9+MUm+
G3A+r9V1gMLh4PH36BwjLj1HwgRVKdnfoAGbaqBPvjyZVDTqb2ZVNOCGh4Bc81rDe5LKdOLNxARr
8qSjDL5ez355bLufjUbBkJdA2yda4/roMyZ4auttiheCDEU7QBiz0fcM/NgSO2mkIZIHN3BM4jc7
6ndOfIku4nsbcU8bh4epp1GwyqsJhT/j801IpKxUAWJfYzo93IXu/GVLp8/nbGLW3MxsixXnFRjb
p5zQY1MQXrsM9LEEI4IOqC5bm8UCzbJCsMoGou9oADeDFK4e6YvOqW84IHi6h/xGMew4c6kAXX5C
rPytbxIfHLvGDCmzPwAJ9DFiuOYhA0uApDB8+B/WjA+m3MRarx7HMtJP+vW85TXQfwY1WvdXMb3J
R1tsxUj6rpiW/YT8Tqfrb4tdfOGdv2u0LnPd4r6kZal/1Yh2pZF0I4vr6HSwN5e7BbknTPtH2n14
tY7IC0VlDw+XfuLfShOHRxtHjd5Sz0U4+51I0LcNipk2vztpxUokMU5XRGi83gQSw9t7f/Gbsirg
Ov70WItk40S38nACzU4O4KLSAm18kC6Of1G0Xt8jw5KZfc0zVAvTW65BOoJ/yyW0wy96WDTHvNEt
7Ve4NUOhECSnbCiWRLMgaaP2xFv97P4HHiBzMWneH90mivbMXMGgFBy0Nnu/46Dbf3YgXydreoXj
DAwYF1aVHn6NaJECrwzSyRSo0B7rWSGAcvD1c/U+mx5JUJ6riGcC0gg0uqMitWTvF56qHR+aHqCI
yiCRUrYoVJgW5ublt50FcEONr3Xl82N14mI2VT2n8o5j4fq3m7m6tHetjwSoL4S1jzj/7atx9o91
4udBKvXb2S8j/g3QmUOsEEkWtrrG3xNWucJy3/l2+fQtOTWP0c2YGFZE11kVQANH8Rbp/I04b7kj
6kkS769Ytvu+8jeRTafPsqtAqB76Lcb4d30k7iNuR0TUUD04JeL9czA27ypO9NEVthFkOOYu3NI+
4bWH+KNA/Xa9OutrnTPI7YPyclinMusuhuk5wbiT66LhSpfwbPBn5DU+sJu4njBvUNaBUHmb2O2Q
UeCP5CXEMi17n2TAUgaWIaaoiBacHVDIuuGTIa4xxXsJPQJH2MZGUYTGSFMphUsO3gseAhP6Lsj6
DkYOftoczvSjp3ehZlTOfp0f9VhxWgnUeMN6RFO/oO+r+wwvUOA4tSc1GHlERJ9R59w5m/KNP2iG
IK1XP6HAMMz2FyRGYNb+3yosM50bmT7K0HTa9OiwDuG6EcgxmR5tY0FYdtRI8BSXWookeeDAOXjQ
/krcO1rPoLe0PIa0omJpY/LdS573nMdnLV1rT1/Z5i2exE2VKXifBr9A3U6Hvu1hWJ6hXn2g0yYz
GqcdH+riu7PLTbxKweEOwkjH9HMXBwDdWfyVWPVItIUMpFtnQqOq436KkEOUfdBw6imZI9DXJp4+
PBi/ECl9AxW1RIZGIxEAylKQlKIrvXXXXfBKuNr6PGvDamcL6l3hD6qh8owe2Gc0UywIbDNA7Iz2
pm/R0t7iti7IYotZDdJutkXSnUKlofYO2Hd/XRFnVb0taGCkmU+MT+Zq9j0pylHxKLcROVfELcFk
r6MQkQWPzygT83WP4+/f8ZQGDfHL1lfjQuv7IR6tCJFYuG7WCrP/YtMH8JWseEPXsjyOJYwgFvLF
0YDS2ylj7pJXVg9G6mrNmKpDfvTp66IVsoBGKopeiC7wNgxRCeQzzQVWeRWw0XSSYoG8umxzVyMl
9K/BTlASUdaprcqJiocM8+AW3IH77NAM2hjn6O/mYj2L6fG/xYjBQ9nvX2bVmo+5HS/BMJGPqvu3
QuIIP8vXxJV0VVj7xNf7/cDLvWNDp1XT/KjhIr/Fq0GzlZHJ9HGKb2HVQxg3CnpBkWZB9gPH/HRN
6PLTvhTxuby3S2boVmaIJDBMV8c7lrAqc05Uu+gxBrARyIndjcc/1QvxsKJ3pyRXFo2eD6geDrP2
njt66PQfIh4f9qjzp8BREmni472MmwAWocsWeo6D0H7lsy2Fd1qtKjYCiYnS4D/zhz9MxJJSOdVQ
dW+MWUKZPo0kzcTd9NMDo1Qa4iKF0Mmlc09vGLkgohR9FRCw7ag87unkPKQI23FsauLO4aY4Zurb
OA84U8gRFyTo1+xzklq9L8oBarK5MTpgUrx0SFI4c9SOz9AIGZSDKU22iwzHRIhXp6pml6BikJjy
eCuUfnZWzn/6/P/pgPe8z2r74wslbkbGJ8AO3nronma6B9uz+BvWrM9H5Qu3HgZQshrhEX06Uwjs
Q4VtJmIgfPW6lWKfD4Ls2shszqKV+UcDN0dyshzeAC7Ce1emcZJ8x387SzZZaihnpl3hLh8tFTLU
2o/Bmjd83k6W6Ar9RkODk9TiS+YG6S5bQMyfyeLZciqmyZ6mDezrHxmNOrHeANuTHiUSxjLsAIbn
JcNM/2LG1J0tBYJBRD/BXsv8UPK+2b5cHvpwTVyShuvBF1047beFcLD/U7sZatwtRO3c1F9YlHmf
/GnosapxUOLe4BQAxUXBmR9uOmxfiY8MUt/8pAzYrBntCDw6SifI0HxE9EuTY8hDD6X1LoJZ2GBJ
mWRmjC5x2+nKlL9Snxj2dfTC5E6zNvmp9cumIBLojLGXrY5dcm6wI+pd8bY67B4+l2G0ydGrVf7H
DGjJ6PjHj+AadfM+slZTBUOAy3fRV5NvoqLHtIOq1pgRRc3f4uMps/0D7BYcnew3cq7YqzkqXgtD
l2jRuJnxAOIYJVPsNiRv6cdKjiuN9JmQX7QFB8L6jTcXhdL/SRTeAvfYNgOIb1VGr+f6/hA9wzgP
W+4PhZdbaNGRIl7H63Wk/EHvDoqsd8KHKp1N/N8ODXT0P4NEikY4g51RP3BrMClmWBgKWwiNo5tk
oqlKD/+wBdsiRZ7+2CExtA4AFm2xZa3ep5KI+5mpjF+naZO73KGZ8Ye7EpaVibCBYeyfRORwR85m
U+4zbniXJm8A+UOeqJy9AjB8gmghC4jzlhLyEPKJwMZNjormCFh/8R5YRV/HiV/qyk6vf6G4YKSG
UXDNRvGRGzO7+elV3HJxXVX+VjuRPxLmQoFMDsnCsPpe8g/xfjNFCc3dRmY76uX7f6TKqymEy/1d
+zTdX7ok5Dt42Lz6No/plLflQsMlx1rYYSh6+SsDQJhkQiHkD3cE0rkscqwZWIdp06jy+pwUr4Z+
KTPPcrpnDRZOfVl8k7pqIdzJxQ1bDTXza+Wtfgy4OEcMnaCdlZdn2OiteSf2/7ouBdn6ypTvQusg
esSs23V0kfieiYpm7ywXCkVGLYN61yDBIrdd+FmFuWM3DkC5WJgyLYD2djXxwG+KfwL1dGPr3JU/
9nvukoPZ0kVLkZp6zRNlS0eWwPlA0xBxWZ5Mbb/YTzvWqUd3hMgcIKAIRjnaj87wICEliqY1k6mj
BBIb7nnWaEXglpMj8Y4BhHZeuAFF5pvswFe0PeRaaPcvofKjV2ERHCKxEigRIduh2QPLHQMC1L2Q
tNncuj4NqLVh9jr5pnfUSzYYDz3UXlb6nev1gl9e0QO/qJLetN5BJXxUNagSp4Rrxbu7EYP6Y8T4
Yu1U19dQmXdQcmOdcVTaFLDjTAiOjF3TZxptY0yQZleHOMeyf6qL7x0jLDJ10C/KEY++U6UGC5Jd
sLt4+KcZO9FlpSfp6lvsC96XRGst1WKlpKPMZM5iQKymacv8kfn6igsMJbLyDO0GiZKWaqP9ecb2
huVJ7SMmM1g553ttNjz3OfTpIUQaRno4PK5nVPq73KXEX/rPTfulO9C5n2y3qPQjSanpR4jhJIwz
6lkjSl3s6POz+T3BW80NPC3g1bJLutdlqCQ5SJrexaxA/SwbxCym3Xq/wS0we2U4Tqv9fXFom1/S
dbanwpiRlrpGLjvCvAC0XeU9w2ecSLVGdWJw8OWYgBHgg9MMvgV4HAI8uGsDip+A+11+HI/m2iNi
IdNjzycL+Pg3GgAL7dAEG4nC5J8fvpuvq8PV/KgzNhUtUbMeJ4+yvIToZrIDthUEnIFJ9jZDjxO5
2k0t8kBuc5taOLgLlbMcrZJFgDXU6H9VdUuQcnmUH/5x1apXHHZ9ffk36sVuF/39ifFTdigFksHH
JKqz+ilIm6oYt1UmoTXkqZGdPlQJoqkdEo+SCTltN6fiLStJgeOGDfXon/EX72ujqv9Y4EUZ11n2
foT1Twc2oPS+8CTX8V96S4gwl80EK9dOuDj+txQgj6dSp+ha1ciPT7QCdiY0OIoesnS4RYuh8RzQ
FlJ3YvzsCoXOvQHgLvb/nYmW7LkK9NgIWp8XhLexmzOoH+2hbdaAdbFIza3nL6C3W3q6x7cmiM3W
jZ6mlEavMp51mILTRJw4owwRPl742Y7PiLTyoLKWPnvgHmeJY50lDYzqKiVh72n5igb6x3hrBACc
4icqcWAqKUaOyuiOQQGJ10Tzguedr/6MQ/cajj/JR/XbtRBDvVWscNEXwX5VRDLJma+J86aI5uXz
uwBL9QLrkjvQr8ywazyDEKh1qJMkP4KhGvnpnl1efvbAppHpoOc9vebO0eZ7Py7wCVaEtLALqQRY
QFsJaoY5vy2yDxBHax4cP4QdMXv51Ow6wGCECa6WmJCQlEJZhikLw+GdmiwyxgFi0gd/BZLFY3Ou
R8CCmWpZOJFbDmNm0uTidAo+jStpZ0TVwJaLcGzDpzNxnzfdiFCmHGEx0Uge/IOrLfDzsqp63ba2
fT/FUyTcRSBfBysRrqq5ekQstVed5PCWqjxTBLbGfrL35bR/MM3SFvL58k3FYaa0mWwYeb++h+P1
VBbmlhcOsnQYfhMmtGkO+48aepKN+914DOxss6epSinCiNeYqY3wTF/bDhWvYsElrfiRRMiCbuy7
MQnDcPRfH3cBXzAzAJCS5PPhkG2U/bZJSZLptV1qjmVxfJutVwwqC9ORAuAjAOkFwRbDB57pkAml
XnfrhZJBiLv8nQK+WYHgUFCMkIl75MmVu+hV7CM4eJgwBF6QR+8zo3C88BHw88gLh6QOBoc4x11g
QLsPdjcim8I1SCPAEX+sGL1zNeO2Dze1pTyeiSQrbdOvqt6TeijxnBxl4t9UQjrpErh5C8oHWARs
2+SjpG9tbL+6UgeJmerX7O1Am0wDOlCGK2QezSbYi0g9jY9RaU9gQEvFjIoXtHO/+yWVPNf8QRGA
T/q9PkXUTCHh+O9fNQzmHUtx3535LZqFBLLAlqtjuUFBUfNcuER0Acu46H37KM5XNTwQOZBP2Wdp
AMNeKXCgX+2fCwPX16yxb4N0HnwyizqJQJOleQEbhZ3GAaZIBYLOD86xTQGswrIc0LFxhIGuXAOJ
7cVlMnRLFIuyFHy0L0eopfBtx6+aLWSg2jujljt5q+7QittUPOGec6RN6hWm6GIEkeKDFkJTsjV3
38y2ccnkedPrtfPWXYTgDXRHpy9z1WVQvgLUj/WrcroCyzI+ujsRMtk6Vz4tGwff+Kxwl1IK69jF
T4OlzdrmYyOFVPu5KMenTAaCcwtwGi29Wf2Ba8DvcUhTm53OTRGWgNGFaQ0+P/uzBsXTUCiks/DI
j687oTVYs/aAFrBP9IaLdiDf48wNgUHAykK5tUX0E30GhHp4CsRfchUr7axRmnN8e0Yvo1rITuqa
8i/1R85Ow7y8UtnUyv1CtpRIuYh4HN1//bbMrxs8Ee0opCD/cZF294boctth5S0DUXrTg2W71R/m
X4absfpqK128xf/SfmRwp1Bl7jJHyRCs7vc8LSxEG9Uzh4KrNy8h/3vjwx5pYqcVJrfidacq1Wv8
2XiTR2f3OjXBaCrJT8gCeLMwA5D2oXN7RLSC/g97u9HAkeYqPPk4ZPeNWSawXUMi8yrMhNJ7DUjj
JKH8fWRxTumKHMV8UWV4ZNBPm+APJ5eg9aFWysF3nrS06PVoQcARf3OtC2969C8TlZstrfjkZFDr
6kk4lwxzjzwUREOCOtV4svdb3wmjFLkS6BI/n/HIN5t5PhifNhQFIn05/OcNocMxB5vggxE1O0Pl
NEpMqxRwzgB5ncsvfiNtckW1c1FK8S7gBDe2+l29ihxLW1iw/ZqsqxOWmj9VIwxKDsO4BNFjH+po
bgI2LR7oIWM2ItBuwyHUiQuDirTBlKdkdYMRmHHkVfWJ3Y8HvVqC/7M9dYdwJ0eiFXr2RgjzLp8T
dgK3Hr0PuMXV6cNozNmM+PHWqWFkvg8FeSRglHP8dwPuByOUGdxBCn2TQtsDJ0jZblbz0PwpfzqW
8j+fUVP37J0FfABxe0mm87PESCp9CpfmAmZ9hgj0LpzMZw55a6NhbRr9tWhtcCMFla1YJtQ5vkXb
m0uMZNBd46DnUsIvGX9CKLNNuhIvsJ1USlk2aTFmWPnPoQ2cEqoaTHsA1nxn6l0L1U/FU00AGu4c
Ez0AMRA717tlB9txMRg68PidS/9kJbt/thyTvan9HiePYZyZ7uokFNqUNSeMvNfplyWtp3U2vVd1
+vymNuOd8mZHkpZ3Ce2205EYHFUnMGaTHV79WoDsu4eXQa7RSAhehHAQHg7NdNtzTP7PJz3xolCU
mcq5LcpMdGykEpCyEBKRZA5u7zwhL1eUvmD2ZoOzL86jXNXGskVPUrhI1ZZPv4eGev8wjtLFFVSx
jKTHYkV2uITlgUEfbkHTLlt0xoxit41EbBgUjsF7yPNoL3RaFQe2vv7JeAsqKtUzgpZHY7UGcMrN
BeyEmOfeX8T4RYd5P8JUH/03gP6ZFLGKh2qFRLKMmItEZMrzsQMi358L4E9u7Uf4+Wm5/kJNCZlE
ahS7RMf+wUs4QcpOL7iKaXf22q12rwcE+Le1fjfgGlEkQBN5D71gHzYuurSxY6elFKcLY76mrL61
hU6sGjN+m7TPovdVIiZF6SX6A8s9JLppw1hZpUSq8QOu5GcHZTvIuIsHe9lxXIMqEYjGU0QZNDBt
JZaELowfQsM36hRnCc1G9eayWBKqMa8mTByPfy6esJBm3r24TcfrAHMlN9OWh7IovocXOSs7wJpd
SYUPcnSFUFHogNG8VhgFfeNjXQttxpN1QCAb8s/yiWWUiiMLXh0xWydBsRDCTOHG0BNbNlXb3+g+
m5t6brun+XEP/qwtDNQb2SBQgO5+D39/M1Fv8xvJaNW88Vk0k3fIeZyVikCjS5QHBbgIlxNIC62t
BioQIL8xi4BHRBzBgqbLcsGb7jySaFGJ3bQyMX4v1vdSIhKLgGfxwz5WeDWvdTctPBNuhNcxeHFt
RM6YwuGFcmZavzcd/9u3GgXCuCOjsHo5PpF5wszsC9O7q2OWGadEzHCabu52CLgvIWkxh56eTECx
rZBLnEcZfUlBmFbXECY0chjiBNMwop0AvgoqrK2xvlAa80EDZ9aNSaCvSAOGb8ATGLG8fAiN4z5/
GoxFyhzwzuKYJCcAPYfbrJgmfZ0f5Y/YvpfNxHZwztOm81xl0fQT6ZQ/fseCFikq3zOIqFz9fdZl
UpxqcWmEih8hsm6GDRJQa8fptqyH7Bg3ZLg9bfUVWxy6ek66DeWeirCIogkdzfvOywP6kw4LZMPN
ivf9fr4On8a5557bEZ3uNjlLibqOixm9BNbFx81fWSDUiLICHMc9TeDszUXxI2AWh4t686y6JNIX
yt58nQs2PqFA1IZnzsJXMHB5UWR242m3co2YbEDIOyg5j6DsF4R+lgA617GRfEyIqzG3fx2EkKLq
w8dCvE/Rnic7fGJefGnwwXCHXIJd/4e1kzPcGGr/7L/DLVio/f68pLU8XdaGqzQzikNvzEUhe93J
fxK3UKV8CQTmOsxNKGmDR7XLSrnnQ0cidJaiw/24kRrz7zd3uTVq88M+z3TgvSRVGPezGqNh2x+w
LBX/hgvgeDfLg0ec0NC524onkTW5PilncmeR3ZL2HoyGErOJ6nxkUprXDCUe2ZX2OS6RiYaK09TT
bsGNzN6UC9tZfT04VLHNdqEyty5Kd4U+9xWUEqiDBm73sK29z2JbKEJpE2dOHqZAZy6RTJsrOWj+
nrAHODqYvIse7m8To2AbggR+FOUsA8vvVuHswoS5gTDR49wzsJ2Zl8K36p+rjw+3SLv02cszWUBv
DY6RBUhbUHQGI9EBUW2UpaeTqmTuF3vgdL36CVh0ECXSTuoX3oXhZS1grwI9wqPF3AJiYWQzpgsY
vNlySil+vkiPvKVR02MGFaagXDOxKCdseHK/QfNuNDb8UzBhocvTQyWRT0430wdjtkfKGOr7WEha
s4zmZMghKPqy5/BWN4fmYENaUcNm+f6pS9MU01vG6YJi6MkMeQmB+KXj4ypAq61BbXh6zurtY37Z
dzWDaBe+1UvZkPzEtlp2vP8J5RONIJuIyamdi/8wuQbfViuqHBqocxa7c3V01aYrqxGPvhpd3lKe
kvMoG6lhgEM24qbRn5gOh1JOuDgbjUByXakZr8g//herYehS/DWLLs4J41A/HB782Th3nAL21mhx
5lXZqEDppV8+W81tylNGrYwZXgUx0M0nsEndKQS4zzwIyx3xxjQnhBu4sg8PkVTU0lbNHP7qSyrw
CN/phj/uBMg6bnzfTz28ce3gbE/id+J3TlpowB4rtHvIv6TFTbctaTtX3uSh56UAOIzQYRGtpW3O
BMgWaX41uKps5MJXMWtWFOJN4f4IJhP7IyyvqUWvhlrLeHyIj8rznQdL5uxS5JC/NaBL8MeG14sQ
a/P0H5pWzK3Avmu7JDnd41AC1TmubvmCwSbrq5ZUBbuWE87SSldbg6a5jpPLfXnT4lM0xBmjkyUf
uo2wLQXqIoK50gqQ97ah4y5WZIcyCY2TZ8s5MuaFhIod9S8nbdqsuD2zkhWGbYKU+OXfQHChzPEq
a6oai+OFWgGkz/5FL2D9/DkJBrycIBSEaz3OqZIFAgwX9edmydq40Sxy0HCfUUBw2XC+vb+fZE5T
MUq6CU9Bl1UaLuSQuN6Zr54W/fzTqOJnG9YgjvWGz43kcGuz4QtZ2N4GLah/2lDbm5+napKyCShp
YgylNKY2BuIVhIsLvD418Yc6XiGgEjXHQ132GU26BnvdS+w09XVqMNSvMwTSw3TkEDCI7R7gGsJe
BFB7NDAV2RxjyY7HQwEuuwRxAJxNC+v0B7h0Cfs8U0fMYeKO+kIBbWOpEpbPT3QVNPEqtm+rDNFH
FFMeTB4KAO6DggEh+PfnBNmD65MoWmhoAhWuwaPYMz10QHLqRneXU+QPBd31U2dfCHKyLzDifIDF
nEk+BSikLS5GPKuxRi3mAmWdI6fxhsBfOKPCGvlxlOOUTqWoV+24T7Q+xgl5XCdgJizlPdAuHdV6
0cXn1I9ZrvYJZjckV2glKLgGD776O5cI2/NfNZ8/ziTe9SPUPekxMSwagd3OKfkKg9awft2tK3xj
Z7he+BmJeE6NxMSSuW3PpWo3wUL4Nb8pgZUV0O4fwQz1pVTfWB0dpouJsbUjERykD4B5p3wvBf9t
WGcfMNWVd32H03zn/KoaSgxpfUrmdZugAqG35WYiX2H8UIunH2a10Va71hzNq3PGMDrOP09jXWBg
RaF11yE6E9dty4aYbaTdKommJRKkhxR6U0tmQCPrZ1A0qfY35naOVp6cFapuCQZd5I5TsiNGaO5Y
LIkYuIKxGl8cYTZxy0k10avULphAtcJ0pfj+eiMRqC5VowWVHEjtM4x9ieXgBuiiohluz5ueAzmd
0/B7XFuvGct2tNfu4Jhr3AnxeESGaEijaZdhwk4lS1RtV7ZEeevmPun28CwSDnAp1BPUR1CIrAb/
s9QwxfPULj6dzWdjR/5y0H5HEfnpoqbABvPGI7z0aj1zdlhca7SO7ELTEPPG8htcx2c1F1oGjn6x
b42fk9sROGJZIC8JZz5ZUIX94743Q5tcB8T0WhEJ7P9svKP3AinL5n+akyTYD5RykiauE7f+cnGE
gqB6VpQz1gCM6bws4i1hoKYxzqqXewTSC6MW3gBKzjMMleOS9sIHpEszmbASNzCC7Y3tZ3lAD1uC
nMRu6uaJLrmfvNYghMLk7AuANdJo3Zo2ZcSlsPfMYGOSfxSo1c83AjbS/cIMy3jMAgEt0KLkyR3j
GRezMP8TQHtmegeHZuPMh5+kbvIbpE+x7z4J3HzPpvcIEDE3EsTec738lTuF1ol+1WjkE0A7R83U
JTOwYFb3Ccf64PdKSLNJxRzcsUduVKWNi2HGPx61ysPU2XPBgqZlcWfYJvD084Y8Lq1pItAwt1SO
MRTR8y3rqJiXFYGVmd4wFxBon4o66NJryMPpF6t6u6zbo7oMgkYyAh9NMsOIeiiBWeyPyM0mAYwB
xFF3+YVITki6kNEbDLHkjEuY0yvdgue+asjwPBFj0Ppwq6XLR1kBDn+n8AZ9Rh1C/UxAHPeelarB
bvDGwfdKSLsIi73jWkhWhV9PN7qgRHeihQZxYzUoOlPH2AMpiHf1yY44t1aQWUbj0GvrcLQt9oNw
wxCWusZ2jLFUDYfupgj4rZA/xUXMif+P4KKyvcC1lX+CLnZN8bB14fin0hjiVcRN00ZRxQxl+NAB
/hMznknLgAJcoPCxj3zWXqXPSWwuFweuCHdUUGWmUt9+qYpXcpapKopE7rRmTygrHn9EQ6vyCtCB
+GeaAy10Y3k6crBEHWpqVKRytxq9QMnvaPlbe0QhS7Gudjtn4wGvSDFZoFTEfW/DqloMoUVn/BID
P3OXtADWT3U2hSNeWm6NreYykD10fILn8D3v5VxH/bcjkA69hxH9NtEoinInRc5w6ao2in922Xr9
r2UPyHsG72NkIPyjjZHser8kwHiTwOdUCbCRRb0nD9bpFCICbwh9S9l+Nifmomtg7JWufYg1Ex82
23AcfKaMSt/vLSOPEgQvRtDdBkAC7q2loCKHnOyVSdoPXnoFXC/R6AD1c3R/B0f3TlDOAsld3awD
q2+wbrPdWU/qqvUhc6G/c1tpWIDuYjywhexucwinec0nZm0wEBMP4ooHKsAnkrQqspyhG311xU2y
lyD0k12DSCr/+bCALLUz7iGWyEMXWytbXLArQCP4YlsHQag1lBDm9yuQ/Y5VuRyqIEvRSjr+b02e
gsCXFFvV/KIHCn++sUOiv0BwoahmC09p7+MTroun1s17nDZFn7o6NNzVw7+oe3sZZpgAqGRe9u/g
9EuHDZHNhKYOSA9DpljJFe43fip1gOdmdyz3enb5RDygq1TsaH/FGiKgn65YUCoq57yDh8EdOYkI
zGhqSy50xy6WEXTdeHph+iNv+PiPJb3c/1Hh78e4D/x3viVMpXwDE3l3pg3hsVW8l6JFt98G7qr7
WCayBIgzlgsqK+n9PFmTx+16KogRBDA8t0lkfKipqSUb7V0oZOGt6tf/B2DOVYwKZvt2m/z1ggo4
e51K1/GmHoQMA4F808/X6RQ2winm6toUef4RcEKmqRzsxg4OvgkTZlswN8HB7p+xQSQu1Q2CME4+
8mAwFfjWAdxyzWci647iK/uurGjBSkCWn4yt3hWw0qlw/GnJSNv/0pGtHC2iNgUZkvhnKgphFacp
AV4Oy23H94xQq2r1B4/LS2xURbCZoCjbgjXtaXyraxYLfdHqahi7bSeMIdj8XffXx9FOcoh50K4R
1yRApwUQaSjPofyFwQ1LfZz7DJlEmN8acHoWcQ3Jl2NcMUhiWNM/gEWsXz/WwTN4r3FJ7nGeywde
H+8wQ7TOXwCj1hYTXtr7Ozae4YYnGvl/EnG3poIAB/be21Uc78X/wq5vQcItUO8/InXuNsRZCRwZ
apj59e52etAK1FcuigXHbsCDbvgWpcscAJcBP+4T21WDMDGXtxXVZJih8rxPvzVTf+rHAmVvwLbf
CwMuRFrphkJKnMnajEnKY1pz3WRR7zP94ggitrKqp9MycS7HTrTgwjl0lWUwxDhy7ec7KpnjrwsT
xzckorUuxew5qSW+lOwgxP3m7l9/+vv0y3MZvsWTEeTh7hW22YRLSeSbU+kVpeLiUmsSeHQFBm1i
Rm0KPpHXkIhXghFrTEtTalEzHH+2BxQ4M+W3Dc0lSOjO1/WAZSSjByo3tuN/yCOFJA0XZ/V79Z+T
rUN3YyRRt/cIslN2r7yNfkeWSOGgPzSp5V/4NWpi2rMazKgTrh+7m8UPGePLmWHc7EZq/a5+AJp9
BDd8NF9XyYGHqWDPPZObCn1yGs1NKNddjQICM3DhNOkHd1aHZdTSQaSIuVEh+A3NW1lm1DhpKlYL
1v+54FiqFJ1y2r3gcz2TYBLv/ReaSoXpCwMO180LgxTQvpczn9Fdp3Ppnm1ECHrTmGThjfoDItcL
+/cdaU8aZ+KslpWGgcwv9Yob6K6yWlbP2+yVqahvnBSibJq8IJPaZtTtX8H8TxPaYLL6ygjuUagJ
Px/g+Gk2RupWImJErseXA5Fj9pQSn78kqu1YeYegboLKdB8E0qK+h97d6auhmV6qVaiZMIYNYZNR
NXv4hSfOeUKyvMMmmgZqBCUZtwLz4dz/49zOz2ba7YumdREAdKfcUB58+JZ1MELyAAS9aI2U6Iop
rrB4Fjv4yDOfcmU++ya95rsNihC/e2FkG7Ufdd83HLVTD9QRDWLPm9KI2pfv7riedqJ9kvmcQvHR
GMeqQUFdo828sfKtjachz6AGYaL5uGsGiH+YfiGi4SrJLveuR7kQf1RFwLLuURC4b+j8KHM698H6
ePZDe3DWsjjrUYYofXm3XHbANzNDl6cB0ARMYrlJrpK+DcccCcWrtqdsnwB3zZQC3vr9hPY0sJd2
5oQhYioyyABdEq4HcoXm5HQ1fuoK6yx6jEirdnWExAGS85AkqKFkJiSWkPpzjJg7hUprV5mEorBi
kk6hSgBtcn7zuioIGZGTlMijMFhpV11+QqfDNO1XmpmRjMEjXRk83GdYcJH1GV0rd6X28PqjxcA5
P2lbr5WgD468SpW0u5qlR3Fi9rz6NcWzomthfiIlZIadePECLXRiKKjmHkPviD4mc9Ww/1VJFtee
GUwOWQcwvK1x3GZXhW+HaPmzFZ20k9IcX9qk9oYGHPxyLCz40WW0fUSOO53VFqkHeffCxqbXKe4N
8xrhLBweloU+1XjTZKnc1RF7NHCI/+Bdfau/k+BgbN0vQHkv999Rzs0UPGsBUHLu7julgMllvWnD
XIIqRB5O1PlJnNDH3ooUL0cbbzwUJFvsStB+CgrrTdLfmhF5t92JeG0ydMzSQ6lmtPopkGrSfnrf
piSXfB8d5T+g12pE+hF1aO0SIa7j7IveGwn4/4qrayYMq/CK5lzrV1hi7RjdAFiY5BT7dVemrdRs
aIs/JOKFhu9bqPsv+M4ZZiA+77SlehRo5Nb2qabX04XCiLLVBe1xbz1R3u3rHBMiRbGNdIaq4kP9
Q1AMuCAi0wdguW6I9+P2XfYP3pcuLX/5JVXtj4AHiTbf4YuKBhGhg937yfOSn5ey8Jvub/+zK17v
e9lby4rYv3hCGPlx+/5GdrfBjvCGOVf3NuJX5Ns3H1jWxtz6DQf+ah2SerUAXxXCXrhR/3YQl1k9
i/garV7/vPgJuswCqnIWccHTPlwuyrhNEN2t59fQbUiiMPXKK/AfeeiGNU3jrVC/3viLVChEILtz
j8EhM+I0xonyILhdrXXEDKMdRcSa8+uzGCSZmYRaqNFRFP3qnsGKQeq85e7XbW68qWcDl83A3LlI
JtpnsdEKRke03Y5yR5u2m4bY4zw8iBxLbgFglnupj+gO3VV4mNCTlmh65v+HK/Tk4mm2HaEWWRCM
dsAvxBOyaVmGqCgl8BRE4FECv6tpdJzd56H2sJIDfPHVAFDB0LpK4IQO0sm11915Tvfooh9N7zuz
hTgbSqX7u4DRJJn/PxLYt7ArqvdaWKiO4xneSjJ8JznsTdoSyyoHP6+6pbrhU1SNx5yZxSMDByzG
nw0NM2FJ8YgT/mv9vu1R8maQxZRr758jDfwwJZGL4tPm38uD5SZfYvUZsaZmgP4hDLrhBdjpTCd9
tMi2M61SiMg1POnKxtSBFFzavxsagCnz08Guq7agfblMitruMPPVJ1IMkHcudKNBhRNG38F7FYb7
7gkj8C1vwH0RkIw7GDRw/NrefGeuCuRY62vFYPW8PkZ3QlDOGPvmBLCz6SwkUAf6yqxQZCDmjuUD
8ZRFLtNEMIt8pNwCvdVe1hq6lJC6WS0HGwkP0OkSp9BQzhp9PtdJytDJ+v34pil3g6oeL/GrUkww
XOKIyKzotl55EALyXoaR9MqDlqNafOynUx2TSVH9qFNk9WskqfxKJEuQvOzsACaMHo61WnPr4sku
iwki+ldPSbNcOq/dDw2eHVcpeemirewoa3aRKFIFggALYbPA4ay7CxpbYj8oqEspzO3+Ml0RMO/y
4OOryZWZJuDH+ck2gZOEltU4UyTFy7tm8q8TLmDm2Re70b2EVhaxbd043mUup9O8xuH7q6wDlBYs
GAjzmL/pVmlkGjCfP5ttjxRtHHhcOybNwNxIuHtZ9CSY6CyeIk1bQhIHlHwQFcDfNmKWHuf8vxbU
h5cS2sixjl4aNix5LGV5sxBQ8BkwIQpoVINadLlRcaPC0FBnPQOJM4Gtm6jDchcPA7rdMUx+acyN
PA+OY0ubKytSl9m3gmx5xAZ95wqtTjSZJnxW6sQm+E6xA4qO1sH4VkrQY/tdbaPRWXT4qtMUtcOg
YJk2y0q7baNFhTLkpMx4HFNkTVedBhnvCNeeiLv33RCDaazmTM66isCPBTDBaYg1iF1E0uM3outS
vBOI5euoyRxY2C6ot66rrwtuhUOLa4InYHNySMJcbvAB9FlKQo1PS5u6dQKsyFssF1BzChbbxT+y
sBop8CbsI/YlpdaA0MPwiEDgSihKksqwGd3RmgcnJ/pSGaY/HLY7sMN3IjJrbUkhNZXKZPhpp61W
AqUFyE++H+X0/KwOCjZv988PxfnVh0v068kD7e0F+WpIUrMJXdMe7dWpfW9lBQfMXkyucdvzBrUV
7WbKxzKFWW6xoZBluOwhQj1iFFMqazd31PxWML5bS7u/uHnDtf6HTy/6P6WV3JifjkhOpHPm441h
Yg2keQIXHg7bILckqvo9VLYgKTJfuNu2QP20TwYxTfg44zhDQKSWZ1pp1CyEmaAyEj5+AMtT6HhQ
dxah1gVaKb4Bph0bpQElQ/TfCQWWJEe08FMd1KS/L1wtdiCd76G2EpEf9AYJg8pFTg1aIITtLONe
zpUL2J1YgapxfeGYpkgbAWCUz6VFqoSVdYYJATbXyGYFkHVdnFyVwEJTAdiKa9ik2+D1AYqTpT5z
kbvnRYGl61ls9YtMMFM3MQF91bgdPHxocZnOsFRv86bldrFevg9DO1IP8qfw9jyqsd1NLCWn5DRQ
4YSd923UPZCeprCtZBNsiN2/75bZ3kI1gbTQs3D12J+NitfBbxGdCc6NlBoSoTfELbrFLLG1qioM
PDRd2/fDlwLrOAksPgCaS4waAShVMVGg1PAkp5kGH9kDXpFg75ptONxg02b45ECQ7DnA1/DmwZ4W
NcyXj07MeiBcIPylHiDmcHOJH0w34NOabDEmNZcfQercsJHC15iSSDCK6/DZa97aZnttZa5Dz9j0
bzCU8l4y+0gFjCIcaCSDvl9/BSgddytw/ZXZ82ivjHp1KURiOfnhN91izdZs+E4AaHhncDG2OoND
rmvPZVXdRJsbLFZknmbTy4W59lXHv5RXS65e+0utJo9J4RmDpaMAPzEI9ElCi738OYB6mQRAbQSA
9K3GtaKYQWbgoQt1cVOjcViK/KEMq0v5L0IRwZZ9BAUMKzOd5hbPi+vkTFnCyMHHHmsy32IJYlOJ
uMyCalUYbwVjjdO1z9laoK7dWxtxIEBbXhWGdKVPW0hhEyz+c2QeVCSeRih155G1m2NxIVZfF/fF
+k2GbpUForczunqwzTOoZN3/X7BLth9TpmkVHPdQ8/q+fKvbq1dW5/i1/NhwSWRQS7imwJkYKl7q
DfQ+CHBKpp0/jU6+U107lxKuSL+gcMMxpWwDDPFDH/c1aDeZwMguddV6XQAt+OZq3beAL8AlTS5r
FdRGbyGWTXvmTN1FpmJiCPB1/fgs/TGybsmkn4dsyJLn5EU+/YYU8aosmRfs68asBThYrB3zrls7
NYdWGbSjGSMxfekuHCS3sdJQa7AocHarlZjKwcbb38Ol+kZGhOYE1nxjQ+D3heqwR/62k/55qby3
kfzpxgsdU7nRF9rNfTiqD66lwkSushsPKjUeXrTKbjr4k4rSZFMAgMkmMZofhGbMSF5VrqC+oYrY
xxQGi3K4SYIWmp3SkK0AlVCKck6HxpsfLYbI6D8+y69OVOgrVTdm/DVyilfOdYqfaQMlts8KpmN0
AzthWrQrQV52JPt2B3Y/lLXCEQIZdFnPk9H81z/774Ix7aMhJtUMGa4AZzfs3zZzD9J0wQBzBmHk
o/TUvRq5QzUdxPGITXev2amT4UDv7JyZzxunm4JQRkrLBfcVqff9rTCQHrpxnOaJoqfUZWu6fL/b
RmR8FiFYa4MwzI7ST0bAgzYBrvJJO/AExi6COei101LRHTJcMo5wRvlA7PEL+YFSV5CSVvfwBj2H
wmX3IcxTJN1qSEcq5Ai+97J6Q3VJ3XswRNiLYCUPGNrPVAYl/RW9DcpvahFg+e9gpocBrBGUgsPb
24nDh8UfPQ3hldfoMoJWiCH5WrkrqlrwpAs+Kkze/X3VFiCjqirhaQlK4r4WpIAgqQznAdj8UJyi
rKre8m4FmVed6wfSsKrfJDN7usIW+g1GUwCDe+VKlZ2l1GrLQTay1lcByI11rUR5ebfRIGPY7IZD
0ydMMpD5rQq7OUr0EwhuWKVSaxFFTvZ78Dq2UO+ToxFTiCObT4Q5hNQJdAsaxKFabtEPMxWCiU2t
cuf0sq0r66BT3fZ6NZnn3G1xYrjcIhbeoizBgA2oM2PX24qD+aiQyLzldSWY0LAcAEsvEVSAAD+q
+GqLxtFA6zPa5FmwPnIxSr5wFX9kHDGI9c2rTxZd8XKeUxHofY856y0jrg442Xa0C5h/vjJC5ESv
laaBan0fzV7LyxybELkgNgzxysQgXc3XdCZ9Wt6Syfmk9EnuGg9G+Ms1S34R8P3+CRCvkw0SZP/Q
2nXmFk0hyIARBECa6qP5QBo7r03jV1J6n/XICO3XYAEBgjzIH7MiIiCTPfeaMVSKtKBrAd5Iej9j
iiLe+JxAEgIEjJXhyoj2kvADedMYYidshTBB1bRDltTcS90TPwoABGiUhsl8/HToCloePJDCu1O9
ggGDBLt8YDcJYYnZ0kvmmhKrcwW7cQmeFbvY1juamDV2GwTTCKHwPHFz76ULa4IMswABwNaHKBxq
8sUq7wA66yx3qaQX7GRrrZvq4yS9xUS9at7v/FDhLoD4VrSvwcWWLtXPFkYHLZlaqQ6856PFRkhr
pVYhSdPEvJ+eGg2bba8AjxdI8MJm1AKpcHJwn1MOb8DNksXQ0np6jKg8kNNjZ1z5NhOjOg+RfWxZ
CNKjfkc9RyxsJi+DqlvBXa0HTm/2vygwGesrxcvN0VTpzjTTXzzO7sCQhtrp1lcmbkbYauwgJUgd
+QKCuTYXwR3LIddSs/grhSMQfWIwo6BkiB+kkZlPlVizZyWV7Unxj+87uiDWm4c+/aW8rSTSsi42
VRZnX8a8mLet6yzEFKN6uyV4OIs6aaupOnavP2v1YVYF3cz0Y3mXC/Gn0Rji3vsGDugH760I7MKG
zrfJ05RaDqeWEqF7kF+KWnZpVJ8tC/bHIa9P5KnToTJNK4X5iPWj/ePL8oUE9zobD2Sljzd+0uhN
U4X5tVeT1ubZfvC1C3Gld3DA3md8WSWzlyGHkQYr9M/ZWLUnyhR+nbw1CyOfx1JplXZcEo1g9PxS
5s3GpJ4hJwqrNSOHKI27QLqdYCcKfIlYsfqjHBMXlrrNIXLCYAJpVINJjeqDKwJf179OfyesaJl3
WdVPko1N4Av/1W3SvGxtrWWITCKBpclYRe7ddNPdjTkkob0zVDcIHqu2qGWAtlyCsSRNKT4kQO2t
zMaOSz9EaVJIUJqkmNzOOsZlPM0zGpA3XIATBVe77BfF3SoEKzKh2Ipd+qk3JpEuUC3QBoOFRJXj
3kdrdYht6vjhYyjlYLNgx8nOuMdfqbACulUwF+/ztm0XNfjPCfJSQ2ThHRTd0W7F+auLcww2NW6b
MkAZCtRSjLz1PxIRiIwJX0LbJODPcBwQYKd85Hxjh50tS4f85x/2inAwUTQB6MvewIJBcAohj6fu
IlYE9BZFUqcqKdYJ/0H3J66GO6jbLUBoZ/1BypKk76UJT3TJI0GdPeyuH33n+vTPUFwRevVtyXag
3mAYuHUarMuLu1C1MAz5iZ9to63diflfzePBLP4szjPm19d2/dQ3OHCYcRTVNfZ722kBqjjdPO7a
8SVzYdfkavFau9e7xcmZ8NtswGHbUHyJC7ZVtlRz02Z+SgreqIdDMPTOYyalbRGnjZRUC9Rfl1Sy
A6dQpS+QTWlIpKGtJUEqA6v75Dl8PtG3F/TMWEUbwjYb6KopdbnSxrgmBfLaXdA7XrPOH+NsXcaA
N3e8VysaHgMYBuqQYQ4nrzsBcLl3sIM7iDiQu7oZQtgDhsaDQ4RV6lnbifupZ/XdNTmSKp5x5V4k
g4y9gC2SjJzi9EBCL8S1HnUCPNijnq9I/TZJbsV8/riWuvBs52+gG+gaMOcnRj6CaKIMcO+QD1Eb
nifTuisPLLBZjP979gLGNhUBa3jgqwsyAyFK2tRUprZR29zq/yqRqIdbBSa/I1ukXIb34/TjnKLG
dDApkAmAi2COXMa60lIS7+vP+fQaF62IrM42K/pTuB5HwOOBNSRmtiTnkxllb9Ub413Enft+AZjp
f5zU+p4KWeoT1VoUhanwRW5WmzXMsyuMyddSzxUvNZjUmQcWpdphuWmQUSGxc+4BdnRn9kY+2C+T
H1U+yD9Mef/pLHsVATQO2dN0RxFrg09hAJ60FhRB0rfOtNCG3c1hXgVzbt9h0KDd0wQz8hFAOVl+
xPSf24/+Rdri1wHF05B7iAYcV5998AIctkWN+pNGA7BvkxLCovGp1Ja1W134uxqnSKAakXswUIyN
FZgjji6QMKHp0svp1FDk4G4qWEWBCTIYjcYHY+uzOI0ehAm21LlDEE837u3BD5Mqfe7mr+X/hdXD
hFA/O/W+HD4EvjKnbFXAlmp704+5ndDgIoGUZedaqNI0+88X2aDde5JyHtUfNzSKQ6Cscqe0QK9a
03mLFQ+bhPlYOI7cJbEwG38QLLSPa+d8ZdhnYxfQHU53vZ/u1NpuaZ7OKo+neEMa57pIut8dLLgS
wOBZDNmaJN87AH9kPLx+1Y6A/1KRG55LZ6Lii6prBGsuqA+wY4CYwhzw8Nx6BRJKRJCIOQ7TdDpf
E5mKVY8s7q124y+JhMj0lgnwLGMtRXP2E0DYp0/Jb5KdU9MjGYFMe8712Xn+we6vChsm6q7gp0QI
5ceBeq54bhj9Dj3ZmiKWxdLAfLBqMnJz5V2P90JeIvtl5Bpu4/YnifUTVYeidh2i0hwGmCPe7HZh
suK4gvN9c8V5fdEuZ6vm9Wk982OEaSdeEjnUME/av6/RVfyrhFjHVIS62nGNzM3uvXs8z0ZdERJ2
JCmzaYV3gbqyg3YFDj86B4kQylx/OaNcEe3Vk3K8J5kXpGjFHZgpC+G8nV/kOMS5TZ95g1Ywepo3
ZBL33hpt1Ky5cm2DIleapHay5SANnLWtoX65TawEPNITYSX0HPABF12wkLSjHUH6WfLfhJ+FhyUW
aiEihLEzSElDd1vZBkQRK1YaDHzLVlVbZ398Qxxh1Gd6d5c42qDqktlh6tLieURx/airxPScwsqK
i7CswcsBih9TW4j6UTNsj8Ko62yXpp0kkvC/tyhz1ru8u2pjqeuSHDCWukZs6OqjDBP775kn0zBW
lLfhraqoyTjCytCV/4Tq1oHOns7kTwKs+mn7q/Qg4AwqXcVtS1IWbPhoBHAiGCs4TvZWage0MFLg
GGQ2i5BZ/WeDXPexrhfFDFTV4eJioLdrGPwmE8DHWnvJ9ASEJMCg8WQ1iyQeZqD9Ff4/cG0GuA9s
Lcj4DItTqYtj3u184TMRjt1P7WQ1JxmsSlwNMthG3Mj1DbZ9fHg+ialCI55HfFPXb2TSqdo+edsN
xvr3t/+EScKW7uyVohM4ExzGMDoVdXBn7I3z0/yaIpT0goMJPza+CEZe3TZhAy76OrKMgBlQTlhh
Bo/b2+lxBP68dYmqaM1PpnWoFPOvBDLOu6sybx5Dn+JPDT4k/2bLoQzpSV1x5paVDQzAvwU50hH5
ahFcDx4H0EmJJhpvb4QoYLE0rXe/0Nj+g0f+pNo2A3gzRfvEnFcfNktQlJJz01S4nDvYT4uggxhp
rMsD1jkFd50VXa+wECUbdnHUMQcXhRH0lHdsH8DTcnBZxsVGgF5biy9viDOQuVxQh97cvnhFcDXG
hnDRWC3je0rly8uV7YJv9zSKWr9XDXQhVN3pQGF30HKe+eefM/z5Anx0RsrQzhxQ32KxgBFCeuJu
ffc0Y6cKMqHpjLiGX1e2Rk48nL6r0pdZ+E79Esm8K+k30brIxGSlGMQiw0mxrH6VZNtbu5+eEO9g
Bn5WCHj85LMz/QoBJ9VZtfjKkdWkQZ7v+bg2WnHWhfJBQg0WqRc3/r0KK/wpG3nE6HUzFrqOXYev
B7yeDAE45v3wxePOpg338r+fvGch9CGlnG5uUdX74aD2qW5rU8OuwCIAzO9nH82YHgyoeRhddiCG
hsp3BBUBd8XKUXt+0NWa2S+E8uS2sAQ1oNbQDc47dHLD3xpcgh+Zv4KHUtx1aj5LhLifU7kjMfDg
sjT9lzp+wlFdfG0WBC1kYT04+kiC591nHlyVVmCNrQIZB6h6JiYrNJ3hgHjNXANb9+UJNyM+E/Lu
NMaRf6WoXjpLKms6ad4pujkUe8AZR2TB+t4+CTbIDo40QXrftEzgo1GlsFxYWLJLqvkzn12wi0B6
RanlTyQXV5j49mfXNu5+upCI1ejmoCckk06VAHWkfK4pHKZVMhMfL0eoQh9O81RiGxKF629lsWsg
jMzGWy+qOCd54ZWA+WSUiFWsk35dff6sSActzeyfwRdwrmsoNcJtDAGannMPeC4UrhTBVEi53rGZ
mvBlh+Wlm5pmLHscqOjbnDgQ8IaUqy/49vQPg10kaahq5H5GkceU/14PX3lbJLWFc40+knuHHiJi
ochw9u7vTSjKGvFCpngWZArKRplRsnQFwxOxTlGfiO4emrwzzM+pApb2Z/rJWuGv7Yh+X2+tZgeF
BS1A+WudwQC/EdKTn454pKN2EK1LjhQZpPIza+R/5Q1uGZxAe1ENu/FvSp7pBUkptnxd1Ngy2xVA
e7n++mroLYpIHDomNpvRkoh7jZlwI7ETize2CAxg+C4bIk09FylI1amXENRUyPTNgl/xzOUwGf80
CZj1jT0Pd7JSr2R8h0aAZKqzY4eoWBk4dSjmcfsRWE260HI3wFYOAzE2uIR9qbCyyBR0Bfs0lL3M
Ohlvm0yIuHmXT2dGn6Tjom8u4A3cHRg+b/crwc92prcYYmECplSo9xB/evGF2ftr4bPexCU6D/TF
d5OItzNDtuH/szg37Gwqt4WbjDcnou6nWMu+0WHEFqnSTqk45Dwa9mCYhqOylJ2r0MFa6DL4imNJ
dChLQniEbCXdovP/zTXLtXN6Ta+uQYkIrUTWP8R7RPv1CHQVQKbJepwnTy5sfp3VavzBHhKRqPAS
xbFg6YcX5Zu+CyZuH7nUnZGmfVCg/xUZ5CYP0kA0WyE8u4ToDEDSMhmUQBtSdCQWOvdIpletWXpC
xtvOEh0HUyoYG9Zjmow/cM9bnKdrbxQB+KXszs0mymyYMTJaGykxzvuNh5NQ8w5i2iTRh1aArrcZ
9OKOtGUTsl2bqW7TjS7odyPIThdKp5XbeES/f0c19oDPlUgfzcfrwNrGOgR1N4tmu2BY11WY+lZP
N8lpAUr2SC6C/DQRx6uZ9r1bSDjdI9UrwMxR0hYnH0IoSJon1iKFG53BQyYbfRHnVbxjyXanF0Nc
2L2cil0j0Oh5+2NsnsHGu8VI4gixK9DJpGmPOpY+g561oM/FRZQbyw6GCf3z1EyyyvygqgBYREdc
d9h4XhRDAGE8sU+IDiAG3z6GYX/m26xkxGa7nq1CgSp2Eh/bvBJB35EvldtfnC4K7YeOwHswDDMh
CHSg59Yhm24b8MPk6ZWX8263DpLEgSQESztP4Ou8FV+1L0CQqKL0zil/MDpRwD3gLvSjE07ardKq
hHFptFiyZz6JJS1xPEcYjC7qnccQugnlIt2GBhGTlP/bzOoQJgaMQMsSJ2v69MOCVZ5HiqQI92ZD
NFc24gvvg4fUyeNAv4w1DFr0iOc6SJn1gRGMRlzzgPMPfR1UB/Cl44NoxWRV4LKiV2BZVlgakRFy
uvXJtMNvQ1NQYrFD6EKajjprJg8BBlhZ1qrpxMZoViEx6BF2o9PJ+G34vSjHo4z2s0B7cmseulHO
UZJhDZHpOH7uZKoT1CxNCL9ftXDWAsv/ULa6t3EPi6EHo1arw3regtyskwpfdiHhSlws+1LSQrDr
WLtjW1cbHayBd5+uv/IrJ9ojuHkzhjNOFkgMZccIoRgPrWZdgngfF/44uFdISc6IzirSXzrmFxaN
7H4u1nOe2oUJAm2IlSuWY0W7rzf4YaiSubbLzHpdBRdZXqU2bIhqmj1fnHkM07j61m1aRwZuskXs
B/dEk+Z64+LWtnDvH5fTPDPGpq05pCVxSebplySmu/pyhhzFKJdqi+XFafHKUxI+R2TZFvySQgcX
G5165jk/ZRE3YJhnCnaDrHb54cfd5x+zNYcD4jhkfjSXqM4/7kTitXS9gm7VbGyDnpj+uALqyLDR
KnmacmKZQULCN602LVV67RoWM15KCttFYv0fXywEOuzApdxgzNJsdxBHUpHv9zD8mOar2+47bFED
MU2y8fd4uThb5WceXMl1CW9mSlKwqBUBUf98p7cx95w4irgTf1hJzspSOy8WDHtX1E1oun06iM5r
0Hj5d8XWXOTSwSooMub7+azArj963yDpIvgNBGXZKvWGyU7sNTaZvrowHbiIJxZvsRyvMqYNH3lz
FWWLOVeabOF1oryAvzVeqs3/QrNnS5CyeYMHOsJi94Jb972S+ZqKY9t/c3KgJL1qU9gv3qVeVTlb
GC6yXeqeITrfJcfe9mTcHgvBYjS/iXUcgO18Gjxw4Tw+57kS/72dKoNd5tbaU4epB5dkx1hR6DSp
/mK7i8YHxHn1klfe59gFmTZy4mf+Bi4kcRvTDZcxX+Lu/l+HZT8yRUqwW23lOitcGYUz4M2NkF5H
hUfYmgbTCQJ50SPq2Aa9YO8rzgAubYEmVNAbifsWMPk+jCY0VtgqR1axkqJxUmempZNZRpOg9FRo
2fjAKPRmnQu7uVLpzFkmlrlyZm6bI8NIXyeaiVN4SFlOJCRE8Ycr6qvvDU6HYGROyz6G7F25sVEJ
3EL+1Lk98q0JK+GxPrHAz/D843syGkL+9sTliXDW9ECUT/cZ50ObMhLxEH8w4cfQ0d6NUB3wDEfv
xDgDxADs4eRs2caxAYvUOL6nypj1G/gaAsK0RqXys1cdjVim83sHjxnT82AbzZVAafRQ4GqjvDLQ
X3+7xjrcjdmlEHx1S49hCUa6TS1G8tEyqY8Pk0Yp6yTFPCs8XE9z5x0dyqN6jwhNYkRXdbT8Ytbo
mC4AfmDYP4roANRxl+Dwu3EFjkUjW6t5bkv9dZSlVEOAsW0OhdiQRCLUkx31gejxnVO3sgFxkftU
rP9lpVVXLNlU2jfxokmgzgByXnJMunMLz4s1saF7NfgZq2tkint5oN+VK424U3ZCShUVR17fynHw
SXNiOHv7XpFVGhdLGttKK/E4E/W8wSB8wXHzLpReZHXUO3rMkwopEuzgk98qxjpon4KA7T1CsATQ
EJftCQl+ArbpqlCAJ6Xd3BD7XCbWrIo4Wibdyr768MppbxnHwS0z0bhAYrgxvQTo0uOpgrWIshFz
r1t5v9jwsUrS4zPg5nt9gS3zGkZxrmjlCHx1DMFXgT0s8SAnijtZLq45xRgFzMH1R9+9O2PD4YmU
rIPCIslzeRMVN7yAFMNBw5q5Js6omHgp6toPAQPs1MCAXMMkcYCrAZIZuA0XeaYbhzLLn8rkrOv6
PPsSC65+T01qnEp3zUzy0cXnYOruhGSKAx/HUzVw+Y2HdHppUzP4a67v7YPii4CQmFGOB+wpgP4G
pJxOBS5Xb908jEftqLosVOCZSM8oIEaaF0SKaunI824/Iq9J6eL36j6lv3I9DexCoS2kkmWBI/7O
0h2HuiJ3d0hkv/72pgtxpdKxooaAwomloHgJ0DO3UnvERGAm+lhRze1PbeUv0mE/o9p9HY6IWvUH
EfBYp89OxcyS2GVL5Af6G+XfoxR7JO56fKphovjaagJPI8TuuI2xib3ODBBuB2oAy27PR0hbXY6j
1Jquv1rIaEra5+9qVipVLg3fubM2nuXDWR0q0ncJqYnSWYcPJwIilGwZr0MDgbGSCbFubKEKyObE
rqijPUE4AXMbVbhOcnMqIcDdkBp/lu3sz/VYZDC3v0vvxPVqs8+GHcKhLRnDfVxjwPsBPY3bBBjD
MwnMsq9mVyjZzTwUU/8REAqULybzV0F+oPtkswm4zG4VlskREUtEhs4UStlx3t8aKCifUi/U8G2J
MUu6cSGLjRIWaJ2byQ+L2Hlloa8I7bmq7cevtKFbuBaeMzRtVo73ZKo5RO7lHAAjjvIjRYxk90+X
PSwbyZzfdUx0Rr7bWTQmWTAAc1h8ytj2UABcap2uMAekqKFuqiEZrwbBjYs+ck7YFRiV3DVHUzQo
jJCV+oPYGBuCpJbxtMZhvDb2wmeU+CxDBr4c/WOzxmCmNiXYPr5s0uchhzDARyWdl738ua+9fkUh
bc/PQehAPhpM6+QbmZexhwsBoVBmOcKnKWQQ3BAXp4K7dslz6LEG+oP7pelc+EOj8l3/CLVohDhe
Rbb9pSUkEOyUp3fAFDc3pc/oLdDe1Eza3zj3oVlzsC6NJ9H1V2WLxFlKt/Ftl9OwAXmdxnXGxiiA
hOKcvntcehm2Y5vImZi7r0ZnLqVA87XPSHlSyVznbA93EsW3zMtcbbVq7MjZNYh7N9X95+s9fPL7
th6cOXXX0MU2bKdnDbGOXqLbiQMSHR2sCg8BJrh+2wahNxcL33Z046pAl2r9pu+puL5pibk/xGZ3
uhjexJabRerYUhGwnCXLFwg8RltnIZCtNzcjjxaOvGu+T413yPvQPJSmKNgc9AzUBfPWGhymlH7m
fCJy+RdKCyoZK3EJVVQu+MRF4QyBCU22vBVyUo9R3jUIn3CvpL3piDM/emWITgZq2ZYmuqCgKfui
rt6TxvFEbEsyMRvd9f/R2MGw4rqkv36Gz3lrl4tSKyNO52Ke+XImNvd1Nei+8aCwI4MD70yKbchq
S6+dj59BzL2HDlXTJEzwmeZdUrlj1CxBLnxjoKeB9MKmaxICLVpocarsHSwXQA7m2FEX6rp8K/t0
inGbEAp70Py99o3H+tRdb/G3LX5S4Q2VYBzWKKlGuR+SGhSkqtm8bLfunupwEZQEAh6JHuaw9Un9
SxPPw4Zc6OFTnmoKlMn1cXAACapYzXgEgj2BWf+iuYuIZRsSE0IW5Gft03qCfJhPyO4krVRUdDqJ
Zo4s98tjBVJ/SfIbJ3RZ0dIKlN3uNXGBywpfZ1lf74U8n23BFE7yh5H0gVS5x2aYOMmdGZCi3No8
W9GnikvqDskoWPzLPOWUV+/TK7wTpTjNLWoMZWXtBEHSTxWlAvUEDJD9uzIENo4Q6GUlOTbiyXwa
F6r8wLDTOJ4PrnW+eoXxDvww7/MDEmekgU2/V3gZXux+S/W+n9mk3hQwBVrqxg/EWnU0YPpz+MW0
1WQNEOTDnmYvazk/UasDS8J05QUoEWezLgSzWBnbs8aEqoAGGeWZNQ5xJXQeadYSW5KJmD9yF6aG
hkIq4CIrlP0/zOINoIGo1sH1BAspFFNhbyEQfvIpPdyXNWUZfSBwuDK4CXnxkoX6SosrTvQTWTyV
bPMkkLGjwb13C9+FFLdg1R2c6G93XXTWtqynjnGq5zXu//c6pEBP9ABDztd5jwKmlEg4Xay4GxV6
oC9R8ybBrkk5JM9ZL4QC9lFIU4ZxCE4tBh9uC9lDyrgGURVfNCKXq2MYXz8sVYvbdfewovHfB163
FO0YvqrOCC0UR6aUt2ikIxXAvNricSfu3vy+Y27XnnC8bzv6kcZOusyuc821D47M3Y7XzVO30U3z
8166hu70NvWVx+zC1j3OVZQPlwSvPU3QA24YOEYc3KCVgPgPKYR1zcr/E0SFWcQAjQe3E/YW2vEn
2Imt4XBD8ivYzwoo/QIta0uX0wdwNwtF98GiTUI3p0CodgqfkZgUJ5fDtU8MwZqaKV6HaHbvUX6H
YyJkoCtJFCzvpIE+WzEcwZ7CurvhJdwlpIMTm/HfQkDoAkBxuzzX6Udi8tJQ7OQwGeoft15nt0Tu
fdEPj9mAo8UYeKplA5YREJwxeTKIZUYe5gkHmXJE8Li0ixzjHYrLeMoUQVlH8I3C+RLlrT/0pAGd
B1tkRZTh4zttw442SF7J6oQamk8VAnKxB+42BKeizQA6NRwK4oMsxvrID2vbPUAhn+1XzDUmojv+
pMrQ+D/ZGu7N92XxcIuLfVlvxPDw+hAWl06camjMoAn0ezZRMl9xMdXf7KxasRoGENAAlb2sEC9R
fgduA0xF51Ibq+gmvE5dvhTShqwr+ExjwaTc5rf19ClL1CPaDBtLG8n9mHM4zupWAUY3GU4qG7f7
4Gr5TnntGiTvqVTT2mHMjCX6q163DnnJ8iwsssWTepYHXGDtorPFiGQUjb4i4rt1NdS98vV8PcMW
r1VSeXF8nPbLjEK8JooFP5xSDtOxI28gSznui8hjDb9Pgg0xLLb0PcIpo6bqsJ1kujqy2/mmbVgX
PnPuR02817764nCymxi8gImvvUl/zM7N7OYmEUNhiFSCoMMbN27UFiSh2g7HswjfBgWTuGaCeSWn
y8Qlx0LsJPdBAQ4tckfQ/lN442304LdQl9WR58JqeL526zXVBH0uMDamx0tFOg0rUPF/9oifZ9fF
FLlOqX1UjV3R+3LGNC1agf4ZPN118HSdSf2PWQqm1otk2foTmi3sFA4OZH4fQ3qmFyNS4xaobFaR
JmT85xS7u0+/eGHLhUmqjcXwl9XtNJKfC8ItSEwXzKipbwuZcnNz0eOdOtQGdN6r/MGujrnAeYBK
9jZlEHdE3iYrIgvbz/nUmvq9XR0T8rfUROOgCUvsw0HhKNjOnZ93iFcvf8OFsxkoi6gimaeSAIQZ
h0kd/W/RVniXlKhpbXR7GwGjmRJITnpRxGvvbYI+uBkuBS40n9HFu66Lx94ubAq+fJVMPqfOWKSe
47GHXmimJjejfW8E4WCTfuQQXGPA6AvUJHN7TkF2GzrMQRVfL/roAQxHkAB7LgWOwIxZjuj4/Nr/
KUpeF59biWPBEh3WLtMsaLBKd+xTu1Ia7aMP9sUwpR7tLEcF67nTYsYnnGTbKUH0CPILncL1Yvco
Bmjy87kWZTXsY5UJ+Pev2FAONQV8m+uKXlFYy41rAVJWMBOjxEoXOQ1zoICpa2wRAh/YbkQazDYk
nsVQkiRtS31Bsp5RpJOK4itqaKrFQQLZv4JCxL4AbA8uUqBt0uDhQAnaHLiu1McPmHq+hrkx1aoG
TYlI0pk80bDuTD/ZGWsVHhPNaHyW5O+BoHv2lCRkWWw03UaObtVTJBNa1JsM8hyTJNdwQUrDOr13
qIttpzbeWxU680FJNnkKq2g2EbHTSpHrhI1GXO2FXPS0OcH1mcA33UBGYRFcaQHvynEadf8Bq14K
8iIka9Jx1dxYEjySrWdsA2IlINTLv26zLHvPkjfPz9nh1CEFpIACgXvqWkX1fOlUHh0oNJeE3t/C
DEUEafN95Rss6itcgNFmNSDo4P5Q+fg4yj1mvWpF+gjT/VoC0MlTecFjVRVknyCnjWRH0XKKLFQv
6Nk8kquJEao9HoUONUmY/c0Rn0mOSmudUwho8Dyab2GuRSoakOGHUpNqjHkLdR23q3eHZhrQFV9v
CQNGv6ZFrfeUenyysZQV+wKuIt/GFmA6NHi53eqovU4PAxcFe7lAUtqjzGpL6Xjz9B9KpE/OgDjI
vMwPZyaGeyOXc+sme525VaetKherB+AYm0XE5zaktwGpEkavKBenNKTVi5XMH9GbZalvbGz+bYK4
YlsoO9uJ2oFtE1/w7vr8R5KkTziRqqlRpH/kTHfac3LbzUrYVuPaAOcjfZ68JEFzs8aMuCh4M4iL
RdSiPC3eLWwkdGrZ8nfnKp21ObvB3vgesTPHjxSHHU5HdJoSeu8bUYYeJA/Wq8Itu+TXuR3TlQbt
OHMoFzF3qxzDbQtCVN9huq5/T2Gj2RFtTefMB+WREKBGPXSSBFSphKU4mlMKC8pDlM7iWArQagVW
0jIXDJHQv2qsv0bXkPxQIoyCG1aeEH4tDfjCFvm55qMydNbXJ5KV8unxOnukA9mDvRv8ihbw5b0N
8RrQBmZ1UHA8vqPoKiLnIJyX2NIg/y7rxkwoBXWg5IOKCxh+LCvD53bbVL/BY8kdfTgVXjfbVS0y
UMMndPGXHMQ9BadK7RwN/kQRzSklgT77UvGEit9ez9AN9VZJD41yemyTH2TAyszywmxXjblXLt7P
LOeNWqgl1PMdr9gPmUlJXHqN7SGAp6IJudxhy3y4aXUMf4e7rV81wTtgF8UZrl5yg33pDIQ9qPRT
8UNSBlLAqChf7+0sSYJluEimSR1mdYdJkNWkDOkI6EWgyihk/EjdRnyIDNXvn1XbWMZ7hLQZJEM4
BZ17rkt4RHqppYDqkj78D0B09iXlrCPDPdCAlk66vnIjNLA3RNhAyi8LDiNA3m6LbHynwAcE4Q1B
QPQSqMv4hvUIKyxT9SPsyu4Wy4TThQICHWbgPJ/H1gaqB0bBirMhbYu5fiB55e87nclcmUsrpe9a
j+yYNaV+uA7c2gkqsE3YyIZyrFT8cxn0CnyTN+urybIZvHiqXl6f0fanOxxwKV8LwL/EIvPRJ1gt
x59ZUs0mdLaSsHrhNVYapSZgA/4IY0fZEv2fvft9xfBAFfpez09oUE+zTaG2cr8uNQ6IBGd4TFPN
ssd0c4Vgv8VnKPqACaZWVedm/PptcVoylLPW80jM8iwhfWHOv1ZB3d3lE6yC92Im8gy1HY6HCkDT
WXjDc7iKvNlJpdolLBZPXONjKHGeCSLdvpHh4kooxei+BjbC+ZUecyignwzt0T6hCUUqYlXOyyKz
3XZVXjmTvQgZ5zM3lC7JHx7X9fv24zk5zlK4/ybWSEumngU7/AszCwBIBQmgNCotiK3RgPJFk/dP
IrhH4RjBO0767X/NoHL9dIMJ+WehMEwYi6fvOpsNcVvw6BWhJThpDX7At9C7hlw9Bm1UxzaPdnSS
hEj5t1efe8WOAJvK6wVK3+1CMksHCxgtDYGEYMeCbkkk3jutPnQBpiYS8XGBVjlDAQlf8eF2dcgX
w7sLLKA3sYGl4rEBKBM3RdIwETHHYI1NTDgZ7cSv1aLICITidDyi/hVvVcOpTJa6Tn6ZvgsnJIV0
IYYoB3f1GwzoPGxlmkBmw4jekCl06YQ3w4EImLesb7cPydED53lVjfMUqAKoQEncW5yk/rQluvuy
tblDI5XQIfge6zzQnmJeqOatiPiShm1cZU5iIKhHyC3xxOzvKoOzhuH0Bw16Via2MbEbuDx0gEwm
82uG1HAhF5jU72scf4vk7K29HSt0ZLCh4VYm6t39JOs+8r+0g2eP7zODKDTzkybARIxCcggLUcHN
DximpdfUz3rWxkdbmLKD8fTgrSmAr6Q55ndYUNWU/7XpuE8JCKJuMfHLNeNaarZKjsOYmHM2AyU8
R/qBmVHKwRHVodYDbBNuHvb86a2/5A+mwysO0Onn/eDnkJp1vNDMdmQUWRmlXGoM8eCUpsBkBAEy
I9sKW8VK8bCeEXxioWkAnnjhuLkpgSVObNlFRzmaffDt2x7yeygOMR0LTbtQ3Wt0qhdBb2KczrD3
scm1OGigviy3mhhIHxKdjcxawG9o+StOE17TK10wWEl/dCyNzz8pxLwndlAel7InanH9VmB2v0c6
B0QXOEoUoPsnWVn0lQXpuqvekzhboeLabBV3v/t/myvpeYb7Nt3RFWDA6FiHqKjZy0LZcUPJp72w
fQfh1PxGoIptG9bMMrbeIlcnlavcDjd5PCsUi11i9mDzA3w7zkBOOejPt195KGi21gH53Lkpv082
R+nLkRyhl9fakJwKHh0aPGUF6bKgrbfuQtwVYCWa1AqiKcq3ciaAParYyyIempixhmMcsI4j2uJS
HKVGFiXXh3SVfC9eSIYmVUPqgdhFdAD0loeBCs1jsuUKCOsHNnIVULxfqHIR0vwS0NoLnFK09M4Y
21CMgPwyAfE4rpPEIBZfz1rE9BszuflON9lowTXZTfyKyD9P9mfZxvrqhwctbrG22VZiraEQV1rV
oAWG0MtNGjaKxivRcY857d4qGQfbvSm6WVIcnwEnBgzUAvkCUZrqe+JpEdfsmddUBojUHIqxOUl4
ASsF3UjQ8VsNC2xHjw+1I1Idegf8CS4guTFTbaU6cLkpWLaE6fLXpd+E2MVa+W4AWt1LzdrhVmaa
ObVVlPrAyOW/j5+4iQszC9AphVVE4ep+/b7z/2KzCyHOJ9j9YGtImPyBjxqP+yKUXVFFmOZmgYU6
mJgKh3miayP8TCQBEk4LjrgcSHGOZPVfGAqCHeyKWttcgPa3jVFKrj0NShKcCgKBgK+eWnxk5VsK
uWOf9zpvmD6jbUNcFEpK/zqFWp8+z67DPXgMV2VD4ya2opa17ZknREqPZEdr5ZCiKEzUGuvTcRTb
FQDr/93CQQRaQKI821r6q52C5D1bXfnnZ35uTEYQBoug0lTRfqoR5gMNTHyXCBIqZ7qEow/wH+pk
+G4Ywr93NjZjz5B4tpg0XQT0HcWeoaNVRSATh+gFFtdCTZi0gwZfjJVBYp7mFDPlIAmCBiyVJe8S
ZZk0krcBJQdOSP+krPR5zN5kF3KFe3Kp0VkqZK1p8q/K1nVlUguiiansF3SR3waQ9MtETAjGLGHY
Jw7/YiPLKoMof2pRKG4wkEcCsZNze86Lss0VTk0+pUfbJUPn3awXEXDN9PFA3PqyxwY/MTMU1XpV
8fVpCYTiJ/GlABKOPPnCQOGLMX6CVKRPi6B0lQI38JbNEAGoAMFf4PXBgmpLDZYlo0pajgVGHkfj
mfH7tH9HrX/lmg3uFD6qcbxZQGImLWjbxbp12CauAdBeOiAXDzdwS0jS+Dkl9wJNKfsXXZZJsWVv
Jd9U2SyLcadT/mJ+QSxXamZ9+llt9dfO8qM5pmf6EfQeOwxeDDLk4QwPrKExPUgx76PnE7nhlcUh
vFjMroJVxCh045uPenqdzEfagUdA7dMHFwk4bgP7B+myxlZEMrdVgXyKmpl8f5yEJLdKphSFylUr
zh+quO5prI9sYsA3qA/o/AXdPPu4RPLQOBT2NC8pFIFdiuFhS4vRnIfzmjBCtdnIcmjFuaFmY/fw
rlyiDkE066CpeZ2/hfXAlB09xO5AAYE2EuzqNISu87RyU3ZiHcp7DdDNOFiF/O5TVtAb9QuPQL5d
Ht94Zyswwos6xjPLfh0Lxt0kZU20cN50Rl8EMUMSQ+dXU/0pXwUhWhIK4IsT6hC7YXxWYayApr/5
CFszLFP9RvwXZwYnHFa+RfV60VyBkwjOmapeyxpf8Hw/ncI4/PhRETSvNW2rWIMJZrIPL/I4jIBj
P9km+xilPl75IC2xxmjYdyNpx1sFMwREG94+DGM35s5c1B1tTN3OCGftB9z1KgmP7kN23q8BDHeh
6IS4XaV8G/jActgJLxD+9p8bBPfN9O1Eucb87sNQdZpQE2IfqDXOpZXMCpIImFkAg91/NNwpqpaM
MdY8jovGNre9+UsS21WLrU/jrArGAvc2Wm41GfE9Lxlqo0tuxxBP993CLu7grttKic4zoOY3CWZM
ydK7epFWnQdrJickg4RC2gfJ26oTXL9A5EDmgQTTIeS+NTHkHXbMqrXa+cLXt2Yl2YQipIHcuds0
k93uyLKcD2hhc5YgBFYYs3bDeqH0oQd/eg/mrYAtfxn+jkUU9KxV13MJfcPLtpJCVU3rfKR+lynT
J2hwskcXzzoXTcEBo6cMG3OlFDuxlaP42Srj+pbSqSvJweV+e9nVKAZLMeGXOQO/1kB3IK5JfsvJ
QAfUWltTzCW8Etu4cDP37pkYjfFRZYKLRmDiAeO5Zlmo5wMaC8TDzkPyhTiu0rpB/b8RejnDVjJc
tfDIVLoqCulPJd0h5dvdFNrmyylA6g8wb8GCUrE4jlkn19wVn0gZeiUAsycZbLg2Dy9/msuyZJsa
Mes1YPWUXQYDExjus6kSntun+3UmIFYXS/rI3QOE8sh0CIIuSIyzyubxx0Jt0ihmm6wmdmyqe3NB
fZ8XbvhX27PFlYYZTRTfgRLKO8FM3rT4Qs4GvOP5qoqZNHFLmLSKTUZmb33GE4n+6NXOXj4+XR+R
SaVYNqjCb9RgFGutG9DEMj6CU+FlXIPtXqAU/PWaClEWODQU7pkaUDnc74hqV53uSRwNqlY0D85B
ln/g5z8tr/2Pzr1jeUgDZDfBLvHPPRIb/AcDVdvZXPi9lS/zW7Pw+smoBsqccasIBN4EOSaF3zDy
mDpng54Acnh1nmMUXG+VRlToqIls3fJa2nz/+uFNsyZnvrMcXjrCpFMTZ8IpN64ibnRY1dwAIEMP
5kaMjFUSD0TgUVFqwp5LWP+rMA73vOAXbJTz5X7e/Li4Rx/M1UEbKTU6+ZqXcPcoS73HMaqpBagV
ZJQtqKARH8Gtfa+SyfhGS6Q5Rogn77LRCnNTMAY2HjfVJDeYvvNePVe98mTc+vTpHKu2U55yhsTF
43RtT5TY5ZzN3pi7R4J/SLu1JCIfim7bod2JcSle99J1UX0WU30qIyOu3VEA0TzIiZ43ydjQhw21
NL+6qO3+CUZgQuuqxPnlPU8HI6FdTLZQwkdyTxI0JMmHA+y2Ae2TG+g3+USldcK7tjzWLULR07bf
sYge+kCfIXzL7WVM8nmnhbE15bmJ0Kb7Ly3nKanmxfARq74ymRYuksEBo/yQ4T3AyauR6S3ESLau
RqzgvGWD1WLfaQfX/WJYcu1eCu/Y1uf01LFIyigjECz9Sis5n/tI5zR/XXI/pVDdv3u/3EdaaCTa
8XLuYfLII55oqWIgcAMVLxCpRgSAhDCo1HKl1BoOAZbEdmDgk6YDILTuotSQs8x4cSQkpOjHGtAX
UfzUtoK81RXY+88L0IkcGQseDZicsWd4Y4FWXlgdaI+IYYsVbeOM+VrPfSziNalZTu2iqnUGt4zI
txzTUxg7itJiX4SH/xb2eWpomgbQOfKD8HKWnI7KiE2CKMN/8wrH3YrLViL6XTROol5APrTxotJ4
CBa7JaFCnjGJ9v12Bs1Ygbza2xnPlRw+mK5vBSjnMN8Kfg20DbmHQBWWMe0SY0jwsnOx5u2cGCo1
GtAHDY9OkwUL0fUoNDYwiKyK+jmOmeVt3Hv+h6wcZGGKXFy5fJQAdk4k+1GwuW8UNDxKrgRgRion
qNIqDAi932mPlR8SdX2PVEObEVWfMmLDxvgAe9NcL3lfrjatrJYTMKIAumBsjWrz9atdX5bhAD+7
bJgjcTMFUj/JZ3+d26Ra80kg6rOvcnaSbfdZUYHkTLq+rAxWPBroTvoFR/WWqM/bHrRe1WkHBMHZ
kC6kOiRTmWg3NQeBJ5JDTzDY4vxgOzho/qrZLGSbZS9wcaCidUxQKKpmvyx+w+bNy1WzqYTk7Rwt
J/FpHesO0726z3DJBl+iP8P1bLzvvvFZliBBXVuRp/kHyO0FlEh+41AX0Wu4luNDEjXZ3VXg1Mmb
oBUR/102tdNf9LIvJHPm2jC+1yl6S2qNcSpkaYp5a7yNPWes8opdcLxYFFnIYzZ+kyw12XFxv+JI
E8ZIKqLeNTri6hYcLdTstzz6Ih4ZFDmm7nKXS8+EufUvj4zgXgUjTIOWppIsHk1bmY860iqV05qU
fgg6AjBkJiIfGse9tP3ZFACTBYKllST5twAFgQrx2Laj2eGQBr6eYaeH2PkTfMloOJNEHChIy+bP
EwPQu328YDTfrT3noONMBDj50FJ3+GidZkvGwTaAG4TbiBaOUOSh6sL3HGn6zTnrTULAroYtSWXv
qAfU9MauTfU1N1tznYp1VDN65HQlo+ifOpFla6PGGcJMh4eLB29QfT1UJN0ulgk+rvDa1sCw1D6h
K13Amci1kywSKwq3bcNHjg1k1ownnvIEJENRwouZVCDIwdt2gvTq3xtGwWY2VrCEF4ek5RbsH0rC
ZZCf4u6lDK/DynCrFEBV/Y9tqKZlCjU8wKFMUYxLcXp3asrU5vzPsP+fHpObQBZv+Qlkaj37PhxQ
TsX/NwhPjUGDyMAuXhHQEFE19PbHSKlokAyHtg0I3Jg0ppVh8s3bOjdZCNvkXrrlJBGAXQQVi0YK
EVNfxF6+PAUKqadyvSN4X4xFUINNA4WYvje09unviIhrYVphKH0FtPJQtUZ5kfTPsdRsXZ82+lqR
hmP64B8BSwS142LBoaDcRsp38m1Gz8iwWc/g1h/xXgYdTKhvF7nSbFRw1nrF2MmZluE12Mp2jw6R
TT5MsKnbQ9qj01R5pGkmaofussOuF/c+sgA6wjU+4yogKDIS0db7YlG0zgx+RFBtExgvvHzwduJz
NNb0TJqwS6NBZygoUBGJZ124st9MtZKXIu8Ms4hU8pQlj3XeXLvsugtIG/3ScxErDo2ymgeIC+TH
/WS0CIbrEtyJBpf2+GITLhsWowY4sgekauxy061sgKjiK+N8EbxF80wMHRI5CmkB70utTcigeHk2
zA/HkOFOMFEj2VLe8UjI41hWon3XEgYKw7ME5Yq/fR1tpDoNdKAxeSYlrDa37vTE8SzK1SU3Ba6L
mQdapQAsIEYKRiqaqFsGpzISebA5r198832vxhK7ZGQooRQZnMTCX+G+iT3QI1eKZJ1T8FGN/Viy
GcSfZYmsCLiu1yeGzz5fDOIK0Bbw0a0YsbqcibwZzebOyn/xogJrWklENdoc4pfJmcsGVHHo7fEv
eypK9dmwxOO5hyNgzdsp6CPiCgs7rZ4Sb/kRtbWDuuuEaSEWoHeFb+m2MWKGb++dRZo0ovkjNgVj
FdoRvPVwsJytpU3jEkiuXrjH+85qiCUXjgXjPFcQ9m6Bz1iVAJAm+/LosnSIrNyrfrUHsCKZaa4l
CevHl/PVy0irgbCeT0KQn1qI9118Aev76cvRcbvYcl9OSzRYhntKc5Z1+iEnQged3AVX1VuuVgQQ
RoQK60xP5drT+Rug6uX4NGY0r4XhSdqvh1nPTuk0/LmBwaQODFHsq3VxeB0X6du5M9Wo36xWlvxr
wAuW2cRP5LlTcIrnsVPan2TVsFwwaTW/LzVm3xsIik+wVCXOF0wkmZyEtjM2dYibkoACRtbP72AW
Hs+I+FL/jbur6wPg0GPVb+tHP8JMlqLUwLqVp5Btxu9VhhlHdlx1IE4fGPJxKA8wJZwfhxuxg2o0
BMpWGttzfYzSBGDD5z6mqpJvO4627F6npSjjFdWqbFhVWlD8p17DcFxeJTS8JehFiVSPh2EugETB
W9utE3Kn25mpELyeCXCF9GxkMUoskZG7U4mCOvetYH3g7YLmM8RdhYQsXSKbXAPnWI88Epk+DMrw
aX/3N6yWeabPYDd48K0WabaswQ4SZ4pNvCuFM9cwn4u8y+yKtlQ5CGeKbJlTKRgHrO0OQzArs+XE
4gpfM2/qcdGEJl9NuCfbVf7E9eDnXlMB1qjQE05xibOWCBWI6W+tn7IFKc0UCFMcFDE9YISQ5PuO
j2BLQ6UTSKTNhtB6RomOvdsxYFKa02GpW8XjqP3+nc6lI3qtUh5m8T2QIvWXlTMp93VXx/PfdOJ/
Yon/+MnWbWqOBauAwT2hNbAlJMfkV/HkGvvy7GHg1zk2I+36f0vNcIgdrGSCK4k7xtEqK3qZ9EW5
oUiWWJM11JyFWtkARaSNWmYzcoIrxxBR3Y8Y0S2iu1FIVbhJIh5CI9jbn7DIEH5qDTHyDu1HI3rB
W3vuKMvPXw0SumGiTFPm4rUPHj5Rww1z9ayYMZbPmec8sQa8tyb5R6iuLJhNTLQEgp/qtPG5greV
fio/d0fuz/HbcxAfO06pooJle3DE8DWGPgSkgb8KbyftBI/P3avE8o5VUMPJDfLBqxeS+mmUgrT6
JOwKLXVEQpx3dU3zDPw6QUSh3CiXt61QxWqw8aad/tise+tXW6rRllXqCKgnVX4gifQLirFB19BN
x+zL62P18JvtMBUlwL0QyiQADMrZkD/izu2sl99Rq7Orp5/r+PXj9WJDoITW6Xp3RhutuBC1JBEh
AgLCm2AGC4vV6DW9Wj3pkhQLJkyvm1aZAvcIfHrGHZs7ydKLlyWAiPg/Ol77hVYOYZoer01HOC7o
bA17ACN/EdfWnUw85pVe9ham1irqWckqckdsETFhEy8SKawZqFVUxlJRZmhx7GegRcyqh9P7VOaI
BUudZ1tKyiqmK3MmZtRabe6m+wLcmpiWmHYQ1zDlQYJt5Pw2ZxVCfRKa+UcZpL8qgkq1vs7aLY2T
voAoCYOZkU8sepzFCQalynrTTh1ZlQKW7StRvRqS4Fe4LNY5/0P75n6AHXXEiIBYnB7seS3CWCZo
C1Q9xbPS+ElwIgSz5ZE1bwPMpDDJS5npF/cz7O0PEUg0cd+0jUT+Q0FowYHPYl84KAjim0k8hBoD
pL7bBCkf719LawjgysidLTRvBY5PKgAgfyl8zg1K1ZE95ZgqgslADt0n5fCbhbgRiK9S8PnLP7xA
k4uf3ZFJIuAunrkQ2p2uHCt+hpSYdO9QaPHjz37oAQWiRFvLVpvrFakjO5UPzIPH14liSHi2ogKO
2GUkKGjmqRz54617WHVIeBiRhug/4aRUkwnx71AkqfJwUlPJ2l7vuLlwMZLm7H4auOKWS3QcORIq
PqkFxYcLkVYICmFnYVP9v2+BZzjPli+Xgwh0ro3+7pcEr44UBOKYPRCTfWxRkJ4LH9pugpv4WI8n
uegV0oOMdqFKZHpTMtlBib+cnJpO7THn/AaDvLYJBS1cNnq2Fu70Wkge3nEOnKVqCikk4pEetdfT
Al/buWzCq+nLG9oJ7Y03seC1CSDn5j6n8tT8feR8b+7ave2TIsKCBD0CVvuJlch7CrjuVW76n8uJ
HjoAWf9gyu1klbehPvMP0D31DxwZRgUnFcizUVsnY+ulal1cgNQn8bOy0vPKhIgFT7sYvmNYWRIW
cE0kKT205tyUptASXaZAGu/N0jq9ndZXynV5cyeVZps6jT4LzWnat6llwbxa2D6mDgTUIgAfGi8b
jMZF4m5WRuoCMVLwK30ZhW8e/6AFeTMNIGKXVt5ESwxYgDaLITdDKe437qU99uuEvRJGXpa7JJvy
v9RnS4knob6+GtDtUtzvLOXX2kBaET4bIacZtTT2dcisK+YG0qHmT7hsdd3EnErjBkpJdhu/VKlh
BlKKEhP7sDHZ2yz/yAeeJ0MWqZkoiyrkcWUS9fOpMIUUp08Ht8xDOUZx706gGtRJgBB6bvfal3ft
KGGAIT/QuNqNB8oV5Bux+1oryyaT3GNRx8jhzSjQfeb3SRq7Iqw67ZSTwuqAzweyiM63TjEy0Pg9
rEcbwyF7jZcSDB5/TF5v43yUzWGINV2Z2BTjlaC0O2OFcyoKj4UDz1/dpi/Lf+G8khCc8ul1bQO7
xb0Sg6X7x5M2N4zeNbqnBjrCRdntmDeFP7bzWpsG63DEG7orWOeU9lwbt2LUj8/RE9i7dUODbXat
xk2eQVWeE57VmouXB5eKUoS2hcPoc9Lb3I3SJjDx5jhdqgJvJ/dqOKfuvtNe4/K/QrTY290bbNul
gkU2jyhyOpmY+zYX2CHBKxEFYMzNkciPnME+Hhz9ddc9naDM2TlH7PO1aj3lBhF0Up28W6QoDc4e
OfgTrGl83clrUT+LCJbxzaAkS9C3ZuihWn4wQS3011w6/jnAG2tZvXHmtGr+IDX9TO5vqTMEvlli
BXw9v5d+N1xISMwnO9k2Kw/Wl6zQbn6ACTGxSuY6q3kRtmKBtc0eRcbNaHPG4vM8W2SRr7YjLRBI
Be3fSBfceIYJwv4POUdx+p8RPh/sq2IYALQNNuNjVb/+eQPSdBkV7x0EQoLwIKi2ZUmqNXA1CHpG
3Q1Zukid9rt4mcz/MKrs5/MXom5nIry8bvH4yEb6rcn2/pGkDIVeOyDvkR8MIzMW9GIEVGJGT4o6
hULBmTDGwwVYUBFxO1M5/N0Urc/Ry41LJe7aHjReMbHphal2hO8nNuq5WTShfMvW0+Qno5PK+3xc
gjo411TD+/J8wiuX1w81YEZXZjwoKtHnZhYj7PUa/SGlz7ni+2KxVT0YBwh1dIWoQ3luN8Io/SqF
rN9SjzjewjKu9gIO5gjY9LbCSa5TMydfpqvdQXSXsxR0Xpy/KFl9AofVWy3SFDV2MpQgV41jNju/
aDmpf/HJ/2NLO+mAA9HtZU7i4nbbx38aImKc/KEdDctpIRlh937ZJ2eNSBjk14vhMEsQHta83RYR
asWTAzpod+4vNd0hRXwnLZfDv4hrBX2MNUAzNvs7D9FVVClYAzpssI1/CJSzspOvb4meMQIWd3OQ
U5YBDwyI9cyRzQp8NMea9TjMRFZjmHRzmTvUhmcfR3hrGUhncrBFw8Pu8jhM+kR84/LUKdFPiq9G
Ip8keFtES465joru45rsa/6C2B/xR5tjQcNuTAVwnKdRebfcR7RZdOPkFNDxwjbmvcl96Gxasyvj
aEeVBpssUWP6kBNGZnS2LUXgXD02I6qu5nBbgKdkeEiY5O+8MdCPMly3BxgNOti3HP9zcTVlRPCx
QJh64qhxAljdpCq/IKbMHsybW/vhjHfGqRPYtmrAHkDfylxSXnr4YUtV3xPTSaHINtT+fZAddUek
R84AZ7LJ7XGdYMjXQ1Y8PDFy0QtYmXFiuW4IViPVx84LqlVS6q8kmCJpdYS6ixBFOMPPgzPYwlgB
auf9rc9eaPywN1k3OYynoPrlzdlVH+ja+QxV5bZJV+BQiDamvVjhJgP+027fOyaDGBkVezZjYrid
hUIJRgg4e5UiqgtfehrSolwdJcQFjgm1Q/KA4CZhzUZrEVdPHDpySHZ3Mi0kffgLg2nS3bOMq177
MkW9JtgfdFNIlKKh5mLCIzDqV0TDtRQLUrZUNUs+AnkNhzq8tVH8+B/jyUzgUeoNSnm6BtpXyTal
HCimoTBuEUdHxTWVfiYp3r55LNNqJTng7vUEKnXK61uox7kOg6svGIeOv+tE68PSxrnk3WHtww6z
cqURKPFy+oH1IxKQJAv9yfcDt1T8SJYiK3qGtsFPs+p6q/vmnSZyu7HhBLHYculjGDBIc9//G4vX
yheGUFzjMm2W/fDb52StH4Kkf27nwKrSCvp4NeVA/qc3p5CiMM38Sh0aY5sUL+R42DY+9F4rNeFP
JPP6KOtx9kXyvdoDqr5x5FURbB09vh3Ih7EaHZ1ua+7E/AR4RFYJ+1ZNCBGvRFu2CfCrcxpYvgye
pk0ZIdgMX/7DxCo5Q8VF5E5zdTIzjvYyiZ+0nqoC3XHjSp6xmB4GF3xewrTrOgCXwG0/RI9q/rFz
jwxefG9iicSEPmGU28HGCJEpWD51jIVOPWyEH8kneQx0aYPhQj4kBzVHoiu7xtX9D2vs8DVQJV2M
8YEFjqa1uyrBFAbIKUUkkipfoJ80v1faY9VwSSn2NlJtfYU+xUUA6J8GAGWbBVH2I640B3IlAhQA
gJHTL+W0Xg8E9K+BGF6kdJrqEYH86aepfJU8zCxr9SZ8W3AO9T6hOQrYF1Kg8LN8LixKAQRWLqFe
BoEkryqQso8Ekw3XfAEEeLeuVNUlt1CNyL7SHXnrtqwGTzHqNyWL7hC62gKkemaNDNwWod7BPeWt
LpOvqMo7x0Q2S0u+Hykx01LP6DVcLe58kYqejN1JMQ1r1Q94712JRFEsOKZY6RWU3myDPTDv5mt9
Q2cb9aFsmA1NUVDHehGYP+xjIHvwM+w+jBEYCGA3GD02Unkb38gkgLDYkfWRuCK4+ZjUEsGPZdUe
V3YDFB7l4Xx4f4J/HJkMpPOtr9pfXPHf524H39HSwNVSo66sE+Sw0AfzhBE3cRbhOHMSUxUzFfoH
K+vbw/TqGsuHcZaCUjrJw3Hi/RbGvjGqNyyW7HHv+DqgW5y0vx/f1gfIIo7tSy4Go5MawPzVZMJ3
smRr8l5Qpgb8Y4U9AC514Jy5Vl8xO4cwhEzN2SZ7kyCvb/2hPvAVDY6S0JIwFpYV5wXHjo+U6F5u
ixB+YKwDwm1XVMM8vdR2H3dtGOQaGIUQC30LyT9a/5Etp2pGTgXbRg3fPOHSZfGL4p9rtQAvDWzn
jZkYAe+L8nMrEAwZ9GH/tv1GB8yVmipSZovT/KHa+laAJ8Xf6bbLyE8UqlMJtRbCm712Je/uxBLn
2d00thTkdH3aO182/xvSYfmABl/ebNzRFI8sCc9JmpU3xVj7YffISKUr2okliwmconfi8t4v4QYf
+oJxKNahNNZ+0PRs3uuMNmciXqJMFFq3xcLPc0u486iwLI704k3Pxj0jkx93YJRwLDAMewWxCh/3
ajHuEH2xS95oUM+H7sa0KHkOY7XwP7Vpf434CaXhUP8mG3eYLA34jfqQiLkhQg3dL9hhNmhoN5Z9
Ig66HNHmfRwxR+YLClAiNOELVtVJEwr3t5OhdLSuqCbU8Tr48yoikjkXcCiSwiP2yoAUSxhGIHmr
QxjpUY3D/XZzO/yzNY5NP116HhL8NTzHx8S6mst6Jkfax2PCuPw4nmOrY5yjSW4xlXeeQI7+r6Yi
+zDxfWW49vV8MBYFKuW2XMjHB6rdc9ouUxJZXcMkTIvWpOMDidCaQDzma/CZgmqJXj1bGjk1WGVV
83QSOM5E3WNX2mZmQQ4V88SzQQyyA7c7HWNVaWUPJ8/GIbQrzre1fWw5nuvZERTse4FcBlclUN/q
FXuMJSpnadl4fr6jPHHsFNGBpd8pL+rOuEBlyHdf7rCtFeNDyICV25+IYXq4j+ue4+BlOWEMHAMG
4lcEOE1M4ooxufh/vwjh4JM3tRzpP6ItyhXUM26YGMCeBjQ31yr9Vjc5/WHxNzmJ9wc/8NFr55ZJ
RgWgFlCWiv2hiTKV8fSTST8yyzm1Ms7qmPoqCdGq3nh0WGepkZlOTEXKx2Zi1xZEYDcEWWi02MRb
YIRyFizFIr+fQXdRbYFTL/NPUDH90lKK5S4OGCtXr5/+PBX3TLQlpbZNgXz6VkbFKdhHtpODE2Nu
Vs79L+IEkSpjW9bzmp35mfZbUx0ROebGsX9j4KueFuk7kzhOBZAIEDy9LaXuadyqUFkxcobHWIKa
ASkvhSIymbHsAL1zaYX/zdAZReYSQFUtj4LI3CjxelHgUv+3XenLWFTY3i82hj8TkngVf8eTJp26
YV1MseozsMj/MiQ9kkon8QRgnqmIAibj8dzXSvVHpIkXbok3AApL1tk2DoVs4ltOm6OWspPAyJEJ
C65bGiA58la2w3woX5yn7qplQIcypPQN5xZbKLLP6NsdYMt4b+Bq5ACGx+++HxnS4Cjs3CfSf1Ah
/gn064XBkCxyreBUiPbzfjfpRXWQ6ZIr4FTjwUxNKenJt7W1EBgVk2GDQK03Xz44Y8QFYc9thudw
R3flSkLW9LzChFFzVqJUV28O6d9coBo1WdQn37OUedQetrFT6r7XiF8nL1iL0f0RRSmYW4rpemQl
Cphn74A56OLrikAorhKi0v4ER04iJFdDqjSWu6fHQnE8/U/xaYZrUJQkiIr3UrDXclhPUbIFRhoi
WlPLZzppzom3k++jRGhmysFDKUH8HuNkbrSu9E8wAw2MlyNUeUaV0ic4j4Al8pG+RWPee4vwrwnz
fq87ehwSr/NH2GWpIwPmS+iRwvBXYKphTX9/05vmc9lAdQzZ5Fr2oYuQj9I5zmYAU5aMCgCbkrGY
mQ5fvkASWwQzT96lepVyL2LNI4gT9EtXp645RY9tHarRJRtIG9Q0Otdis+sEIZRYeUgYFJNefBNe
Lm1AoTzb+N9xcWWej7ZKG+O50pzJxrpQgB4YY2wbI3nt54HStPK9zw5TRtlfvzG2ry5SXlYeikWR
0MGxxNqvQZf9Jydrw+R0AAtCB3abUhu9mX6WKMtaztaNsc+fC/cOsXwxQAAag8aYVbGF978GXo26
e/5/0NlDDdH09Pz+juWU9nRU4uHwbdoIBL/xjeSzPMmBlTiUURd8i9qa8ZukTlHfIpgXm+xdAyYm
iwPrvvl9JGoOK9N+YxxD6T270uL0tkTzVX2FfQPV0KNACpMj6MbxZD/TGgIvLVfNoD7DqlMbfn4T
4bAaHhGsSlEIY/+a4Oqx/haqeQnusOzP5afYhQxIzADktd9/auV3FLKrZd4cEf8YxkHU5pQ2sx/X
tLlTlGgEpwjXFFLYqIsHEeEy0hT4exsQJGcM6nDCs4tU6dIrytR5gQBrxq+WHGSQBeQZUBretobe
miUHEZdFCpUVLV3fUs8hul+izTEIJOYWGbjAOibyUlZFJSfgQZeCnWblGI7/Py++MmIQbD8Teypv
cRn/bCYi2jWjlnXYYlBiRls8oZjlr5mosBlqvRHJYKUPIe9jhLm0Otyv7gCSYm3GT/PKdtkmaZwK
YrWVW0gSIr5miDxkqq0htXPt0oCZIjlN+asr0+EwJz1NNMh8ilPN//TqXrRNFiosUFcqwLWBUlwg
9doMn9dYYVqF5yc1ZK6asE0y2xMbIN8WpwG1VVAKP3uJjd5O1m/ngBTmXs3PpF1TQUIzTv/h/DWv
dZIPMUYTcS6DUldKks2HtSGu30JMLJagjsCx79R6FW24Rr44JAoQd/k2cLPq5FX47EPIgVL6Ew2Z
LTEBVpkqhgj/1Lp+to971MIiGYHEciNGJHxShz8vpyL9O7CAlzDXy6lE/uemGntFVZWwIU2ILAqn
oXiBiFyH1tEFWQw3nE3IDq5/M1BGf53AAodebV0SkrNI3nAjHcnaItqdoztc0ZHPFpdE/WTPVU5T
RlGZjo8MXmqvYQ7tZW8KeaxTG5qIsgi2l4n/eFgmtP/IImYfNarB3HytixzhdVjbmYE4H12ygaia
5KDh8+CvfMriFsK55IFzJbPFbEwYHnzuBEH/0E97jLjFQNkf8MzgLcGdb98O7HcDmO4qrzIT+hQ5
aw78sJOi7PpwSJIJw4ErAbUtvptlUDIMkd0pUS+cqui5rnE6yQtYru4VDml5jRLPDGpm14hF596t
MKhmA/04vJ1vWOLurRA5F/4z3PhFCg5AGl6oeCNDTf3DG5wD/d0Veru8itZOgzFfCBK2FwjSUZsr
jQ7NSLrO1OT5KH3xgJV5fen83Bx6s695jAKhVQog2AS9LSZYF5WsFKr1fLaE5KFJtolhSgeWUyje
iAfagPjcO5k1MrBMM1ABCrrZUkM+FxcYkTJH7zY6hwKzjZoGouKF498EnYRLQLFThh3WF5OuIOBZ
GYWeZkJLM1VIkG6uys+yD7a9gV2hyuvdhhbg2byAtize5Jjm8lUIWqEY44cGExk+z4JB5lkVjfzy
N6StL4G3kqvbJo9dXgpJDKzoRLm6rkDoHmKozhH1Yyy71FEmTzFO2Nw7r3DG1cpTxLPKTrUe/OT9
HPYXBaaln0M9cINEEERGYP1we+8AjGXT/wo0y1ia8FnrDygUyiUF7U1UUf3ldecnEFLoNS2tpMVa
pyU9Ixxq6fR59VXx6E1JgydGEsRhxOFPBEo7RGaeLHvaAQwfxEOornjvaZx7hCPSUEJ0Iu3rpV0B
9kJOgwf5w/bfFHFUd4fX3c9tXA+aVjC78POK1RCbs+fWKCh2d0JuMbTP5jtuCSF3eF2nhNFqwuUz
TO18/SKGosQ2NP4S57VjyJ6mGEEl2dlj3QN3BfAfXp1l+/CwWpxAFLD6vOvvnQrYjOcDZck1X9B/
sYP3YukwFpwUhSnK9kChCGYQ7OtM/gb6Iw089vukzcYpNFPtDntR8m8ehpBdYQW9+I0FK3fKiePM
zuP4Pzz9VBglpd974EMTkb9KEcsf5aVrZFyOrZpdgAUVTJ1yjLfzEc/bF1/DYoVOhPevJyhq1EeR
QRmk3HrILOax85FZySPSCxxQzfVeYQe9I5E+tliWqesZxUOHJWpSZyi7cmx6XG1eRQy5V9613a/7
VKVRZJAbYHH7kWsZ/JoAov6EuSuuLVzzfTfXAsq0EUOfEc31Xq5rNKdoELgqMf1dLBydNk0oKtdH
zx86Y00F0AAy5HeoEu2rl5mqLkF65y1Jj9vNKEUm6W8scmcpOy9wWRvhs2B3GXWtJo518uZQjcz6
p2glJRIpUbNNpGTd+erUN2EpxOxHt3w7tB/K65CkcWqA3A4mPjNUdv3IBFqNZNVat6a/YWRTQLfZ
ljzTyJHtyE9jod2uM6UREBYz4vefiRkoR1VR5vPAJwefu5SjUw4uQTpuHU74novrptVdcI0UpeyB
668Ao0qCQS6n024GR19laZ0+s2HWzJ7IhMcHDU6Gtwj1mJ3BwYAESF3KbQM+L0Ip4wSjahO6YaaO
JQflygtLOntWnUpDO1E45AdrrZXkLI71Mrpck2qAMFmng5hVCNpv3QU0Dg0G/wGNNTwTveGt1W6e
dXtoQyMA1a3Mb93Es3gYWg6BBGe7bMWHIpgd/rP5y07DCCV1UdaUD0WdElXbcWKAVbAdccM1Xl39
AaA1U/TwzKbNJJCAOLPA89O+mTcw/lsAmyNTQqt1NTJBUXBODaoBpLHnUOahuHwVBNLRBeVX18Wa
aH+FjEM9OtLqvnggf5WszSiOj5hzBIzdoe9W8E78uHfzcMoec2BOqqReToS3RaRT7WrF0jfkbuDU
vDFp+ahMjA6uX1b2ajCpd0bs/YtqVs+nsz4xjy+Yd/VHdK8pCFWhpPc5TTw9M57y21T/FvojsjnT
k8apY5k6X8luqBuhroeZp7WnedizNnZV6YmyX9/05obMqIS88A0adBpTUJ4kqXjoGlHAY+PC0q/I
uzT4EvWzzqaI9jzxO2hJNyW9+btub3ldXVygMGGpeX4UZ59whiSRtsNvdlBZZuGIGq1GwV0Ob+/C
vvZ8huwyCcHvVSy1v/jL34OoiLDhp5ZHzhJtoiCYvaba3UQEMH/rZFWxoG6iDe1HL2kYM23p2Gbp
QSLxClk9cPq4KW62AzyBwvyE6L1l+RQhPUliVLqoicBU6THBSeBeLNOqkY4uTEn14Ztc7eyUm0n7
TKLHZHqyFtYC7mOXxJNTzM/BjynPolh1DLogsGT/Ul/Ac6xrx49N1J1nevQyu58wQK8o9+w2Bh+o
ATMOfOukaMFFpxhpxdfVcjd5S7/sZkUlwOTCsW9ItQqtKMYHZlMXWe31Dhv8wFtDWU3/N0py3O2e
HfDLMNUJBGjmM7BGRN+59wsFFAhStKseyw9g4P/t5BhpZDnIDvE67vWTAJJX6s9LSZq39uZwanW9
PsarJl8G72bRZVVOB9x68FvK/h4wb1Zqtz2DtW2O3tL66zhhjyd1GAlAi6TpH2tTuq/wtIPV6hqL
trqaHl4QovYdb9aza4HBjBJTB6aepP4gsbv1HeGlGmM7yjXtMTC9vPss6RkVMs+8GIlZ5qgQZxgr
vRiPAmFRNHZ8b3gfmvBwGYfIwBKDGyVTeETMPWLO+Y70yaqvrCfi+CF3BWH8gstm9zYyHTZ9YG8j
KXgYw21T/wpKtnSllLFDrHHsCGqELpG31tzhm56LHZSTAKh6nmlK/O/P8Rgv6QnpIq2Sgmd3dNwZ
cFmRJ7HJgPMsIfDK8V1LbFvQbaraTJdK6RISE6KucQl2fxoxS5e0DXzEONpBeYtnCO5lza5dQqgd
tWCHiegdbPeqovxmxMdhlZhJo0umow4Bn/sI3ZKd788XCIhetmKl7uBCQ+61FSZ7WqYYDu7ZgA+a
e9TYEtOkc2HWqE9saQQOmrpsI9PRhqJhXismusFqbDduwybn3LTx5uXZFDRMFShob7kJBFaDsOGT
4noD7a0jtkOTZC1YOveBR2wIU+60Xzfyz931sRlnbZyQTqNWuw/SBsPCt2wH5CUqTuvjHBEh+A5q
lht5GavjcXgyGKGSJrT3Gq7p6eGCfOvmDN69gcIaVJ0dNOeOyIhHB570k6/sVFdNEaEUlZp5YtJZ
c8eECCZhdesR4OPlYuuKCevrVrAS75KHch84zjg6FNbhH798zP4Vd/TTFTbWftnq0BMebthTtIuF
3JEPchqDU8siiPxLV+yItJiP9yKySKOguyc2o4LRF8AR5chxLorhBJDoa9SEPwc5BFSqNA9I+Se6
A2gxaH3wes+19D9GUmaIoCyjexdk+tkB4gleBvlT2JheUPBIoqDGyFPJKizmixDxq+LaCYXqGFoI
zdOvaQwihkjx9Mwqxbt1VyvWLDvGBMp7ZBdUYk4d0eYkHPOHZHbp5YJwIvnxFqY8GUmnLVJFk8eC
71v3VYriEaaW3DcOZ2eNB+sxTd/1vj3WGLVMOTyBMqsW+wcfjIZXfhr0r3cGbjRDH2+VOi7qO0EE
XIHT34IAFwUuWCiqoq7n1anLKJuDqn18GP24JVvOE5I4cMVSktozSjC985illQ41E8ssZ40RLGIP
OAUCbo0uFCzutcjNHwRnauIZefmutq4RqgHIF6ldrqSO2+8kNWhHE2qTvPe90DhQzYfSrKwd6Gbj
NsJqc1QT2OCEBj4lzK/kboynjUTtie8zLm0umu0/p3plRTfdMwmqbZ9MYNN5ozQw5qh3oYDbBaXS
6bzHZ9BeZdfJR3hcnR+sa9jRQD4xSgvnWtSAyNugXgywYZoGbcRLc1D6FVQhEnafssnQJQIcJ1yA
1v455ijoRGI85Ue6Rv3LxAfJN30WM1ohEv9tEk+hRYvUax8sENSxpoUyywgaBJq75tzQxglx1G0j
vQTpkcMlmzf7MrVcUAGP/PXTLHA6IsHr3Cx1Akxa8GZ98eSjSEZgqA3DE6fll6bXck/iS/woGdfp
Z7G7gX+1gWxL6szzAH/xl8Uu7ukQSK+vavGPtS7kH8AxZ6RBF9OGUCWq67/f/PQjkc6JsjDvoiee
i1jfi7lkSufBx3PSMUkx3AqAGPn2U0i6bHdR/HbR92uBKLAkIeNnVU58bKyLtxzajR5zRYJ+abTG
3XZjm9ygo6NupwE9Zmr+vAPQyeQ6YgMwYqjZPXa+qgKKeCE0rVOjDKUo+9KYzeO6W0JdnwxY/BQu
sIVh9Ll1fgZkHAdMbD0Cmdqg2BOYf9C8Gz/f5loptY5oiVzsnVlD4oF40u2WNSxryyjUVtJmCtRi
pK1xbEsKjEp+IyomgCzaKwQ55z7hVR9RKQ5lpdts9DI5HdavuM7/HIsRgSLV9MdZrAxUoZrGWNti
3svcK5fHVvmsfd438n/fEHWE+9QlHCL4mH/UQSZIrnVuTUkhKKe3oeW+2Eys1ZDlDFaNjFtRvf6I
L2bac9vgPt8fukyaX04+0mmBiFjEBzrZ2MQf13nWdpDmUCP230LDlASoc1TkXJYHw2pK8ncDGgWj
0bt5/mNCrCzV+mxPy/kN7lal3q6lf/DRM83Gy8/anVGEDq3E8j0QYa3Uaenqa4RzdP8Zkike33c6
YLZrTlnTGRrbODCwyvT7iamVcOdcP19wP/u0prd4ANJ0N8XY2VOEbDqNdNvAjaGL/sKm5WwE246Y
wyNm6GTEcosMF2kpB1pD2OQ9eGDyjEmcECM9CrSSVCZhBtJeMRyjf5uOcIJ2GneD3GXTd1dPUCfc
Q91RXwZox6TcGmY/nuR5CZH/NJ8stLK9ZRfqUrXVJVVb9X7BuAz8GcJSRKyipOKgr+w7qW9Wuogc
ZPUNX/6Hf4cLpET/Jje/s6bnhzCc7mVc96MU989R/1FSf6RKsCm1sU0k6uusl/4AlMFhQdCzKEcK
WK/6YiQsje54xkswyGwJVfwUAM/gQgMtqwnaES8+qej1iTgZJ8BK5+5tGkPejOvM2Z2eoxWtCDUj
blnEK5oDeGEz0rqFRSvh89NYsx+xHbFJJG7C0Xjp1EpQ/cxYrjtCvETbEEm6jX2y2rOjDtb1QUjt
LQzPTxge6K6SxcgDLJ8iU2AghXEIkqKU2qqS0ry9JR/iA7SX1QbGlGfPy9d2p3LKFwY0WxvTjKCc
2fYtjg0AZFG2d1uhP/Vhd17LS99D/tR+Oz0zGRTAFsCFVmUIs93srnObrpXzpgRMs3Dl/oVuiKrX
1y9TEcR2sbNKd0Uu6mr9qazEgS4i/XdeTmvbqu7qtVSnAxfLKKR0rlLiU47CGW5HYLt2f8KvF9Ye
UG3cNoETw3LfAxMSBoDyyFgBu9vT34M0ItAH2rDiEC28kV+dEFjS0B4AX+Gx2z2V36+K9AOHXQzC
QuO4QDkH41TNbLKy7ovsnGVQtSja2ANm4lD9M0m+gEnfqju/w+flo0wieltD3Qsv7VIDKVHXV8C7
r4ZiglOmyoljjsKAOA+BAHUM1xMcwNV/kAdt6woTI4uZxDxKl8CqD9MVQIR87nZGLuZNcVHP8sGf
w43DqMBYi0aeD61IySXItsm+/22Jx16ZKFZcc9JmbUnLlx0JkI5rAeVN2+ioka83C1WJjC+npvXn
x/8SZShgIGuYMhfC0SwJQjZKW8AjqY0epvjN2UaWdIeECkjOwFDXJGEHrbts0+anQXxYc79RIiIN
dKNJ6t2cnEpwCe3s7Q/CsrmSdM73OXVPhlJHpmyllX2wiM1EQWME8YDXGX89829ai6Vl3QDS23ea
TbJNMZS+cr1h/s4YRtrMvFGHVu7iXBdE9XeCO6/I/n/CrpCBiLoBUnEcikqBS7Q8E0Sz6aP/cKD/
+suCPCXQVdkfQNjHUA/7aGS/Y0sHStS+52vmgCC+3RmHcAu6xbjjppwgiaLBR82yVRBsEB6Ywyau
dSiNseR4FxX9KS+924KRHRs6o7HMUOX3i4/7V2Z0c91kyM4oKQyGray9vS31s16Y4RWPtAOu/UAF
Mx2yWp7MzoNaZJV0q590/9aM/yTH4IhbXoeC/vlAACPEec6ihAz2nYv3wiV5uaI1kt+oGgKKgL7g
AZKI9VF37r/dzj8WpqpeNec1r1X8QYRg4h3PeV42sLwjznWPZ4MV/gsSj8wXL9tK16DEUHwqQJ8E
R22fv7kWRDMVpCmUTXO5bAqy2BAMdBP8wW9iEi1B3Ux/u9yhmwnzSGWGAHkxEEXqiraPadvleA69
TzqbCohvF0wOqoYosvqKCsa45iSRt3HC4RI5AmDnrFk9DkPeWG/P9sEhKuKQ2/iw90uHdjHP4jx5
9TbUJ+g8jTRhovDhu0vff8XG9SFa4Yf4ueXCstmEMlU9CQbj45NJZ7N+16XGaWAYw28YjEwOSsyf
1kFMBobXPhsu43xPVgAnWVZcVuLM3k0NQAT9HTuUem9kZQfapGtMtP8dmb4vteG8/RaGDzjPDZKc
q3krAJu5YlFT4m/QACGvgGTdRSHbvmM1hvjnQDl506xJFcm6pmcWG2WHBlAGi1tXsE1bqn0szyKU
NZ2wrhmrUcGkUIpU+muxfc1Pvnc/Mi203ky3o/Vg9ziDLDPFgpPOiHq5DRLM0FL73leiKxl+M9mj
zImR7rl0nPFe4CZOYzJ/YwGhphMwDdpz/mAFF7JDI5ahOOKUQXSVeWyGr77tsDhM830cMwzU4c9O
DDRATIMVW+fJam4tak/179khVd59/Hep8n8BizS9yooqKI++SX/lYX/SBBKIdjOdeZ5UN9cJSUXS
pmY3tdNSDobJn+q71XY652x10KdGYNuHycUUy3a2S+RpU4yBD6RWDAtjS8X1f/zafHwg8TpHHm7k
6vQ6y+8+rgaJ61Fa/X3PbOuGllUxa+SeWndQmNyAYaQNUqAvVgrAFq5jvk14MKLN7mLUItOdBad1
GPPXu1inLgFJv9veB6BR91ogAQMBzXAMiVV06cvaj4ajoNiV1qvQhw68HqE5X9KRKBYAMUKP+JP0
hf60fNvYqTje2t0Jbvu6lIjFaoViVIWKI9MdiiKhiiA0Y03bz1HcK+srTa4eQNRC1f4ig48JWNpr
7e6d/ka+vD4VY+LCa26YDvqRsUbcMMHgn6X2Tutx8INGKYiwzbwQZ2hv2XRujALfotTWpoSw9vKB
J0OcNDwEgcjUtrt4fsPeGUQMpowm4yAbWyXfAaaPlxe3yn2Mhqswt67Vn3bY/BR84QwsdJLfWaeX
fVnlH2W/ozJtaWHv/OG77Z/Njcxssp0BgV4lDr272K0stIJeFWpNO2ptiaG0f+HaAgAZ1c+huQ6O
6Ac7Spy49JdnpQt8aNkUUb6iGQQrVli1HQbiE52KP+Ku8/rUocl/zrsupIgHuUMAg8sVgnX49O+H
cjVlCBq+JRVV5pQiPEHvNUDdg3QIFMcybrAdBa0e+3Kif2v0TwLUK/SwOgLtirvjqs9Pu94hj83P
iuNQSCuFO45DZwlFMEdJhvR9HZ18LNQy/LKhMUuO+MjzTeykP/MG204Y8f9vOu626a0e2gRuLaqA
xktoWpmmI0NLJKjACZP8RWMQiSuV+nAtC6fY2DiUoGSxzY2Qn753JWcsbjXt6lTqCUXo0+YFop8H
uwxx2qlCeQUfEZMRRD67itGZfw8dR9RyTOoqJYMyAaVjZU8wao+CCJe8rZFXdj0BT1vnRZUeORIR
UvjNlHnU4Wrw6SvDB6PxMQJ+gtyR5dX5AeYMsW5aVDN9Q4bXwCm1UaKQuJH/H3xcA5KmgU4TinOr
rwkICDkVd5VbnklkuJ721Zd6XWitS7gc6CX8ytPllEfdFK0pR1GQtu5A8v1dRSOjb5uuWtpCF7az
Ocgn51cc7S9UL6/gN5/M59IVNfNgpcGbwJ6AKOOT1NBvfKqu0xmWBD0DKJ9JRuVB2mNxBtHlI41t
U48tHBKNaE+iAC6mb0nSOyNNBSLSMCHGn3p2HTJ12ima/Sn+yff+6H2sbl+j5GCqAujooSG7izLX
nvwVV4aXm1qBS0/t5wr+cA1/RFVb5oPgf5zZP3cnJ8NQFJ7nPbXhukSzyqPvr2jxIq4PmWKXcn+Y
QSJ2OOX4iShTgaEARf5WuWfdalu/RnZR7Y8qnROtjR6yAX2JT3oy7PNNT/CwEpnK6Lp6TuPyQZrE
0F3X4YEM8fvAjmvXC49K9bKzXXThakcNnfANOolViw1Ci02oewGQQ8eHKHPM/6Dyz1I01MbC5Puj
PJyQMcehGob90WULVH+MD5MsYx8G1bKgmTDILAbuvPha7JAlpkBtYx10PpoxydBzSViZONPuWqMZ
68iZMZzFXzxQ2jYYeQNfZ0tX+Lenrk33/v+Ia6QjcQc3Zq3hpn+2Oebwh/ufsQ4InaoTSqwMbMhL
haR96bvDm5A5rfjnpwmp503bArwva5PDgbXF08JuZ5qyXOF4MPdp3C2wJdJVdkvOiNrERH3IHn+C
hf5j9eAkURH/D6EzTsHX9m0uG0gQq9ug0D1PvSFGN5mn70/H8LVMUGtF4ZVSmzh6hqITzaGW2KMW
sVQlsMZYF4pnMBxdPupcnro96wCV1xkfBqktV81y3exXTxm3iz0hLXWho8SV9HSBSnBmGyHOJcgI
uvUeJ9fqoPazn8/qAXXok3eJSY0jq+hpZr/TEhTkXNcPkH+f/0jbMYn96nmlsAH/UXF1DerioGvQ
48dA0thwy3nJaganwpbe9Z6nYUU9I6TSf1XSU2eZMvHmoL92bh9AA/sfI9CZgWdqn9kS+Ja//WXQ
Bu8ojubYvbOclay4KeC1KpIKo+1xKdyXuDSRY5x5Wq+LlVPGO41lxr39HqPFU+Mc8v4PniJRIkvn
5kR51IEykliPOLuZsF7M1a8+RpzERukUZJy8n2u/FkwSh31wNK1cewsVHMcXRqX9fbMCUpBg0DqY
bvAGwNt4cKFPhdA/vzx0w9ALJIgW65bHmbLsKyYySpzYO16J9cwDOmlH0RzJqKxe+pYzJgyUE/LW
xf36RdaEoh9ok2MYlE+pDbGICZyGf6PYYw2yjdSOa1wOVeOv4b01P7QG5wU/2pYU63ydUvFcyaM9
zEqCLxnTg6JP3NlKbMfH1CpiW5l/QKLgIcYLDYELc7/zMwuoDvCWiok7gfWb6PoBP4jc5cJ/Hfyd
JEe6CpeKxOcC0VIyqXAgNaKqo9+oiUY/kAdIN0fFzvAKRHUPRc4bhBwBttsM0cY8BGwIer1ImwQO
coQzJNKWFhMtNZygHDG550pbBtK8JcFZ2sBenv6zG18OfBoDkYF97oVfAvJV33X5YVz5ePYWitfb
7WCRlyJXuBkfPfFRWbaquGY0nQMx3QKmVPmXTAVWk6PowWvWXowxvQLJvf/Inh8u2T5IBFJr6wTt
Bf1w62EcDOEO5F1Y4z9lfjJjxoNfG1uwAafu4+1IDWq//v8CT7QJ5iWgbU0Lso9qf6EYoEJ3hOAq
vskU+IFthwc+rti3gHvymTnymYycwAT3d+6TUQkClMYA3T8s7vLfrPLikCaIaYEGoPRCbWZ4ls77
/qlIaoqZSWaYMiaDvrdW0tWeW6nfhtVvtd99lOS7Hjh5GhFnHWJVIaJB8WTCD523ZT9a/7cSl3hv
4fIrT90grgw58dAFJ3YvYrH+JcvvNF+VxG/ejj/0VXU6zvnFqCHYgXeV7SfZ78Nyfm45jN2fnmv1
c65a4c+nomcnE30/dIZNAC1YHx8O2IyZVkNmHvNz0wEls7ENcySu0ulyTyXlWWTFCP7U0/9bpvQa
GPJEftIB4GndMUGkiYJFlCc6xLZwB0RgNjvTaBI3QPFoYm1Dwq1TkzX7fCF4OzM5V/9ZW/FSdtSE
loG+I1W+PJ7pTY6fARDKs711PE7eK4jz0B35yQ423Uss4oRPPx4fsKdmif05k3n9P6PmVvaPhw1B
Gvvrh75nTtVN8Drxl5cfTRTjr05XBTKeo+HjOY7vZykL9p9Gal1K70n8pR9CYD3HpO06L8uCQPri
97TVaOxLyv7BC7YvO+DzMRSQ3aE5takwf6mVK37slPY6ic5ibAn4aUZ9MU1DbgnqUMgf2FG2SLUC
iS/HFMk1qTn+2XBNvKColMmqjYF8X5tOJiODw9jLuuWUSfRMxwgnB5Ig13ZfQG+/oZMOUHGZW0QJ
X0iDpEoeYCjOxBTmxnSzs5pnjgVpFAEMdLyDB1CduSCQWIhCj62sRcre91FZADyrts1IEoGxOMVZ
0ZQvXGRAgXFxErdGtYchrO3w1NjLKdShc3E7/dMW4U1qMDa/eILmP4QmhgBmjSe2w/ZDwoGy/xdm
PAilfYnP5JuY6OEsy4KmrrY5uY5i/ve7EjyxCZfkCQuzMf1J/Yd9PzYwlPCpuGW6WK30kw/XjbyC
82QnKC8playE5bevxstIn4C32doo4hdvGgQo5z8IXvG7jHSSranBT+KrgsbNkrSk+HN+a2DB/DTC
iVb3b4NI97f/0STn9K5sb7WwhHi4cWAcyS/Lb/9Ssz4Ips0sJrtk3nlpJXo0xZuSK+EXUV+MO6Gl
iEXZgetmIiTg1uFsH1Jx96CzqHL+XtL8d8Kk+Q7NV2TuCeFINXj0YaMbxOfxMjbOrGB+Shb1NcVK
DP/quvt4t3g3gE02XRHARkWnAezvfgMNR+7Ca8BBZpK8nAl2hrSs58R6VvShxuU92UJ0MlClfoee
kWGesVSsb+88OQI8NSx/mljl3ZfroVIQ1hKgrhVi1RsWsY63DvOwtfwcrS69uUQ5Tpr3MlqtKoRt
9wMYDlaFq7VOVvkkqAGL+Uqpbw8c+qDq6P+hrsI1XbVvesP6wbteppD+hWlJDznf+aH3wieGrO7L
YAwN3prgfFtpE+Sxh33KGmRkRHKxA/NeJ+7Ru+gsbhO6RNaAOE+fIbdOx/lMUR5xR1J4RuD7jNpy
nxnj3Q5m+PLvUDeG8vR4s9xhF0jDd/XOLiyjWSURWzXVJo+OH5KDGeOHxrgZs5ktbicF85KQSpjT
yUbVxNAlz5gDYq3lQYXS2hz/fPabaxVRVcBNjXtbrITQzgASh5jR2+DM+e8npQP4a5VSnqZLu4k9
FdbI/+3beNKBZGZy/e4CRX5fyKvtL8ys7uTlHhLZZSyee4D5XR9iKBtPoZHyjLmYPJ213IoE21Db
ei+Kpg8ghR2+6ofJ8rtXAQzH3NXVsZtz9utdNI1xePQV1qAMtjsK1zN25pEIfDSfASSSujNqbx8+
Ra2j4Y09Nqwz2Lwfgf8NvfooiQnVxIPrzMPbYprbE34EQe4V73kc5pPYu93A9TMWoGoeNE/XKrmU
JuF7Lk20Yr8XeqlcxkSYlGCeiIEMbdenpEKNb1VUvNp0kYZxQS8oLtm33b1DsdodOFCvBsTtU+ss
3r58cU3/fYBhC4sPU7LWcseBXyuatilluxZUC0f01HIRx9BsffIHw/IGSjiQhDD+znNC+5a0s6ep
eg+XNYeBQN44zkCHqVGfcANoSIgkCj94jFgDyXUGU8GXlN9Zvwware8nva3XgVWuiVxaldvZlWGK
Atr+rajEhRtAiNnwrHj3txwSDNamX7Hz9I+91xbf7AR8JuTLxCk9HaS31VkTJC6TSLB2TPtDqQfz
wlkdgOy52svUzg+ORYNhzfZrI8zaSGTfMlS76jK5eK4LsD3GAOycgsDvv0WWHZHGqa0dMttvCgqD
5VQdFceA3TKTbdcIc8hrB3lOngk16q6kTmzQ2RCUCfsH7ETiLbKpTavk4kIfDDPDt6HS9G62mwGV
xAFlmbIeQ/6PCwZx1x6VN3+sxnfRDA5lgEJlpYdYVxl5ISkB2DZ/sSADUxuQY5sj7AnJhyyD2vIm
9xUqm319PVj2pqNKMK4BQaQgi+1jlmDy6pCgWprB2gITdPobO3yGkWgS8bNBq5tIY0zbUIVkK5En
35GXFF6ZhznTmVWgdGydLMAujxAdbFMoo+8XE3wOjHg1GDE1ZRF7AnZB0jybpLhYe7sPodhjDBi2
mUGKs0CNjzRoh9g6LJABp9CgZQAlAtt0SD3DubosVOsdNYVc2fvc3RHNEQlBZXksEJNRwwWChsz2
dQ4KMeHy34ZLSI0v4ltWvOpqYqgi2bsUOLzynJwlKrIWutqIdnLo/0jlVbbUXaRut0ovyS2+2od4
hSPdmg7rkctcqC97tvuMN9XqS9gDbv0R8uR9yP/+4zLKzpuQc+0QU61t2HuO6lfOXu6XRJ4HyVh8
Qv3nR5OUaXmQuxoQ7vRmSfmJw8StmGHzUFcwU2bkYxBYRcG2akanKHATPAGm2nRh72XfeBQeYQcu
7rGpnBz93Er8W5Twmzi6WEmicw7M5Y7IPny5VZcR/YOH8JHUtYDShw8rbArUGdNp48uf/O3bS4/6
ZoHdeIvCevGShk1R5MjXuN8k34uH8UKvcLKdU4GMToGJZXm+l0rINpxtMLHNhfjhw7C1+uctwLES
a+y/Twgn758XegViBaMxR3oWXsq67VhzHYsE4HVhfO57n5x7kwTDdbD4ETbzyf0kBh9cJBmgj7RD
SpBC723jTI5vFm+Fq0AkJ/tcRQWwQlq3hblpk+5epXXIXWh4SGapr6RqFhdMefZF/Gb29YOifbBF
xD3DzYXU/5FZ22rfuo75Q6o1xraBbjjaHAzXqHbio6DJR513sDGZlz8mSQywQd7/7kOGhNVq2F1B
gzBLsSxIEaWiZvI2Gp0x8CMBMBs844Tzq0KI/DxPwNkv3c1R60DGhQhjiBJN1ugZFW1oOiYd/q1U
svTP1YQvu0XNm2ywZmiCzh7wlw0NshMX/CGI8Po8QZpyKpohPDnPM+lcUpDYnVLnGwX99WIQXFPS
ZthlfxSSpFxIcSFvaFh79QD4QG/QBP8DCOrwoXbwe1npwadlyAtR7uwf9cDDgKpaVu9KN/plqh6F
LUhrFZnEsc56rXn/cgQLaWI4ouAWIz9khpmYr2+pPGdeHkJyiChY+381T/p85nGsXVaAEeRcyUp2
XtH+chffVEtA5HOzX7X2G/BbS1mV5cL9lYorp/0BVhJvtSNG1UVWLgInFdGaHTqe6vhhUYX0cjSH
1+53t8+UIYIpHH8FJoddz2YE70iqpKSIYirQ0TDWs5vDmADqifdvi/yOWQE1T+TTl2yZexMZAOR+
tCeDg5qLtYvlVywCtgQhSrUFtpmjY8fu6moTlUmc4iAjcDgbkDTzbhCpkX0R3+31c+07ug9F2tya
D3Vj+yofuZmydkJUbKCKbPYScth8ry0HDp91fketgEmobBYbB8Ts3scMoah2JE4HZGG3aMtFiA79
OXHFnaPkz6Mx8pMpPyKg4HvfDZMiI0FKB8BQcwOJ2qfgC4QxqaTxXYNIbISrZHuwDsBBInzA04pQ
4XxCTyekw6p+MP8U5cNXM1gKc5R1khRJ+ZrTFiff4iYSXaPDfNjiOC5qemRm6e/oArTR8ysMD5vu
FqxkcA2kl6/qE1jhmHN5OS/giKsguNa2pMnvo2r/pwiuPN4IOCgoFjfFA9O6lTyuyEqQCLUJHRBk
o5fAGUOrbBUqku/Gen8PnAcB9WyDgOyiBYI6ko65s76lvRwqoCELW6Bv0bYEya3taFnTAmSZqT/N
v8pZjaF4R5RukcnKJzKXwQ66NxcxDfWnHe/fu/WNw6m7dTeEG2QtcVSGZNB+gj4FPDqLE2CTOCyX
Sw8CehMz2R9x7S8ClNoW3rEwWZ+isUuNxueKeBrJvtc0L7Yflg12v4LfESEwjBmi9yVfo9XPiGKS
cfB+FXEQYx13Fabc9oTv1UExvvgTXv19exohfvoZQL5GRmnFsnsbfrJhrwj1dU16yen3ojpuA/z7
hkcPZcznMCe0+Nm7xyvDzNFtYxy7RX5V/ex8MIjeTOZodtQ5hPT434Xn25Aae5sJRMQJ6JmXh9dN
i/UxF/ZMHZeX8ZpTAbwrUiJjOLuhAF50vGuWVTw0EWg9d0S0ptd+PMg/lTdLzLurAWVtAUud50B7
jTkqEg6suO+JFU7kSFXmr7VZZLVIAFzigDrTKEj+ErriWcE+kuXMXoQWN7KQObtvwItfSJtamjUz
az9eZqf57acece85WANVwpX7baCCa65tf3hUyLNGx+BbSKswQqbqv1fckv+vhYU0h033/TJGV/7Y
QXnAnh9lzeaTfKj1tJnkC4K/ranPP/nT0BrGNgJBACfbMVpJo2WuiPbagJNw+czEPBKlT5vkVOgM
k7b8bQui9RjgAW58NUwudibBrdNhxO+9z13ZyE50cpuhuxabXolir+IOUuSZc2PTYWRCDOs9EFkw
mQi57cIZvETFu3GoFQ3jqNfEYIgFlynuUujnXCk/IsC676gWFYToKPjdalII5+Zge/oJyoOm6HZ/
MJ/vv+iZWZBDkZohkBim7XoU9kbleZ9qgXSKxGGiiJJ1Rdb0l6eQBYW7m+V3KiEhVam7msTZXbwm
Ci8fD+IPLIYk5vHNReHGpfe7cEnHBvkTovjuymW4BIqrsYLU/SqmfKjuVr3gK3JmHmKUtS1pQ0Ps
q0hI7E/IKuSrF6tHZ1sgcgoJvpTN5Q2QMrJvBJmeLnIm37KQSRCtduOr41L9ng9Y98Oa0P6BJru1
n0DyabjeUuET35xHYevLKW/A9RbwfBXYf0vALFbofhkRnUne7gWj8Jmz3uOORYvfoOqdOZ4oJOhq
RqaM1zG+tk5Sf4zQWcExhzAFteDyo8u17C6aE1DErSSoJTkK1VNsNntxnOE4/jcUJy5NLw4TxlOq
pDKdyufhJpR6rfRNyOhCoDEPfkeBa28FTzyH9dV5RzMsMI6tlKoNJirs862hLUBkA0Sw2e5ZaaIH
Y5bE6zYqwzuZBtyGDgsPU4YpXf6NhJUsli4e7Cj7aAlxICbrY4HfThkTvUHuYvwNdxXr8ysmZNWK
u21j7Pq+WjsAJM/LEVC6aGumTh/pmBSyojkeL1ZAxmb6PFe0/u64xOILauJ6/kRDysBJofaVtycz
4oDhSGhj8nGWB5WTv+uOklu94x0FLT77sM83AIvci8xJ/LWotdXY8cFp2y2FFLCn7XdLkSnwkKFw
eM1SZymG/Q+N3FmXS/pRsaxLjNCrCPVr4CQFeK+1iqKYKQSrwM3U7Wdvw+BW4btM96BITmeTXIAv
93lFl7wHEt9u36ZwZmokdTrq254mO+E0u0jVRUY3h7mZHsFzyIYMdo+TelPJJhUpAAZ/JkjOqBB0
XcsuasNrrqHWAXQmfEy4N64KzO3j3ISVl+tghbR/mbH7B7fJbJFKCpqc+MAIEMcF9piB1yPVjsmY
oHxXquWkMCxT77ooiBgnGURusv2/ORv4wCHfvx8RFDVDAC9DugKoYQo2F3DPN5xjAgSXmsH1ccit
AgRf0EGX7EPZeJPZERJBR9D7St+W+agV6YIDWDspoc5/nyItiWfMxVsghNkx7mNYN+Ewo5wm2pjG
W7GbRkgvdl7iIaZamNzjTTkAgWbquDOt3Yud6Mf1A4j6YxwzGwkp/MCd2VzJ288q+FTDpv3Z2Abb
wtCkx1CWHkTtkYaTFV3T8GJzY/rHAis+0RaH0QFAge39x5D+osbRiGO+BsNVLdgwsR2m1dJyBGpI
e7zxW6rrzdQBiQR2w+EvmS3YE1OADnyjLjPNjaxy7BLEbCYWtvyO7/Nwm5T1MUiJDCDDjZq77ahS
gtRkHaUvwJoTtBbTVBtMp3Whi6oLO5Zc99GQ3tnS4hPbRuh7STUxA2PgOwkvCLLh6TaK9qIh6EIZ
LjxMrUZJdHOhfc8gGl8cfb1a1WaN5T5gb8Y4uAKdFSzzD5vax/EVpCxR2lbkcP26L53JaO2S07CC
9Z3r+2GY7pTy2uJhwH+bOOJ9qn+61IDSdVKCJW3kA/dJYGvqkut8rdneDLpYnRUE/b11Xu/aQ1BL
ZI+Dwli9VIzA5TEtDrhyWakwxwuF191QWybTPZVNGhbvO38oshKFNnJrkKgT4oE4Dxc+/gXXwt2+
TwoT5KVDa8Kh7i6Fapz2wrFFLAdarHr8v70GA/fNjD4CvF/xl44lu9dpEb1ZeJrl4DTHAG84k6PA
ht78X04Mx8YSLyZ47ov/QOTn1ou5QL76qgWtdLQ6rKP9nDlVxJlg6jJUJtkvCkYb3c6SX8rZvemS
FKMXK7fe1c6Ahz6BZ6ieQNntiZN1MgrwlQRs945vYv20obroZC4j8/zqrKnaeG8zZAy7AlXa/q3i
B4EFR3nbAgP6mwOT4q85z16HyfAoR+wJCxVQcCel4PiUZCT+3s/OPwBhGpAU4I5yIcV6GL3ys2II
fTiwC8U5U6pzukCJCyVZfIbB7Jq+yaijv6A4J+fWCtzDUhD+ClkmBxSy+4fM039bT5/d/QIVmi/u
dcP33weLHJmZFcRXW6WYUMn3DMDRwzTEteldt03vfYnO6YNNB2lZkadMmLhZHgx9U4NF02+IR7Uq
ZzaJhSKCI3+VF4EN/z37TzreXIAnkmlXJTH4x8trn3FZbR6yVCCKxMdDqd737SAukgdVETGE9+BP
T2O5w1YbstjDGXd+HP43gz7KT6qvgKFxQq5kGEJFUoV1tXi2uAdKyaV7feTJi5Pme50VWjackl75
rPsAnzKOzwd+/sr8/bBq4bbIRDUdd3ZwdPVI4/RGG434BpllSRWeJaZHHt88/8GLv6CXp9iGNDyj
JFaNkp0WeoMH/vzoOla/CohKK5uWM8X4bQyA63M4LiTfeWOv8VS7ryEy+qCvIZohyLbXtuijPU5F
iYX+wcCoTt0GmJi5EZ+YQ4Nw0VjSr9T73dPdRacjTztqQ43G6RME4NPf2XsrrQy4wtg/VhBobtFl
tMb+0yMVC8ryblN45bcrSSQC5+g3vjkF7xCeQO18acgsEnoERT/t5bIlrwAFtzPtMMyRSrbjHbEj
8aF7TjFla+PIqWM5ZN5ZHGQk6nVrVeov8n6eDNcUNP0prq+Giz3EBE3WvsW148oCJjH+D1h1joZQ
NVJ77P828wnWTvCNNZghxTwT83GhSAC6oKQ2XPFdOtu3QiEFa0Z8d8jFmygv125hWjn8cp2qv0+T
vXnBeKRgTCxb8HDcBNylq8wQkXNYysQ+ZTWvp66tfOhs9oKnkgZG3Ad/l+FD6TVGO3qlYWFWuQsv
9DpvPitlqOwM9OvXLpcJDFYFh+WC4SaYQyilD+qAohixZRlLLNtq7eKIS32ev1snsUKJK0QufB3P
naDV0y6PWrWCxrU7EsVjDvqn1m0UcP1rEuXj5iYkp0PEVycURlc0CqJvpgpcfiaBxRJ+kTtNZ6h2
pAQYn2hnXgBbtBZnxOI/PxXR7GEtmujmCiykA4b4n3u4YrsF2zrkjjeGOYlbLf4gt0nZ166IV+5D
sLw9Gt2mwlXyJPtk9L/owKC95AnoahjmQW9zHtg/BIZIbtJjpOBeejVwMuCVJdiDIavqDHJTX/Db
zDQnihn08GFAW5RZm7IaS+HGUftT7R64/hRJJUN2v2NKjKoPrKmVfo0vaKW7sBn1wvoQW19TAlN5
GGPEmLm0YluqZkJtj+gdZQyHMEc16QPNLJ8QPmXgpMFhoCIgOya4bS+z0A3W8p0GAXge7bn2CVj0
uu2VKywkKeJEDi+SUWpsEQTZBl5ZncOqBqilI8+gV1P07Obm7hzkItTkzKXrDKZzAEJWyBz67kc/
zox/fqXDa6HuZbKxd0Ewdr+RcmmvB3ztDuvZyXOFDCprjFMNrrASIGvS/Vu+vjwNoHnWlcz9LfoZ
BGIP/DSja7WXhJ+i9MylrSRmTbBmt6SjR/DMS6sBAzlcBN/CFjM1ou80oVEplNUEiEnqTdch4c8g
dRX/u+16mTMc8ekX3A1KlimYog/B6Zt3gmUv4QUCCgqU9plHFQibD8b4mu8Q4p4kx5NapRGfeu88
vxLt/bMhujGWHl3624m9DIqOBzqt9UsMIptM6N3PkisCOzlReo9Qxoju1VNL4vqCS4WLMvKgad2/
brcvn8euBw1AzNdZ7LaAwnyO+/cf37nvpXl9h80FZTHZwSMU5x3B6/5mZqkhq8j59mU6bkLXRHvV
Ke2iHKvqiQTq6OuVR/uYjE2Br4icT55xRJ+VTzoXaBB8zV4GC5wwZokDZ5mbGuqu0OXITewKjhdQ
9aFUkXYVB2dbI9IqebslvTJlY24B8NTsYh9gAHku+FGDDpBU2B4tZmhiitj1omkoDRMe0pBBWNTa
a0uRF9dqsvu6k7LOrO8Pg3hUzKFmO0AluxlmO4kPXBOWhqzUDGxQOwIrTRsamFy64CVhieCmPFz/
rFkhTIg0j1OXZC1YmHMynLdWGiG+EfPXtofL/RajzTfMah5vn7vzx0bLr77YlazvDiqoEMt6sa0n
AQNBuLDV2Av5AceBCrscWzq6eATW3q0U3KZnvUBr97aMEKCRDcOHWc8x7Be1R5CO7tcwdVTKUpIE
Vi+cdvi1y5SapVoIDIC0IMJVJewzegMV2aza7kVVAtWCVs8afT2kcO1Lz+qsZf39z8vHqGYy/4EL
YQyBeImmcBNv+Kh58uUjGjojT7yp4XNvsu6dgIAS7QQFfr4jyyab7PnZ8kZMbXXDbwnF73s5DWE4
+fHeEOfr/tDMCq5WeTRQwMkYMl1SDJMIU9yh686VBXZNJr2huaOl5szKIMHnjHAnUyWTRzw4mP/1
2M9kk/kr6T9wbNZMb3WhfuKtVEWzKcaJPbV3Oo0ORxr+Y+pX7Y2HITVVJcQzx9DqN8tjnTSPFCoP
6mZwW3s4GNJZwA8n4prM3OhxKOLVdgnC06JkZGmIT1jDgYc+uzjA2x3z0/2LLUxVTL9uKcamG8nZ
iIm7bo2y8B8PXSKp1XYpFwtl4xJmrYIPN29NyDJVE4rnlU5cPydThOm6uK3UUeZc6snML8uazFcN
Ngu8X6JaN7FgKvVmRD9NX8AtaA4QeBIDN9INI4dY78GewuPqqMLw80CxRNSZ1ar8abkRnJGyxyah
f2Te71VIqwnaqKwMI4p/1xb49kAR+wpWecowcms+BUkq0xw3YT5dLYSpuExmXXbr41wm7HXcnmV9
F+s9/AIzf599+JqL31cKQhaLmXTwZ7lO16Vd7lTt19r4cDpplIeIN/hC2ooafEs1fsribWMqBLQy
XXSDZUEcqU+mdvX5FaDLn7UqZaaYXnA5InPATwTPSySfW7CQNj/SHQ3otis6eONCqtLt0njZ+Fap
hL1t544p00qNKy+3plj8bZAjC7ORWmiVywobrPkhoAuLOiKpumNG1gpnfmLyYcbea1dvVzt4gg2b
QZp8PA6/w6KbtmgsghDnq5C8OLy/u/W1Nw9VdJJwXnCJK7O4HW6r4GX9odohBDptr/vi3oEW6EQG
j6MO72/FKGnkAGbsvn2P1E3Ov5HmFgYixvDeSeslE0DMPNBwM6Qoekpy5CFNdXiifwLTwV64e5iM
AnOHyt0PQbkpzcNMuTedIBdIwLMFAPhMHX5J0LvVyaXcx7Ld/fl198vtL7NilSQCIo0KZMtJZFLu
3NZS/NrZ4xCTS4sqYWYkZY76k5QPkJTL7cBrtlKUQF8ZTZ80PiK0t1NZtVlCWm0NRP14uX7iOsmY
pEH5CRLKy43GiCTlWmgJIO3gJ7KxAzek9zp1v9rEGdbSkvWUr42+odLlVjiINhPoSWLl2JRmAUs6
u8qvST0B2iwC+qY+K/fpHaTgkaz1/w8PSu4p8Gg98cJMev89apWb16ICePVIxJmhfzjmUR5A6R7s
HUmRhhZT8KAFmjLU9hc9wHf4vBvg8ph2BlVzSDzYktKArxtWzjs+Udit7y3TAghjynaGyZ2u1D/7
78VeqdIQY/YL6IOWe5Q6+45ry1ekNK7/TYOyoEFxQhEu+Ksv0KJOz0XkKEVKnQWobsv3/V/Mz45X
L5+LvddH3Vm/wbSQ2isTnjf4Z6k+tPR9vJ/n8sW9gEWdCGB9hu8PEy7dhUgEKQfgiLbTUkfBjtRK
HCU4YNYayx0qNb2p3iTxNLHhgqdSWnZON59LcBqqU+H87E4ip/tVV5R7A2cGTs9iP/iMhOI14Mui
kCc50AG21nIa3gnQjGhcmc6olEipmXvmSN8KPLoo5xi12LDzJW5AtyCCsFBlugKlpqciEU/ydXyK
rOsZzSfyDOoEz03ntXFbRjvgcylD+Tv72dbk0/aDEwOCoknn/Vx2zy5futXfVaLpx3WYlAIv4N2q
HakIQpe2qoqRbaJ1Nm3PLU24p4qWzmNuzZTzJ22LUZmsfgmKUT3FIUD0g4NEi6tXTx1bMnGjsTHa
koJOOeZiLgqltFD0QM/Rm1/eCCnuLJAGFW9FWmT92h/ZITGXUJRl0DZBhNKkwcOd61bp72IHU9EB
uTGhzC/DKeHT1MrSEkapoLkZiUxe5eTEIOW6EqooTd5VU35ZKd3Q11TR1D+c5hZWyveZCyqQuvD8
DmtlUQpIzwdOc4H7fI+FtMWuHkmbytVLqTR/sSbVzvNnzZon4d+ZIzFrybkk3vzkSjCTh8kIx37o
hldgF5+tojbwiU7gc8q1Z5yPGaAhRuPBKHwFd417jYmHRrjJtodVFq1bgwxZqhNXUFSObtiVIEQv
nl9lwS9h4DUVuFvtC9N8mgh5jGzs7iXqpUzL6N8R+C8dQEvHgdXixeX7YZ6Og447Ap3cs7Qt3Q5e
NZit98jjilIo4vpf/Nt283nGsIY56Y5u8lISqmIW8qtpChi7c0MVvAkxukEURiT9hR6RNM9fWgt3
2YfUKtDy77X/ZLox0U+TEfZDb/Ql9z3PEUvALBg26X44ccZQw7lKIH8nbEU5yYgUP68kluGA1dMo
TsrJNyUjCMFJ26lxX5flRfe3xN4CJegFj3tYqr2QtOpeSPEdvLJNU/9qhEjfHKFf64WE2m8tZkrH
Erbfwg3FGu8DJbNlsTwaKZbBRXVcrNczxD6h5tDOFDLe4gvk7imAxQVzGlvwq2u91wCc81vLuI9x
r0WR7gvHaCkxtnhhxyA66YoFxAHVzRuYKYTX0Mv/sJOc+eg1rqBFxSR2dewGXGhsF8OgaCM/yePM
NOG1rr9tki665+AL8rzp+HywLGguLBDKpExaO46H3g8bo6rqvkSUZs5a4vsRcnJNZrP2UfLa6O/+
pdiZjBlT+akMD4Rh4lpem27tgtf+4AMfz9qcb274JtRWdLGbDvsfjsxEpwno/UgLS0ApF9549Oyg
hSziDi7rUMGn/noASuBpnU3KpSl0ArE0gveNwcEZvguByeLFcVeO4HOIOPeHRHaqtXhKCIIgMSn6
fqQEIzVHziUsttsyU20hdVoXfeQf6rfRRsKMF7h91j8SjQ3nfVCi9G1QYkgofYksP3Eu+vLC1sCf
dx0BurcuBCoXyNd7Pk3OEuSny41kkRUFsZLJcoSDVGLSpiThXV51rEG3iBm+ZD0xzA1i5HKk3SKk
7gpNXAqJD89BhsVFgRAvHtSnpQcpU79RR89zvg1aIBeZWPJic4WVqAQjHE7/ll3gBTDZABX6dUYx
2dwYiyRM+jMCXinTOTYDFMPKFx0MD1/nvMtszMO23aZ6F7Y1KJgOOoiIdu7pMP5HCLpMlDTSWGVx
+/wNpL/2I/IwQ3IPX48IaSFmjB2FqxjFYpM2uXfPqSaoc3Rg5/wyTfc4lJB7U7jZuUgXqj/p3KY7
wh3++Dgk8zTG+yPBX7706wzLeW2avlQS2kuxP+tkfsftyoBUWDzBj6j0rBDLkJjsb8hsErHaMEQL
aA9hF5aH0j0i9O8kpyAUj5oYYA+fGYEuPk7ZUWmL9PJK4hI3cNNgRpDTw9NBh66y5+o+hfQevuSF
9mN1zKkrRhMGq3L8HXorEO+df+GWVoXd5r1BwS6HuneSQ5ifle3lsRHxFAIm2A9iWcpjNJJqllEu
zHOxh0f6jYkG70vVK4E0gdslKdmPGGSsY02K7AG/wj2D4XD/3NRZSefNeldcqyfLijL73UD4s2zC
qCt8S5lNaH5Ufw5mKLj2ZeZXJV0hyAEGWG1or/zljlKuNEutxrl0o/ut/L52pgUj7mD6ca/tVQka
Jra7Y+1fokkVB8GW5sjS4vIQ8fBzekRVUzlWZ9GS0vmFBqAE4RehgkEGXAQ9a/X9CFcHseGoPXQV
R7PPmBRk+/IVxC/nThq/uEpq/2OK67F0UjOZp5IKFVSoo5h5w1NMSlbhDek/mEkuJK6UM5nYQdc2
Ba1vXY8RK1jFjMv4nfzsJxmJOl9GhOM1l3n5R2KtAt6HoQIEOVHP68kntuQ22KyIZLSQ2jrbLq5k
TT9D6RR+Jmxv3T9xUWWeBH9FxCmvVotg/7gTecH61dTcDr8yhJMOyJZM2HjNbAhQHNVHssEvg2OP
ueotBXO49pmkcqi/P+F6xqAHHE0WqbL9tSwp1LTHWipJl6jntgWR+S7bhrKV9Gh3KHAdywEkbj56
Vs0umhIELW8X/nvgevojezLYYK1dcicoKkJ9fy4/caefYQQxL3GU2Ykxn8lclw047YTF6jElxTJ7
Fi9qJqHp6a05YgU/g2yfRww+3orgXe/+SQKTeAd/zv/Un5wwLL35/lN8Q7muJK05p+tiHHdlq07Y
AVo5YktCH3wVz+3GvFjzqcy6wrLFhfNUmPtNtAWir5RfwTuD7my+uz81xxb6oX/KNfpaIGIzZ1tp
8em+RTOL/eISaiDF+ZrwZd6ET6ic+wAWbzEV0TtAyWHwbwk16+kcg3RlFejgdTXYZSbbI0P30Z/v
Tf4OLUzB89owjZB/6M3A70FyZrJl5QDYH9tVYgBiyLldITO6Z/e6tPSPLDLst/51wcHll9ekzuqV
5rpTz5E8e/pa5a6sh4hW3Iu78NkuauffnNSDm2cKhJq1+WKN60VCQgjpsbEWDEwQBubTFW+AXOWt
gkvwsK5M6vnf6saXwnL63lcDUqldMCYIjKaYZDTZtVx6kBHeRbF5jZdaTWhAKSp0ivmz4LlSmViX
XpzhcgqPzJLJcvvq32fAFuNGSEQuU0tcNkioobMbGAbGw2Wlsww0zkJvmk86ogWVRntVvkO2ekuw
mXHEtVFFu5vV5tDUiYs7MNX7nFKQvasiw/ZGkp5Sq/cbosE1Dyw2j9qfO3J0Mfd+F240T5+Vo9bs
rMyvLzAUyee9D/+0d6rxROXWsltmAbKdZMSV2ZzGbTTyd7H5q6LxlXG8/zg2/XVsGS6dMRoAmEOy
e+f+o5MU8eIZybMsSKuCyXmUPSIxT8KK9NIGppOmkCFP0usetz0PUL5G8iBeCKjlCiAfmEoFJlfx
bpKBnJ07X5C2ThkZgiJoAZuh8n1M5VvkE+qN0ze4XFtnNDqUTjH2mkD37VMMY3uDVil+aNTlZGIu
jx1xq+oxNczkXKZt9VfuP3Mb6/7pdlUcR00y1KaI+RVfJKvwtXOvqGPddq8jJ9HGGmsizDC41w4d
SqVLfaVIHzD4pX8KwOUP2uR44zmuIM4C1+GUXXMlhYD2luojaHZs4yGtmdOhm0wOg7a+VUM6SbS5
Quk0xj2p9XWFs0oI6MonJVYJYyYHxz/0PFTJFZZXhEPt1cMff9gHFgWmr5Ybr9jy4ZmQwfczCDx1
WPBxoXftqgfQ2Zt9SBm+fy0W/Q6HPjsT9CzMWmqYD4fyRr3IvVLVmCpM5knNVugcbNA5wbp4WfXk
GaKg5L/+FTk4haUhPacv8Vaxh4D3M39FIrYKEV0BRI44SasIV0Js+ZDbHfcOqL6GsmmJSfE6eoKk
ybPYIV7/CfpS/0zWSa1sJTrjvj5tRIGSt4A8Nu8i7PhlDkrcyj9+TH2+S7c3UAo6ktkcpDLYJGxD
i7/QnVgjXLeNvw6vpI6bR+Kru6CBM6/XczjqFLKUWRvT6mWnYqqzWxTmNh8IRBjMJ+ZDspY1YyfR
/YFyEEvSz+NIgi49dOl1PquGA/IwK5V6b+f7W/HZDz68eS2unICMDcsEGJ3BH+MAlUbH6phv2tPs
lo9+V0VcTNlwu6grzS9bFQXyNYOQAXvj5etjRvtFSr4/oCzD8EGS4ohUC3QdtOJQp7Psip//wfT+
J8r5cL3eHWxR+0/Ni44EJBJ9WAcQVk6NwjPwpruESTASqUW1ia0UXrTf768LdKpS7MIIaBHvarDX
ny6Lal98e903EELyGW1NssL5+66dEPYA6GVDn5Eb9CdD8EjqmKnJmn1qTQgzEy4HoR3WFNz3MK9s
gzC6ZyqtkE3Pb6ulixum3eaT0hN8sDHFCKap910sk89vIhfuXnbR4/pQk7VIWjiT6BIiXIuaLjWX
XRjFy6XXfZ3HsCNDi6hOQ6ZSATbHENHXt8ny69BTbZYaMZxkEW2vzmtsC6ArDFQ5MNPqA1Dr8Oj3
CIXAWOeOfhhcInuCj3ajGjjfdZYBScFs1BVnCbEUuEane8whvAyArBTAsSBrNzDr/gElBs88L/AB
ccxyw+VWl8jzjiXVAYoI2+sNxBetD6H0ptH0eR4e0bGzbWw3AQKGV/N2sjktoTxDtScyyPJ/5Y0U
t2SYT3Ma+6efV+YuCBBVw6feJfhb5ZCCrXbUajShz7a791EDdYF1hrF3pwZLbqjQYv24JroeCyeO
QlH6x+UEFhEXginBl0CNIsM5gJsHWvfpoNyUsFKQEaKrpL9j9B8xkUQZfIUSMl+nR4W21arY4IiZ
hfz2W83HPG63aGRQPDK5Td9FnIySXLl/UAJ1CKDCfCrLJ1zFPMuXzPpVYiE2KfH6T26frMehhXLH
wYn0vRs4BxnYPLK7cOuzD3F4K6h+RFjQSuWOuwJNkktPvhTZHdzl+z8SlwL0dOjDhWrFivTBQvld
z+TgVxlbdqRQtMFGwV6nBtg4jOmt47Ph8ZrJnnVxa0dky5ai/A0j87Z4VTkZxAjsCNvRS8St4Owp
H3qcau7KH+UHGXZk13FOINdDwgISuz6hbKZUYhXDzPEtIXF4tQXQrOnjp8Y22lLF3NVRlS5cN7Nt
Y5kysmFI3n8/tQEyLWGZQQYKGmun6DRczqy9VyaFKtF5LEb3nL3zjgnrddjTMYriKrAW/gBG5F5e
DaNYM5dSaAdsIZAEibp+K+xMMfIYDDsNBbsdqvdjpaq8IcNieh2CBfnxK1A49mAdLAIYg18N9oyM
acUSHOjgz8MZodGJcMlBBTkIC50vZvg9yf0mB+ZvLl44TsTUjqzO2KwcavZWwJbnBSr6Nn0Y1bs2
wlnL8F7NF3nF28cvEKKhC13++IU2C87ep8+HvZnZR0oK6B2ICaPwVw4dcq2HFIG83x/TM2bvLCGH
/OnGj8zDu6gZYV1lEyqZV5V4TYIFgyO90YRU3aFcCyGqB0tspXwm+5GLnZzESgQjV44gWa2YcSyv
UgNZoZ/GH636op7LByh+ccEOTXZppJh+hxD83ackg03ry8hzaSuWcoOMaYF52As3mOL3tyG5yUpx
NX6YVMWjDMSwms+UtvFnYoSNAtQC70p0mVADt+i3I5xdcJ+lMCAJ+ZTAJh0aHY+aR82Aco7AfrGZ
Tdb2ASb1T+M1R4RYSBT31b/ebNNGFsyYiM4xPUDbKvXQLbx0zuV3XZGsU6Wh6yNzb02IBN8G6HvM
92ZEBJRCkSLVzmeCXvZvn48KT0AhLY7jmcUFuPSi3Gvphsj8DR8nDs1ZSlIez2EwunAiUYR9V5+H
kh7uOhWKOLYIhp5Jf1jvc4yoXWDa3JBY93xPy2RA1B3b8yFg4GWlgq3YOls0VQSAi43cyDgy1pq4
0Kr+deSn1zdruBiZcN1dw+/0okQR0Xla4zTij/6bjZdB49Ly6o6ChH3R+LNJFxHea6ePoNsO7/iF
66likeHaKTRIENIcgUp5+AM7whFR3fcD3+XCI0G7FJHk+susnl/EH74rYK3pXKPqTLyB+76SuD92
PEdx1yzhLrOwfxHWqiuQCD87bkJU+auMijgyvelvB0Js+cFYf2fl+dZfGPrXAh5JZsI0NyIKxprF
5TkUnX2UTriAr6CsWVsVnRgsBLSkQt143Ola4IQWs3DKErz4zMQX7+XbPYn6deMTFEn+cKF/Aa0W
4KWIsODMGwyv3EMWhK1FruHw/dHcZ1NVcGx/wlK//hZRM36SKRxPduRHb+w184aXWvi1+MjsBsF/
SUXKXfQTFqnsfpIn3S0MJ33Vuf1m5zKcbD6px6Z8zJ+uPuDY7x4LVmVb4jrQ8mowPfdBCFaGbDLj
QyihcFvfqYm8wFl1SWjSrDj+0s+wZyY9tJKOWCfy2KQgqEHuzYnc0nYSBYiBZQfRZ6rIUQnLK0hd
xmgLMAVqus45NsEfQCN/KqtOCXA0ubtxpcj3mTNi139v1UHIepLWdHmUCijL30BmDNDkMgrUNV4M
mxLd+0PsI6dvJ+03PxUdiuusv+E5cuwChE0mvaoAHWXQHR9eZshIii31XeqWF84mljsNGHTbZibs
S4+2lhQ4pQ68e8z4wAh1zwxZQUwV8T3NeyStkaUibpDxslb51RfQod8jfRFKAL1VQzazN3pxxXlV
/L1e3prvpDSfvXTXltteiZ2mAig/OzXNbIdABYIiWFkNuLNUYgzm/ThWhgn+7iYi1izjIDDD7aTo
g72iaVlnbmQYxHrTMXFIFT0y2WyUbtS8Am8638RkfZ/i/nzkPd8N+7XYHVptGG/Mt2BLLpGDzhnD
YQ8RRpKVPosg0wwylJgf5Xf9a0boR0lPJ8oGeMMg3upG23VeENdFrMlFKyEQG3E2sYXdW9hAg/QW
umVIbxwggFhBpG/1WOhtpEVA6xn7oMU+w3oezJjPJ3LQn0DKN11CnvtRMzBGFMu6hCPO9ODvAHq2
zTjrOxOUs3V6Ag8qjaGqM+k5whg9n8moJc8kQt0eQD4RUTic2nlBtVkkrHur7p3ZjgMxmy7hFA/u
oWm2LSRH3TTsIbCoMHqZZ+dMtMVrodE1HafSUTCXbcia68w5FV52O/f0xVQrsuuPQc6cEGEV2RdN
Ds6f7wU1qK1CRYKSYg6rlDkW8rz9MrOV2rJIsXSbcsXy5qCc8CfRCwAYi6jAOhAKJYTviESJmk0+
P+5BoQiaO7ni9PMKhXKSTm/A3RgF5DA3RUycOP1FawIG1rc8adIqADJtisjLB5pAo5n0Px+pU++s
t5K//SyGdDZwnImkKBeCnWjKEsCLMmMGeeQul+KbWYow9HoHQozwMHs7RNVNmEW6EeUCpVkTNCyU
+srYv4x6vvINvG3nV2nuli+WIprhLuhZlQXUOOr1UfoM4IbC9/unmGJXl5IUNk7CXk4/kslsX3zO
WgReLlGePWriK1tpFWvkIyM+yfNfi7biJGtiMnA475gBXuh97f7haL4RQXJMLARACk52qA1uwcxF
kWCVTuq05xqaXlQ1qG88rkrQ4qpTHthZss6fLnfDqZ+PtZhtyylM0z3XdywtL5SCFC+BTOvlIlBM
9v00JbUaB9HywwyQhzUHgvtVifaTrmz41314RxLfOJCIAxzSEIpIh47pCyP3lOkz+jbDdwdFeZoy
rAwos2xa7X91fMh8zA62IP3MZwtZd1T+HCo9Zdo2y/1FlqUeKPtM9Mi/tBwEm+KCMTkqhi1ZOGUn
4B47m4Mr7bb+a5rqvbAlULy5BuBF7qvPpo+XLudCtiA2arn1ww/GT82U5GzpcY0tI/nk9ymCYgSG
ilnjAmWyNfSEgP49CVuz7Vh19VDYqYfCbM7lyMz/LELbyHriv+fDaX693C9MaeLP4VgaTC2LUVji
uaolBB6mhD9pJ4o7y8/yqQpJbfblQlcVDj9ANKH3fuOVI/K30/0xLrmONRnwg3wAJbfz/tuM7XsF
Tmz4SWDHVyp3gyIHGQoh7g5VJRqU47xvopSXeKBnc0H8cHzY+s+K5n+4MDg/3H//d5HE4KzbMT5T
/05b93QdIxOAdfJcYW1FMBQy4WFjDQtrL/rHiJQp3baAXFZWY2ZS8fkr80PBTVJo+MrSwwdIEhGP
MPKMvaNVO6meEnAdGpjuTiy5cYTtI8BeJXWl7W1pMVhGrSzIESeHIrZ6U42+YhltG/pdWxUkUjuU
vHZ9JvPMOHsvwF69jMBcb5ZFBOWDN9mQTlRUtybh33BbOGugA0dxFbI8Ix8mdGfSMSvpMb58J3Xy
FVGjSFlRUK6SDf5Y1ttO0/u9fOxX29YfPYu+oq+YglqC/CHqZvBnmg6JiyYOnKwmfWwLCL0/Ycfq
XLikD3BLSaUEFnmxu5sowZ8FsMy4vzts9tRHj4CGIwrLV8Up+drwBzfi8H5d2gHAooIpXUDWRKWC
9ix6nPvAicQZy4kG2A+kVqN+X/C2noU5tVyx+G8JTGnN413Nr37cCO954GRv2mw7KXc63QdzF/Cp
rQTcWgHYrWRvUT/qdvWmkiPDFpAKfK3ApWsBxYD9xscghbJOLHXYDrpO/MSrvoNSZ9zfgU1+Fb4H
ZWJ1x97MievVqFWKPs4oSDnETCZOtvhWfkS0Z9nmAJpRG2sWk3ncm5jO3EoLMzbWExeN/cpAD8+D
c+ITRxjtOXtU63Vrk5X4+sOJQAUR2P+RpNeIK5dae3CB7QO0oByNdSKfQ6oI2o1dUuOl9Ink6mzT
yOQPVxwCIhkZ73jNBpUIXLA49E5+1gyx8ljqtAi9YZAQQeypHynp/8jBJe1FwIqfj7rOYjsnJ/cx
icfC5UaYjbeCbOoX4y052dIIoWD2RWwLVDiOzQvt2pAHm9Vg6HmHvL6v2SRWVboJiiiwSrswXSLn
TD36BLywBMK2Iw9gPLnLC6YaKajHSKAQBmwF4/6oSHajF61stOC8DcXQPPAW3sGMuwWQ4NjZEnrT
Ip3ZABnGFbgbwtiXb4jSrvJN+LJbADC4sGg0xfuX8vbofWJ1tC1AQvJqC2F+4wHHtKGWbqCIMtVC
70ajE2WLWGMj89cRy6oenA0hoS+vIQMN7VJC0tnErbJy32JbR++8vr5OcvTlihTmFgRgBQ69rQRr
ZjCV577ZJoqqizbW+L3zG0pcuwG9Usq5CmyYB/pGSHsDbLo9CTtWcbFvTeqhgliU5/v9s01gx/4B
sfT0NQn/4syjFyACFovxbjFKyr1xs33vpn6nrSOcUMkPr4UuGMKMOEUEx7RQclVBlMmC03kOaY+p
D/o6O+JwsTSXjlUkKXMHtbc8TW6c6vWMXxMx/ngxgWQxHvtwTSOQxKYOdBhax3iFYIyB/3PGwhbl
3QO2aFfRU44vGUWfEr9iILoZ8IP5aXuXILMRQg6Y/f8fxxDXJ8/cJvx/wCoi5aCGG/cbW+TzzL1c
qn4ZIluuSTh60N0aC4HqNbofp+IJByhhNCsfYEmaKgIMNhGsAeobB8JSunexzSGTbTyB22AGcZCt
XTyVbM2c8zw89uwrRQ0LJ2qdzTdq13kn8gOs5RqmR8KCDYz+OZ2IiiCFMkD7c602CPxhRqrQFKuH
RWoy308/m/T1X1HU0QMSqxlvLTq/JZc1T5mEkM1JoDv/U7Cn/0tyUsTYN0mVY2gr0FNe9OGwGa+I
Me4YJTdWXiuGfYnqvWYJ+N8kQNY1AIPPhmWUBKIORz3Oju2D6JWpWt92sW5K9eQQcMes1yZnheMq
x91xIXD+Omb8sjjg1yLYwismkHwu907/2OBkJ0HgptZScZP7oC43bCal5ccvVoPzx8kpaB9pYfDJ
a96V6eHHOf7gqlnzmt2opSecKT+JjmE8ATNg0GPt5BVpNK27pxp2phV7do7x2AEbHWZTvc6mg2BU
JAN4ZPG8brNxEcvgnoTp11IaH8hesg7R38XVVaqHtWBZZJMLh+HxWu5WS1AhxwDpak51tUa3rob4
d13683TdhqJifvk2ulFd7n+tUQ7J4wOS/sX1/xFTs+9n9XPy4OdTY4kO0juUr3PachOwbNQnd5Ab
OB876kdVYmdiDSUrAxWUaxBfSyIHENC/7MvxwbWSQY4+v+H6maI29Ri1JrLuevP0w13m85xKndBO
Pwe9nq9KWstjO8orR74s133QTP2tfnPkq0yp+54LSPUIVC8Z9KNUYfBht2IiInp+pQQ8KwiYT/OX
mv6BNAfQ0j+JGVWhstI8Pw/PxrH2SNol6g70Vgas5Fr+yIqnoxRwsp1B9XTEwha+t7jR7f9vsxGS
GFkCqugg01cmQ6bseYN+H15JxlwuHYHNgA+FGwv9ZJnRcPdgxSd/RO+oNLCESMfqAtNzRTdV4qlg
DNiMnuJKzx0rgQusxTD/l9nQTo+H/Kq2bzq1rA37JBsguVYl8ykZlDWigNPa93Ar807X9ELs3xML
GuNSPLtjsrr4sqXx4/UhriirqNPfdSFTUNyfsXMD+O7pJjdwL9m6pHT3OiqlU2l0oe9qntEfcG4a
ODuDCIvNxB1nCnqBg2dXexoXiTmRESGz2HukY9KOmqoJdrfA4bCFWJLyzR2D3/yd5QMLTizoIWiJ
0BU0TvOVdQXSn12Rs13hgvTdQUEhFu4KD8VaEo6Sx3Rh+96QggwuidDLZPD5hz4U2RWwx8Hxa7Vj
kg3mBayib64K7qRU9f5P7Yiek5j15QpnTjd8kA7QUebVrVvWTGKGSzIQeOJicl9k8fH9ON04c/lM
k+fgsBb6Nt6PPWno+NX+9V7Crzfqm0GL1qftg/zsxE+VitX7gr606ankeapWjx90OOERkcIxVzEK
SnWMIXgqYVuGZuoMXy8TlLw1Cv3hOyR+rwchyKQ6khCMSWe/iW4Sv75S1e13zAav1pi7vPYEfad4
bbWkDIY1TGutuiEsp/lZj5bLWXvnmJxCS9HwgTMHFZx79OcmAvzmKQ5/Zg4pX0CP0//RC/xYDuvU
KY/2KZbksggyktKw7B0gLzSp0WmBHh/h+vrHS6nfnbKeoMWC2mbJSgOZXrqXE/iHlLdqJCOKcTKj
9sS4CS6JKeLEj2oGrDecPajzGlx4dQ+XT6+rydv4+NCnJ9nbvUqRt0qU+h9/lLwpOvhwYP9oYJu2
7LfpjEhaqnlmPrh1SrkeLlb8D+JKv9bt3mquwRq7Y5uHLFHE9DTnTLqxNe5UhJe0slkVkBfxq/a3
zU72szbiP2hnAE0Q9VenZp6En76BTdxdZHYIJQrQ2qWPZ8dKa5F2OIJfqQtdfKoLa6y6WXXPap2g
CMGYedP8VzAYpSkDyXqFQDPs2vDzWSFBec7NpLSwOQ4re8JucAwrSfMPKMZYQnWvzo2C8Mafr9k7
bHGQLhYRJrKLN2BA9aQHknJ6rVG869kbyTjyR3/LeT94c70PM3ZnqabVDUjHYvqEyozcZsGsqT1z
a3B8L2sf6I8unGbbb/r4o6s7a940SMgULZkNCebTQWZDKN0LOpvEJZhhacEfBImdx4u2rH3u5R7v
93E0dhFdeSODP03XfeS09+eh/YY7L0Sy3IhKMkWcRezkYmyOeC9rDAETtOlj73O4ITPYFE+Esseg
cYkHfzkNpa1Xb2oFwH6CWf7XJZ4MdHBc64GJi58JZAGmNO5S+t/CTbAnpzXkCQ4/RVfNt3M37kLe
hcir9MrHI5yDBAvJDizQ7bFAh8JAavD+PUoT9W/Crvb7YGhXEevv0Pf8xDBpuc0HNeD2K5QKlsHy
a0Y5levE9vHfz3KpOkgm8hQOfAvYaCmRBBcigaA1PLfp9SrIojRGUm496an0X1AadlFRe2/9DpMA
YGuBTlgoCVgXB2/5TtoR77viTjmz/9uFbVspoTbmQp41eCBNQ1t70KJcBY14JA+PfqAKypqPKOy9
hzeeiCGjJSA8Kz8CumHCy4SpF5EE/0rg4BZM9L4iYZ1l/TzpN4wpFQgMI8lIe2jqIVXe56LCUy5t
Tjx8r7XbRM/a/OPHQScv314Cem7F+r+dc3SjBTsy57vPI/ix55nN22NdTXRGV3jVwDNip8nM1NXW
a38sHXkHKTR+7qW9gttkxTIcOsGHmXQsb98ktFHNCHgE2mxgB7Ce9gapZYxoBe/0AOx3y9D07oOX
SSq/0kXtU3YmKebZtKiObanYygUYzJMZOaf6OACLEZiv63JpYU4Epp0zkuHNAXaqYaSp49IeKcmI
Qv5BsrrxKXq0SLlnc5QJ1Fy4aF9CGh8/NSBGaS8gOEKnlYHeH16lBalwWTSu7Mi0gN/eV2FW0/Xe
B/VbBz1KRfxwouqDlQ4kkuv1mEIoDbpyfRgTu/4hAgNEitloYMNi4mXBC3U9kEc84zV9UK9JveRP
9amI37XbMRIBAp7tn9j3T9xXUSo/mFweDvDfgwLLNGGzDbfWiCoy8ruJiXO770C/I2YjtD0RvN1q
FzCg76wmF1cS3fdPCiY4MQGBwqE25WbPFGAsMiD1gZkEk/CiWyFgjxhzzB/mehKO3BJlSoi2f/pU
I47PfTqVshCHVin6YWOfZNvzkTD4q4uSoz4TiIJr+TWMaZVfljjCSJC48qUiZnJ4X3MYghpah6fZ
WFOXBPEfl7kqVWwFBvH7bbKAOYsNupIdio/l6jIXa4yoXp685/Y9/NtyTdvC1u7NhhAQb1U91m5J
S24yzmX+8TlOwVDHhka+ktiSai15PLwRnKOPZTDkosUNN2IVvkFverMt8CDd5P1Cmi15UFjAZN7+
vaSh80AlPxAh+3P5LhxIaCQcc73ViOM6hkAzrXPkFhdMA/6iKeG0vJR2cB7yKa/TI49KWHUqnNik
AqjQxeqONW/kxK+tDGWkYsCce76FaBdaj6wX+H5BrY+Av4B/FvhesOLB6ghlqe3d8PKSiTdocblp
6VXhgTxlx64lZqDCdPyHaGEKgLZo8JBDtCFzsV1tnKxfmjrwCJvDggLBCljNeR9BszctymZGKW7z
4kfEZMWNnXyYdkfIdqYhHlkDj2fB0IsOB708Q2RdPeTlpmZgTS4PBi5okEh0hj7pkdrt5g5pLMGY
Lkl1Ylwdm8nusx0HqRV5aYHYsNASDaIbKnyxwKL2lFvma7Sme54TrwhEm4w+4P62Ba3y/ngEN2Fe
LtPclUyI5hsyKdwwiaUd7PEoKEiX4xYplla5mPGGe4NULuvW1CdHwDW5mzmO2NBhArmbg/irCfVO
bJR8rCYlj8WJFGY5LcIgRwcclTfvA1+hylqLv4JsWtUJ38Yl07kTkxgZ3ZiC/D703LqSnM6NvBkG
APJrVgJf0/T+VwrFFp6Opp7hK018P2OrA48/fCLr4g7zM0DgwcyIVUuJe8Be4pHb3Gb62M3o5qZe
wu+mmyMgyZdZDA1Sq+K2ipla7F0uHCYin0Kz3X5D5aiJ+nGGDdaK8aSsUwyVDysb0UxyAZ59Pxwm
YWpgjubmmnEaFDIbxMnAs0qgPpNeN5Rw+z3CDBD+rhyM7mgO5hOzHiPTSRMXHmIkWNQUQzPuG3PF
pjm+9e5BetxuxBH1GJFCfwUm08BYuJ+5KG13ya9FQUtOCZXqAn7gA8pMw1iOCY9zVnwDqJ4XGeeB
y+xdA1o23Kny3AbtrAq4+JnkMcfNciD2337avM+vgd6OqBA5EhUP06O8jdzofqUHPeASm0ldklIp
CCaT9J35QtHDZNqzga4RERTCHbhM/RgGf6bg8Hrd7uVG8m1lvgxBjget//+yu1ZqDTrXNlMij+m8
idaP2JRGlCztfzZO/v2sEdbnRy2LsoqVnhm7EfDaO+cwOkXy2j/LGbyrhml9HS6PiNwDW2rk7L0F
rk7Gg1rkQ9f9JpoU05PoqF12C8ta01ItOTOrosZPrO729mCeMpwNPJNesj/isJ9DO6R3mOTLaxpA
IHqrfKSm2tzrZGdjrT+V7HGigQYHp8pdNi/3CtJAOgjiSJqk3yEd2FpH8cmH/NEIYZp4EgB9vNo4
Ew+ORFg1F5wY/xfoHCfLHMDqGHiAhUVehSex0uHryDirj3itMQHT84Kf3nnc2+GPk0x7euvvYqTE
pU4DJMeH+cboH8GUk393PCi2ej0Bk43cx9SCy1VEiWAcDkSkpQQ0Yz99aAdezAv2OUV4qoXlHMR5
ffcJPK9xwer/zOzeA/43VnYLnAJT2i5eB7my2F4RcEKEY4w287+aQTwsl5GkwBilWuhyt2onDpPl
L5Hm8ItrteNJAIPJ2Nt/QR+vPxa9egV0t74zK8TyHhyf19pVm0q4teifSEvFLtBn7Wcy5fPp47rR
OvINLla0YSsKQsLpfjK4EKVo5gD1CI2ctclsexwwEWz6iCbirDLP6bbpttrILfcpf0fEdlzmJhY7
7qgYnhnNYwJVzD6X7G5rObvIQXTLq3uPdRlBWsq4/GoDm//4iThdnTNGyVXeLhHjZLzZYhYnrpsl
cSwct1Zw04BeORConoApkWgQx7rovm3Q7GZmSnUIthslMUZvetOPdysNwF0vgQJkiYxeYbsrPTN5
/GnrSXN8Y/h3PfY3UKd2r/Gnuc9b/V4hFni1g5KFesgRiiqmbqPGb3SRxneV064IyYDYYj030i3p
rdOqb/2U8qcYXmbNAcL59WMx1xlNFxfHnJcQi3Q4RtUx48uh8qNoStIzQUFADX6hrtUU03S9Og6h
I16T30Aw7zR7mVyL1m0Sowo7hGHOcrmMPI44ZF7zvxzeGpZWbJdicd0dXrRjd7iVJUzJViM5PCU9
ImzVknu6hqcRsMpVAWujZ//pAoIEkFbKURthGEKwJvScW1vK4TrTGCRXbwfR0KiB6JPF5o0zDQX+
ka0TN9nmlrUFbUY+cHcPBzDdPZA17eKeoRr9eHDkINOFmRTGXnTfxICGvi3/rTDal2pFd1BR9QKx
OuKkUU9tJw/vy/IceucmlEuvUj019eGrXvZiGJlRysz0hFlqm48KTlc63G/PirD8z6VbqoDahwjz
ll1g+XvY3H9x+WJ8pas+OUUrF6v2Nrroyek3mBx5fZXHCrMOLhBgJEBFs5P4oxCjTZYX1D/9an8J
z3VB1TCzzozy5raIj4gJxQ22soTke9e70OZqyeDk+PJTkZ37OKCSq8t+Kap0Z28kjt5rOFZbRXrZ
ZjszuGbpQj3I4oFX3ncMDa+xYyHsxJx7M64ZCMH/jGGDIm9C+Bm1pC6Co3DFyLRFAKUr32PYI3i3
cP7qGpjJdeDnGwl+Kx8Cva6oEY6nRN/N4no4vh7UbVBxOUWw7Ve30PGf5H/Mu1Tj6z/g7ne8hK3h
GKfOq0m+SPdcvXKZM6gtN/DtVvAxM084YfBbs9Rcmk8Zlj82f0DdhxpWuJLdXOP3543eHY7MUKnV
I1mk9OTSIKg/xt3VZSP5aqg8NLmXFtVuUAvzJzR7HZ44pucJJ8bmX6AnUm4Kp02zrY3R6179fic7
3dDooi6r0eqh0OIE2yBEeSNcRwDFHvkM/+7OLnqaF8Qne3zOWO+eXr9pqG+rgZ03IWbuCW3OxCdd
trdEoOjtzJP3A8k7ZV9s44bQRHVQIf8s50r9GR2HeLLcuUQgCuOCHSPgK/Nr0YhdAyrq2hBMcW7Q
dQ7jMxe3KjSU5snvAuECYqEOiUNRLpSKSqhbP4WDsDzqaqYDbrwqRvL9vEhdEO2LtkIRFes0PYni
LVLdK3CunXUAzX2RJpsS1Sq3MV+2mY6zTDuknEeHn8VVmzkPqiUQ79ropMgv/0f9+3e1hX6JyJYf
t1YesyqvAQuAiDJwSNPNf3VIcnKExYVFmbCcVWKZFVAewz0EkxdzbsMJK79BEXFbafO9N20/nu+4
VMBHwWF0UwwudcfJH69130uw7ffJMCJUrRKdU39C04q3YRbnp5Adi/frH64BXEdODpqbYDRcbNmW
pvcQ9vUxlej22IzrMuJsRRIdNQfg6km84zf6+NWEUS2nN1zh6wkH5P4V2BMUenvofUY5IhDZ+9Db
VZwqLUOKhAjt33+ndmbJLBPDpwnFwk0Pbbr/2udDIPR8h7QhP1227ZRHnoUp/MLnFHfpr9Ph7sIf
qbgMfIpUKpLEKfZMe7tTwJSSNZzYtMBFxq6sD/fqbejYylYrmf2knF2HyfzLVk1wlVX2nQTza+2C
7AK7Fb3SlecItpxEnb0VQOo7TLpRDSx9/1vg1xWO1trOzBLESP3jjwhOIpaBxPUVcfuiiBkLaMYL
aadgwXNfko18IiLcuyW+iY4sY1DLpSX9OubmzOR+u7w0J+ThQF/tI5t0hGLmpLnV+jYYfUnLg1or
/wGeatOv8jHniiWkbfevSMy+82ixSuGNuu9og8hGqsl+IBXgBIIZL5poiT/S2iZ9qs+Fk4qdhnye
wcjCvFQdgs5N5pw/6bzkegj9nQ3kgGVBxIRlefAenBESdAaKr4oRby8QOuKfpD9fVvOP4ePIwLm/
txT/Jv3XUUANrRLSMrt125325lQIq5xWkzKcabAt268EdTYJDeKx8z1Wbsmbu3iOKWzNxhRrvRJr
V9+BNrR6NL3/7Bqvkg0DovgrShf+rS3Y+CrLF+mlKdMR7bY29kEDfwikVEBlJgrLE8+qTccK72fu
bNU2xJ+MpZw0PUX1v88/okkPWVd5um/x0w8Hl4NZ5vl21fE3Inz3Ay4tC1sgm+AnY+l5VjcZlfru
9YSdItNF5roGCrQxt7pWApxCDNSYj3bjEjlOXG+0EdT7G7FEdaCgA0RT0H6SChREx4AKRjPk4/LU
PiMFnTp7xNbsaZ+82MOWzeVcHYFb9k5hHcMh/TNYRU1h+nnEk8UVef/vphxcPOMtrUPN+8TL6x+l
Ei46ZlF2EdyaCQ6sG0VaevRPGqaO5p731kSZEf/XHPJRKUPMsa/ida5fZKsuZ1ffwukjEKmC/YRu
yzda8IzVdQ6eUqKtnVnZS+/v1M68bMhN5qJ0JWxtdMoxnUp25m8LtpT5iUrXADq/76piBuRUY7l/
PMRys89lTUYbU2ddERH4pSzJ49WRv1vNiFjVZVg9EGWwcIzp2tBtZhgjzkjRPYC6IgYu30uD8pe4
ujmaS2P++iwwY78Mt1tHjwvebLkQMrAgEfDSrXBKRwJB8sopQ0gW+SLOaKc0DVBS2CysIq33h5Ee
7wuNKlQyasBut40yvUkigD42MLyJ1GF0OLt3oH7f5DzaZ2xwjgYs8WYZcDLZvzbCVp/MDIT+LC5/
WRDfambTZaeAPq+iI0P7lOoI/dEDycSSgwE9EMZkZBLslNl641OT/XiAVJi7psk4e+kNCMyGaubi
4TA0mOytVdzHwRQ4oSJ2hYhKTKwYomRueMN92/7zIuQiAwcX8TcxMzfKcvVW5b3jN52yeKju+Lw4
X25ERJL+Z1lTKuQqHCWQQu5V9tZAty14qRg/ee1TDnAXJPgH3dJXxxWPX8cEq8+2xjTkSbSOTaWs
4o5yKpBZvIUBMnYIj/HkGLQFQreQx5lI1z8Mw31INHgEFgqpSqjMzT3RjUb5IQc+MrNQvRAKL0V7
cAZuMUkn+ne41JTTEQdtDsOJOquppt3Srjs17WVQpl0nyjWLneWDlcbHDXwanWVvAsxS3fxBtZsI
RED0ZBGetF5z9J1H4wSzM+RDjOVlbPDKnnxcN1Rx0Bd15Mb1AUJBco7mrl+WU5o6oJWnKZ3egdzW
kykTgtymufr9zMtAAxA5w1XIPAsz5b2NLXi5Bt9N9cqYYY048MU0UEUJJKeq1VMnAbDTtDDDnErl
jDdeH42dCG9cJ9TfcqyYBE4KeXbc598XbKzqsl3m4qnCAVEkzPqRNEP9gO3hJk+0P3yHzWra3CTU
OcQ9vF+lieiVWtG6rQz1bEL/3WZKzp/pGAttjKhTwSSkiFSS0TDWu/YP2Dl/1O9PW1a2CQqMkoBX
ML6XogiTEmjTDqHRDrWDiVnguac4E89RguwPB9mXkFefEw6rPxp5fZJFP212eK5mLHi6Jm6lMIgH
V1s1y+W/UkYVua/LlmlvItUKjd1it/PCDg+opT8EIdQHLkPNPKbnPBE+IjDSlZ7zE43rBKG5HIPG
1sCC4Hx+f2SM3qLTIU29PMoAY1TQfiSNcoImtKycg0+vKctG7GsQOouogUFIcf58TFe1gazeVKdg
94OlGiAlVTaQ2rKdsrx1BDIQbvwh5KSKTG1cX3SL+oTrWuY50kbhzXcRCgAuGXBSOCD/miRrVRSm
8+bv8WoxwPLmJ7MlpeibW8+smDzgWdtgBbCkG2MoLFMuvLdhRizFc04WcdFP8DgxELzwwa0FwGC9
2GAQRwr3/4m+LEc2yFAr9n+x9bDveZR0EpUFw3W5h/+IAKm/N+WWcnUFHZpz+cFdxU8V9V8zzgtz
GGsxBbqXuXY1EycX01sWSYy6Z4qcd3O/VIeeASyvf6OdXOfatDVEQMCWbuhaQQiy9GpEkg03a4K+
caC335OLMYhZcIEim1DD3ohZ6UOHpXmqe6Lw54e5/o/sjWQiG7JbS5zO5ARdQwOxYpaodnEvVnZV
zjvKs5b12klzcUyM3x4E3hNRZk9bNACCMB3G46VSRnNx+2UhOqLjgYkMptBIfIlBwe8ZFKva+vB5
bBu7rrp9y+Omju3/rHdZ/WooPqLlVOg4/LriANObocC3wmJ8t5a2u3h2Xs5NUqB+WXmdUIdBSqxu
6zgGYaXt6Yd5WfJTZHhu1+ouXM2aJAKNRPZtf4O5W6Gk9tL1oIP8NaFXXBzxGHlqUF9NUDtLckmy
LsKqITOHaywKymhXt0kOBiP9OjyCpn946UFudUIUuFQadS30fw7QliyHA+mW6BHyIwWnrjpe3L4r
7LlpTz+7vjGMIon3EXcKmYGehAnsbHeJPk1Nzgqes23ZThi/DVuE98H8dll6y1j7wOUiycEyOJNo
hCIMWMLPnB0tPh2JO97+x6+LKKcL+xYEXj2PpFgHEEcgo0kelzHj6shJTxbcrX51iAtJ3KV5/RQG
gw5yUYoqiT9OzrEE99JIip4GZTq39Ni73ROb6B2pgChxMdknP6SYT6eYEdmTKChe2CH/wktcg+fR
UlABduPSm6irLDqwQlyjZYRTk4vI9CPfxbrrHG3My67O8CBk441fM/wWdvCWFo54vL+38MBy7JCW
qBPU2pQ4smjpsdv3k3AhD1kx5hv5YTsQC4ERokyvlRVcfy+oqpL7JcRwaSAOwIoP0zgnjz1IPFbm
VGv342UkVeQAhfU0j78nuHT8i1B/APAQrmLK75yjtvXLrvRqgmGByELvmoG//vCRyv1qa9gjZgx9
1fyLsqPqQLqJe7qBpA9L7iDIYuFFjP/VRT8Gb07utEaGBfBM08X5PW2ofdEFaYLM4Cfpf6MPRDWo
PpPB+T9InPZcl9cWT+zTjo7Tb7C+cYxhDLtHYWy6UKEO2cy8sE6ImnY8u1468llB7Cg19wK9Ifha
XHUCUN4DRC9/62O+O7OEjs1E6ibRIt795iq+bhFM16B1IbOlJWtTJRXbDu5eWq9uNXEUEVLZsf3b
mBgJhDzTy2U36MWZA1X0q46CB9a6m8+yc4Ls6erSlZdN0keCEEQ8Q5dCCFeTO788bvnFm31VeHz4
mlpXpIErCIANVRwHDCPCP2i4vmsK0s2Xst1UcKzCWlt8GMwUeqUp/YvfJ6QYKEXl9NlZci+jtiw+
phSNPpfF9cmYCC8T4q6EECxx9XXQdijfyrT7uXD8V3jExchfd7JuvqyKlmrOlb8xt+XmdgWjPQPg
3jLtYpL5H2lmw+0vYHPsTnd9mh5pE+7FNqUjV67OfjznlHUnkL7UFauU+6wSa8upWHUY4CH0yFUG
q/T/KC0d4teLO08R39DaFRM/65NwBU5w5iT8jc651y7JdhZiJkvx1shqklGzF5LjH9DBGICXJpQi
61nmAGTv0Pxo1mq2SPXxNvQ+wPIuKITEOU4WDgNWQOKsl8dmviaqbInhZ95qguAFMppvEpzXJ6pt
Xck2X+yF1NavP7eUariNTnPI/LWVD3upCFBdvbtsGIb+FPI2lLyfslDZOZLGl07jvZ/1jNia+coZ
x6I6yPbP9Z4wEn7INf39Il1n3/VEmZ69UI685cAN7lbZEV5jOQBgW6eM6IZiETwjMhqUy688fxFn
891wtjxiqF3kFVVyco1xvfuAWoN8Y1VrZh5Wqv2iYxaypxSHukjUN1qoix3dAi7Zt7FKgBtnGwwj
UphC7k5ZUsjsZTwl78BYzNA56I/k5Mly4mRz9uV/NHb5RXcKBnE2RUnEEHGzM1+J7ZOk9Zlltclc
Z51fEtVRl3OJtEfqW/Fvw08Du153YZKc7PFUitrM87bTNWcTU3Sr9QeLpuTsYvIlXgj2ht9S7Zvk
YcKHbUdcw2mAoOsN+K44mhiGnDcgFx3gBvrHSpPghVJD8+c4+0pFo4bibssLEfsKzSyniheTDC+O
hnXK9qo33SULwKrFcE/Ax2OUu5XaD0/n3zPSN+BFHuB19b5RK0GWQ5EF80vMv2w/nVEG165i6G4s
BVUAvnQbeJb0+AEXlus0nikUFCBGtG2Vjb89UQKCsmych7g0alytf38MJieSxbtVsNOIjItli8LV
AivYa2ukOa1x0UcqBwXhzytAv7MrpUFk1xwjlIqF4dwfw7Er55LMOtLbEVm2RoP4CRIzXPJ0qI/M
zVShPNGcWbYvOgRX0nr1NJ6+mAXGoDJ74epVVko9MNaOMT0AdrGug6clxWAxOD+g6UC3iTnZMFU1
zXf2cbBngxFrRSGsoTgQMOpuLajkZhLAZcIzTnI8e1hZDUS3QRIt1CFCRvobM5qMGrYbpInDirYP
zYkduJ4Wi5Vk1aQnsxxxQZytj3w5f0FSN31/3senAZF+FqcCIDjBS92DOPXTRLCVNepJRvw86CyU
xKa5ZhQHn6B/D/ylEwwoDR1yZUs3vxy12vcV7brSNssKKIq62e0VdpEY6sj552n3VEFRP/XMS5wO
cK3ed19UxcggBzRNo60bfh+LmNpwIll2evEJvoEM7v5Bj/697/dwKlEjq6PXrGfv0Sny44Oq9gsI
WAopbo58+36TnXcF5Db9iKOfWyHIE1pX8nz1OJC8R118xA4QbeyXZ/GVbW3VHhhCJv5ZexBBmiFS
vq88eF99u9VZV7TbpR+PatI88Tg5xYwPvwNr9SVqhEkpmk/kxcOZ7BbBqZdSu96gnE5Jzy821fw9
+NBta7NR3bupDmPHikSDoODiVV9mAmxx4w86XZOOMJB34N0gqte9SH1WKLhaBhMbnmADpIR4/dph
N4RujjNgurKikN3ZTxYbAOAvSsq7u+dTeDGkWKHj9sM8DjikSFnznTCNWA8S76g8ajUjKIhEnH0E
ARuuYTC2uMTqvpn+UVVgLkc2iCIt/s6aH73jkGcnasRYFx0J9d8B03/qvSgK2wKM2MG5aorkXhxP
BLuSnDgMFLdz6lP8MAka0d5pvJDabVtugH9hxeDcvTIFxeHW3aomXiSdLxcQqba2XipV3oiNpHyF
+r5mSA/7iEzEA1wqhsZH8OZsYspAml/N3dzJpHhbssoUuKbNQrO4zuYC4pBhjmEN+5rKo4lH+FPf
garRKM/e4+94YbHPvWi6QHkywdDjx6NJ45anJlhnZz7IkgMOjh6wU6dG3V0obxOP3A88Wd+KrvA9
WoCQUxPlpOK+svl1TJoLdGw4F2g/1zUQnIgFnrY18i8LaENvS+SN6KDkgjvTCLtLXzxaRKf03kzO
t6J4IqvjyErcOXWqlvdAE4aaZibEa0zt/Cc+r1BKRoU+9UNwfEv/guhU8FMX8CqjNCMQVuzvJffF
I+JeA2qn+DRF7XIqEVKP0rtaVv8aBt95fVI0fZuLH4Bdkh5u51W99oZMJpwo9WY4wCwj30bG4gmw
1Jq1o7d2+n1sATbNhe6LcCOnGphFxrXwXkGJW0JCj+2LVgOjJc8WxRVrahYC5t2uBC56stCgPra3
f4Vi4LcDeG7dlKAORCwq90/Il8/euvreRWzjBRvXnGKo2axD43mGEYmsc4RtuuAZ1y6Ijez6BrXE
Nx2K9BLZnc4UzbXG7kDgbFLBgm2szewEsHthkQ7ZU+u5P+PBRuUPJeX4+Q3kfeYDDXD4kEehKySw
pWuw+Yr4rRuevPjVLNwo2b0PzG2DJbxXFYJEIbz6qi3/WXLhNhCC2WXj0q3/CyjgaPBDfl8CYm/f
YXjpNIdYbN5ENyxZAeoczX41VCgjEZz6Mq1bPDD2gyrRY+nwZq2nFQXXtKdYTc7BDpFoUO31FuAj
0FmquGRpqGT9JyHvwTVTBbWvCNQ8JH34evle9S5MrieBJWFOvBrTjjEcACss/lJS6sJPa46jbiKO
aQq5Yg6QtGgbZu+hxRD1xqmmEN1lcXKEXsnHgyijo1gAYXBoeS9rOO7Oz3zTGdrAwAk5p1P66v9R
j3IY1ATeEuy8iwYbeZgjVPBlEnussgsH1pujyC8C4pUAMyVNFUHP8T8WAkzrorDoF9GPPxlqDkhl
BON/Ny8z5RBTwoEc/e/J/KZQDuebOlEMVONQOQdWHICifBjAQJ545Uc8KcmdvtaWPw5ktEQImt/D
j1oHwK3R0JlfatL6D25PArovoPbntGDgYy1zSZrOl/T0tdlsULK5MzXhctJEMSsX1q4s+0ELZ9PJ
oJxTlxYxe6t09b1duiZH4/jZJnIJt61OS3Sn0NDQrwyBAa1lAJc9dcjExuqIConQler8RjyULFia
J/Pykx6lgyZOnc8rURgdEsqvc53xOPBHdJ6FSQubolXjRtSQXMbXB3Bz/6VHtlQPSzeIs9Af69t2
exnD+NuhdMdCNR+WlPcQLm5/CUHetQwTs575uPZ4lBuH7UUzqtOvMRwMBWUrMWgA0jyzW0LsXcj2
8y/OQLHH8acg/FkEzZc7UCTKtMYyDew/q721apOuru/QmzR197TYYndim2rqz5TznPvFytcuNWlG
lIob1dZezy0GnowD+l1uziBPdWDGUtpo2H8XVx2efDhi8r2JynmwnTMDLhN1v3mDKuF4+PJUE+br
TTD3D4PeocqQXF/rmfvu4aP96fBP/QSSuWiDBJzLerrMZusyq9yn08S1fMj6yMSfM0pChnHaYmMR
Eq9lKVe+CASJ9NFQc8rwNmK1n/OmavhiawNiyl3Iblg5idl7VTl7TOqOcp451VgP6OF6M2OiTcAY
7H2u+aFxZPwLK1vk6SYtSTEgpBfV1gvs6d64i1UNOxgkIpFOWGhq7Sza9HxglrNhOnhyz333bxFi
yeUQUv9S+QDkbMxNTnmcOBQq0BXNxoKBHfJjxcHYbcST3maUzNbwq6LXQl+gLmGh3CdmtzI9+wAi
uPdOPZyqbVaaK2q5aQHJgdUFAYm0axbamYcjN6Kq3O3VJXCHmAPehvszFXVcC6yo5mFs/4gOY5vn
OpRTy+CbMxXWQ9Z5/3QU/lLjE5bfiY7tskcQxHb3qLh+wRafZUxa9DszGOw7xPxfdt3+d8039ENu
PaGU5zB2/fDXliC9lemXJcUF5pUIgb66xwIx14KeH+KxgOSwAz/b5c3Xq31eiMO4waXJ/X/Ji4Oh
F3hb6DUxSSPHjga3rvhDNJtYY0ghIMzfUqEYBCJY9Ma7dwslMIVdvP5qc7MG4ZjEH4k/ELkMHQgH
cpqqhEL5rQVfEz8Xn+YVSYJs/WTzkR3S8VAYAedeAz0wceUxinVrbbYA+TgndHj/hR84xmlb00IY
wvdnt7/EmWxYp17tNHmI4QS0CUx9dF4QxyAteh7FVIYndWextLQ9Tq039FiEMkRXdOhetBEcm4tx
QlYYkSLsAB++A07HhXZr9X2NfHREZ24enz/shn6PayVYIAIXZ1UoMdTbCjTW1aHLTKE9/3XcCkDs
ZWZRobJdiEg4TqzG1Xmt2YvLVkUBvqP+sqFhaiIMgm3/tEvL8FoEPElYm2UVg7Al/u2FzcWRqcrL
DXu4ge4w8FjflaeuHH5LG2s5pRX7tSTGSyihO0WISuVz6DebKp+xf0j0Vci3zHbzL8raxydvg8tb
/N01YbenbI86IRVsfbHLVCOYA6irN4qQuihrPSNf5692latbE7VkAExtCG8BHAUjyjXvy0ESfZec
jwm2WXX98GLgkY0PnQxYchij/IKBUYoZs7LuLkSrAoIoRLfam/FhCvdF3m8AWoVglPzKFE+XmYUf
+iP3tAIo1ot4sjlL13FTsRC84aDWvEx5OU8IYHdrmNde7tC1QpAdJbtOfSEti/aZKStlCqGvxzQL
YzfkgOJh2fI4fa7dvB5kvtzSPPJvvdSSak3tiYkrABjcXnnYgu9y8EpoagA05nuvJy/OzEw7ydrB
8sTxbF4AkdVoHgsozIahfbx7oOSq0vWIY2uWwMKHdJ5ZczysJtka8nD3aOu5sLbwkhd1HC4xYiC1
U/i27R5XlaXcpuMmJbVGZKLbH33vPITbLzrm7vKh8J9wi/U39JHh3v6COBL5f259u02m8QwX+MMt
x4mFPC5K+YERsI3TFE3sOb5DLd21j2EnqiFFx8kxYqc/LII3T1fEQ7galP/obQZgX3PLiHY/PnaZ
Fq6NPxs1Wogg2jUgnJrhnXPwhH8Xlc5GDkKJNuMAqi3P2cNzU4VyJUShpZdD8b4LPxbnj5naCtrY
I1/C011/yVedLxVLGHgUQS40QkykUboC1fZTB9oVBAdMpdog/i7hGGwI9+aTS7ddKM1rLX/U/LE/
5ntTkGIUcsD0orLUtMdOhfaYIlxBWe7HkdGtFvJc1NbJwjeu/q2jJ1mqULNG7tbfTgl/UgeK/s3l
YaAYN1CJNVy7Gon4OoJppaI5O0mjehyTOl80pfEhEKfEGiLd+WOO0Q/sqku1+I0nPw3rIwBhSeKY
bMYAlnjO2XfjAFIK546djaoph3IyFyPZDeKA/TEk00N5uNzGI3kbPrDe+2Y/twB22mF6D79rU8Pp
CFGVeDwfY1t+QVCD/h+gdKlZ5P0QKaEO3m/ULcIUZK6Ujqp5hu5kRE4/XW8FNolpkOxsbRBdpybe
CrOTLktMAJ8vaOGIiZJ4dDbnodhJIJcd9aVKpb3pAeIRLCw07xOmbqjkaHy6kNqA4I6B4OsXTYkb
uTw4MSkkBAYfzI8dlYf3zDQ2djPu6LhEdwNLfcaHEkb/3wjnKTGQEeJnbMvg4RUhbdGSTZ4iABcG
wtxDpqAJ3y9ySf/pIXsgIClTR2YDCz70ppCf9gssn4xYlx0uC8a30GI8RgHhRjI3gfx3/27mTjZi
eNAkYHvRBVQCgjUGbbmKihYT741zads/5Ocw9f7E8rKoW/6l6VXaG33Zd4hatAbDw9k3Epd1sI4T
lCBX0+RICL7+tBAEgFaGXVYz+Ll0/L/GJi/HkacNB+BFPb1F/aYcpe5bKqM4t2guNAYloa8Qlg2h
mFSf9gzYfwTh53NNANFGjyvQAXTVyoDUT4XJyZGs2d/KLD1Fm6f3TAkUc3jmvTHJApGuF8buYinc
bV1R9kZPiAQME1W2fhpjySZvfEjEcwlIvN8QLgKpv2+QgmFEo06x13Zj1Sglhg1ro8Flw8xvgMR0
qVsJJXDvnBqODMcXf4TXjpAKPr7cyd9EB5/r7tAmiRuCVk5rqK5vG81U0nt5vrwcLx5hN6RSXO3z
XR5mBfIK9uDoc+zGHd5lUMN1wiF2ziH85VHJanXo/JCoN46+iPYoXc6MCY0TFXrHeJ5P4QqAxav/
FXggUgJHPu6CF3qg3+l791BfBRSc1F01n1LR5pENU8vKzpQiBO9zcCYCOoYSQx0LGz1s8KISssxm
2pY/OTf2h0bQeLsJY7fve0fYvqXYLR2yXkQJswr16B+Y+3RIk0WaVNwMQzRZJ2E8dKJnuZ1bg/4j
aKAehfDsfglfB9oOkSQV2EPUegvkwWMcZsLpKZsnAeW0611bjSEQaDiZXrkpha0JrfDRJf7akoR2
goIuqHkss7r9lKo1z1xtDvppkKINq5xAstbv6BJVCGhLWr9Boz5OSoWq4XQ6sp/PCRv8JdcLM7w3
/mmeapl5P77qO9fSCmF17zsOkGKioyprqamgexT+1gHJ5mmXLSETDSdzS5zhCjk7t2+zzfTxVNGf
LztwwcGNWOWzJMNmgrrp9A8fTmlh8AIuZSXJmqUE3CZpgqT8wDYv5urEcvLU+9k7ypDGxALF/Tm4
V43VHtJDZStJnyGOlDLTUYv99iau/IyqXkFNzM6YjJHkX2oBIDLSmo7wI5303qEi269h9vBjLPMt
vfG79asSGzui8aNOrK9GblhMlOKwV7z2YkPVdgTK0KteLBNtjO9D+w0hBPfFbLxjihomeobtmRzJ
hWvZfiVLJ0ukRQfatG7yoSi2H+JZDvAv4wtWBr4zQD8SALhGa6i/GMHybUXxaJo8LgODhtklv6Li
OSR0bMqRw/P+rQC3XQxhKXJ//B7DfNiR2CF7aOtFJ0qUUuZP6ydKrWvWL87B+lYKA3q/Xq64jyjO
pZf6XIZt39o5YeSS86FuzGVMr7eylEEGeGKLJ96W2hu6cxO6+xgOrUh9z8Fo8xrlyLSlDwlqhx8P
wEAvFWTeEAzqJuu5Yh3JrnwRkohRDKG7kUL9AvK7m271Zuydr6/v7I2WTxDc03cDZ5ti3GrFjsvb
WWu/GYImzPm8sHTTAloEMMqYqfXPZd6o1lO2L2rFUzDQVTDwCIA0rsGa9a6ZQyYBreI/zRnbvEo4
4s1TO+Qzphy4IQBuj8tPmb8M9Kep4hCWnK6aHBb2epc3uOYZxLDI/E1W6vhjNI1prkBlMfRtRMws
PK/2dCjI7gH4NLKVw+G/ZitdgHlv7x+IByBfY2HmkVhd6KagPc+k2CLPFiUQ4OAO10RL/wOr9a5W
9MJ4reATfssy5de/02NxvIIw2c3WlH4wt6Mz5cC5lq+Py3My24dY4CmnPEbxtUTBirD9ea0ypJoC
1mbb194KzizB08viN88Dt3CML5ewivgZ8OLzdV7Vm56v4cGyvkTM0yN17q3Jp9v/38GociKtNgbS
G5Fmzlm2EGUh/crpFbfG8tPFqsOxw3bkRd3uRz5hSyazbzU59a+5eGv2ahIYzm7r0W4HR4vITAsb
zman8NAQ9e1P5cxi/zrfsvmEH0T/Iw+N1CqBAG7Rx/jImUlBaX0KpsrSCCVXjKxhlJySlg/zXfaF
ED6IwVMSbwRjE3hCFPSOwsQi8PCM8ka+rprZUDpyTt9lELmydlqc0hdlVQBj7drt26AOs7YnzIOs
6kUAxTBOTLq2KcWUJmgTW4eWNJEYIKZKj6nIMNsC+E99xmOafZeD6HgDAJlQ95798vtVaz54/lpx
wiuFIVc3Q6rMkxYtOmTiPVqnBKL/3kbi2jvE94C3iwnp4Kstqmwg2H7f1oSwdZQVYm9EUtvSKKTR
MHKk7SjBMtvCr+u3Cyo/r1KfFcMNCrvTUCeTgs8ipvcHyDPyvz4ZCIXNXm2bqNjEV7DkY3V3Y8D4
1MhCkixXih1PgxLk5ok1jLVGDX5lOPxrxBgG3EyC6R1h2LLZIAZdyDwiDHgqwBGBL/ibr8cz58Bt
cDyCY//fTtk4+29FUWcBe6eaSvi3iYsokbx9KoLD/7kmlEDGW2EZreKhLRgjLkapgsilq3ZKNh7S
bCKQKpQ0wcWqGXmSHUEFhkQtM9aAq4XgUT0wZktJk9qraR7iDzGjEORoJq+Fhi6ia1ohlOd+7x6O
mcnN/vz6clmDZWzNF6UtkZxpGxJ9fOv8DL/d+PQmSSLN3oCafLRhYO5ijlawlaI5n3gAWvNRdbdk
xzzNWCEOdOVMFW5kiGTRnIng0m2IVkLiTYHk67A7EfWG9riC46tm5A2qOgV363g/yD+qZ0BPCCwx
TY/g26aDGgcMoNLil2Vgda6LfIGvTIK1nYCmlkvrgFe/seTiB0Q8QbSxsrD3xEigzHqqV5wcjNCv
vPY1HzEoNHQUZT2uk5BHBZ/1OIgKGFKCyc1zes04MmIXCLxM0wzrybez0LPercK7GHdlrWOmSc4y
8P1c61HrOsIWFRepiJBhGwDUlWxIWn0rwBK+IFyokE8epmDw7nl3O7rdPuMeo7dEm38BfAF7DlLb
wWkUEkdx6TtuKxlz4xcKZCfpwTPJGYkU6SOEkELWLvC7OhE2g06jBoh5jL3e1yc6AsHb8vnhQm9N
8UnbBvc8xQAwbJ8/Iv6YfaWSh8XiZGcO1/Hx/V32uirKzEXmF7G4RK/jvjwx/moW5XbVeo9kKYYs
Dw5KvqliOxIhZ/acgl/ILDT86Pf6koAebhR6iylO9jDhuMSe2Cuzs/riE3SdLqEK3XGWwZnBCxO+
mjfjnGqcfd0SgfELtYh5k3Sl1+VOHUbCAegK3tIW+BYZKlVPeIWUGE5Ociy6DclsZTp+gNVW4j5M
Br706zFN54BkcxpzcGSXRDHwTV8/WTMQ0KNrU69vysEZ4BdR6PfcNDIsGD/iHOJ5NPYYxl0qgBJ4
PmcOjxEYACkF7vsvNo4XX9sFzvUckh2jSUQ9Su8N3q7mpwxboVBNB6PABjV8IX/u1x6pjSdpopx7
nhSkWTo4OWr+/XdWwqPeJX7xQmJNHPcDkj37gZO9zsYL1hC99wkIe2mi+45hz7zmBMa25POulXj8
gwIG8WxJ7RYitZ+rAKUxqRQgKXMksqCpqcYgv4tfdmrfB5kzJmQ/WEkposGH0kCOoYhuhJc1Trmr
50UgVpJYcLtN94I3VXLyZQgpcrneKb0T1CcULwhDBMtE1oEDSgENsywb2B9K6M3jJ037xx17jfrE
BbTH3lhd0cdtvAvh3U30RC6+HjGM3Z8oDWsqZE532pScEnsGjIwUQjjbzACM9s0CUWDVzNc+pxf3
q66QrFCf5tyVM4ZuIZrDbi9eYSy1n5e5zGa1q4jTYlBXoYzTwSAMbPGJAmD/q+mc45U36aougcDC
CKf3HPc3EBRsmjI2yhmXRB9M+7DXbtXZf3i3b+K4ITWLyUQpZcBxsyNHnTcBL24025pHzvfi30Nw
pFToUETUpcs6ck1QEl2YDQ3x5zDcXWRoJM4lvcEtO/ZNRDLepYoe1ElqkXE+RfwjE/rcA+B774W3
m9F+8IHqDU85tMopV7y9CKN8f3kIP4jR/aqAq5mUHMhBaPIf/6Pr1WNxhobnxCqii+BuQ7EZ/vA1
gzzlEpXJ3+6rraIsvyMtTzHyZ2gDxpa9W8sHcFkYn3DaRjsjOVPIR3FS0+ekV38aU2w7XSl8G9sR
1K437WXX4pP2Nk5ouVAbhl3Wc7D2nFAkjuOtcx2B7IdmKeTxzDLNv7aKQvtB51mxR626GZyp1+Q2
tUsZR4BdxLJBHhTeuu6MUzlEJvZvffb4bhrKkzTscO1lIEPV0S10HYP0ZQy5L4O2E1prwRq41ZqT
XapSCzFcRnWtJRrUS/x1qROlbYJ05L0x7S7MlkEKN2enHaI49qdu5kNi1EXY4LjmYckLFoF7TJcS
420RTubwtK6ern6+89hwwiVbr2GqZqDMzIVwa/YFTsvlrNpZ60lp61rj5DuPd3V/2lrw/a6QzelU
eN/8RDIbtfBiayIE3iXPq/t1SoeaBRNIEqNpLnKgjtNqIcpbh6CbkJNb8wDboN+TZkvwjmsxmBpl
htP9/dXZT3m9Z1r7WrNOl1C8TBMGtM6NuBKhcHAX7n/vrfnteANfCxlZDZuxEV/5QdoB3FUH98Ux
n2bC+AfcdL7X0xtiArHLTwcPDl7/S4hfRMHYHheUR0j+nzMi+kf9JwZhesSFK6PW4hNl6zLVI4G3
P3bNXw8mxjGkbVLn2UNCU2M1XnkVf00jmo1ka5CMGv49iH5gZY3AqOeFyb7EYnSqZNyraY8vPjul
nBMPRJzaxK+MpShAwEiSzF17UBtG3bEvzcX4mi4jwo9KMs4ygYo0aladbFkz2x2EDGOJIzwj4bX2
InQkN8KH83HsbX4fdHAi23eP0PX/PWQi4wqpah9+8D+cOXxd8fBZ8fATZ2v2YS6jXRrYTKRg5tdl
ijyO3qb2smpWumCm7rMeA1pJlJYrJf20QYeqe6VLuet7F1og9v8hkH6xuuBcHnEORxF0wb9t82cl
UK6+t+QN1fpULxvn0QEeByy+zpKMSpKVILDX4wU27F9AXuxBD/exPNH9PKh20dBX3IM85SNqWRZ+
ux3N1c/JwtqTzqpBBLDskCTgdDZfCgZGwpYTGG40g+Gr/SQObpZFI9OLnUapymP0/lRKEmjdsjqI
pTb96mA+X8aZkvUMsVTp3dmWICi2yuVphPmdHwOumWMmPzMOjqBKDay724lDnDnoNAUQU6e74V1f
wOEnS47w4RG+bt1I7v8Is4skXlAWOGBLu+iV95FSmmLrcyU5r7Ev+1xKSdkBeT8wR+pidobXClAQ
xPENsSouqXIL3NTX7/+UUWBlaFLRRYBM59hU8MS4jT6T6mH5wE6JLxThoq2C/gUkcrUHzQbOoJQC
PIx2QO2Mnzvd5P3ym9E8XXYdfBrORan+uvfvlzBtbcfSqZqLuY/1nEAQLlF4nN+/kysBqnp5PtN2
ZDTuGDe85lNMyrYJE82LFjVA9z/g4RTRw5WHH1a0UxNNlo+tJFkYajYLRU3jza0W1lKRPO+qj9RU
NqHaVYVe9GtObhdO4+E9WJx5mPT2hb6hsJJ5BGIMwsTq/kXArHI/e4hAU0JTjSnLk69vhqaAFobf
sjxGf7Ah5MOvXQHBsCCIvMTV7bFVbKIodBL/x5ke9eOCgbsajjUWNf2mmx4QEHhmVnseLJqy6+Nb
ISK3Xj0m/GM6E9ZH2NI56elDik4SPSE4CXnDApGFkncXlAlBPpSWmgxhf4mcGzIjr6UMlJPfE+EN
iQuitni3hdqdTexsi3+OSTGJ0rM4o2idavsqttFH25cbL2f62F71d9OMVM6T8JcbcRu/dGVy7Gpn
Dt3pw+4Ri3e9x7oG2MO1KH6RQCKEKwTXAKI5lVi/yvkru90jgqeTdEh4hOTzwbqTiBw6Kq+hiMSW
5mezrTdoR8TwOaNuERvGzt2UyAFJlF4c7v6SmMn29jH1uCsKqFjYzhJunez5UElStkm0g442MQ1T
uAiqp41KgF8pb6+NDN4RrjH/1Xcet3Okvk08Ncr0b+bF8Z8jJf92LfsHFsb70zJ8Tk7QfNBgYAsP
OFDhEsFDZ5O16WJC/h3+uX53Czx6mdxDEZ4zLyCPEbtyDe2JFbtl/X7Z7OoiXJMtGu9iSobuugZb
EQHIeouusaOmUtwfWZQW+DBA+QCsQvpEpNZNUJ54TrmwrGTegFOoPdjLXFttp3waJuq3NExKr8Rv
8gbFb0bY4SsCwuXOWQy+f5ACPHWH583WAgRbg8qQHwuS24dDhMwWUIc+AU/NuY96jljj9MXOyHj2
mRDF4Dccm29wxBQzk6pgjTU7mqD1u0iMYnl7fHJbkt49bOvwmNKtDF4cPHEJ7Dl99lLaqIJORzFM
XRaRPm3B5iu4FEqclRieclN9hVnmeSE/oDzo6xmVDGECoMQXs1llQICQqfYtn6X+uDeqeQ8XEf4a
OPorR55Q/mq4DMp3mPWzlq8v+bHXV04R3F4mr6e6wta8QdtzrshLQZuLm7SlmOe7LGEN+u6IK1hD
xSl7lh+jPLM666e0P3HCv8IRPIQGm2AZyukN4+kB0uqG1TkPF/tK5iSqalAe8s/oKyXYIP9vOLcF
j8pLAAt/kyDkOukrV2HqM+3IgS8/7Ae5DHeiW4hLj4/4tshoirxlqt2nIz5oLEhYJpybXnYqAyDC
5BDNnGlcB5wH6t6Re6VorxggGbre5O2vBhYiKsM9aCekOaj7eXEmjU1YDZhhOd2II+dNJ4EABim9
4pmAPmP18JT9wpVGhyRJKJC1eOAi9sSMqmanOhdmwxCFNcguidTam54jAbigT2bdDv+v3x+7cAgb
w7pdX47Kp317dVJfadi48loNdnRMVAjqPOEsumLSecqGmpU5sqEjKt6Y5x4WrK157J3Gr/fTfZa5
LfGJCxQFZNLP1ktYlTbM9Y3F1jdjauN5eW0b3xTd2Ml+UKY+9qpT1Twy2Aw0YDrgcFpAnVzXpE7Y
KiGoDroHuQZC5GdcE60e6YKPbFdjgD5KAKRDiDku+Ku9E7soJXTwofoftTLbYetk8XwugkT+bYKX
ZGZY8yCzwVLfNHzRYK5bKLJgBbURDXVS44tkgndg9RRiQklQ5lChQocV51pawJJf+a7ypAnz6PC3
NRuBFBe8YB9YqnIUaWANWzFtIBl7ofVR6SNMs8WembWZ2yTDpMptwwIPMAUEosdNazdfnsYxn2yl
hhpopsXtn10Wa8AYzXWNG1xdK7GSWinhiAeDcdU3fxsYL3pkFTU+7y5BSa/0GUx1skzJz0i3SC3S
oG9eD/8f7CJIqR/xrvE5r9CMPpf7E0N9X6XqrOwuoH4dCxnogPXhtwENH3M66cH0YdupUpWhboKY
AY5u4bTtNgFV1aIu3R11161IICucNk7EJrg2iSx595lFowXYxZHfn3LRip5FBPv+6JBz/nVxYRDA
LCR3gQl9AnLj0r33haMr2gw4FvhGslYFAuCAmpQZ+a+37pKDeFtLIc+qRvbuHKZUmmIGOs/AFtXk
J6N3vMEtQCNK1KRPqBN295/Uah0qR8wWjE18BJa8NC/Vh4fP56YB+fRKbemZKDMo1a/UUO5vOvaC
kOjTV10Lk1aq84DJ+bn0iAGh7vaRW3EY86fQIK4NDsEezbRhI4OZLvYFmzgVYqZQ1pYhLS5h1UBN
NXb+WNoaM1gik+9KCYccW6Z4EGI357aBs8omkWLFB2FbxVvOMEDd3aCqiAydTb0hM7Jr5Iavijug
kAetzQasZQG94uPsfAzsytkDJB+mIPqzCZXXxzmiWWmNS26r/QHOMyNPGu2Q2Q2Cat2VbjKgiKDr
WFWfQQL+azm7Kv1UMGb+9OuN7SRUhcrYMeFJl1eVpsBSFt6NDAQB5fljXbEm9dbtydXhzP/Ci6M8
pthxGTkloCYhyUv3tnw7OEqYoCHFieZhQMnAt3VRKFye2/zW8ltNzpamPH1GRpoRbKMdZIlT9wOG
OBAenaN28fZZAkX1TujXbApFweJ2pQgc16xOxgVgB/jJijLwaBU1wLIc2jFF44LlNqZY++VcPEpM
cjNwwainzGYZ7NoIs0qsJngloJo+EHE1jU4dK1nZ2S+ixb0lxI+VtzWc/VwReqiIdLujQKHmolu5
bVnqsDVmZ0G7PdCd0FEiCK173ugCAoJOOVKtQNkbVRcUHOhXULL2h1ouJ8E+W6hRIyuWtQTl9DQO
+IxWpoXYqS8RCa4B+HDIVnGLaz0tso0ooqFjyVAlAL9lpElbZ4ZGo4r1dVJafvKxxPNk8Hrzt4kx
pRi4RylVtVmTbxhCkRgtIxDiDhmeq8CqrzVQirzZCcMQccVbM6eeS186e5bEaipY9QhsTW3mU2Yf
5yUzlK+Z+dzIoTIlJGiKG/W9/A3wGlV4dgttphV0m3qqBHn1y7QfemWNqXM1gUZzxMCIS7ws4+Vx
BD4230l84GNklNigr06jmYoq+gmIilh3eS0Zz6AswPfIv8qiYX3ml1CK4XO/9yR+WrmHrxClvzhR
GfH9hddjzYsN1QHi18LiCS0IxMNiib6Jsd0/EMF0qIblc+pfIt9xFpYrLm235C9Bpv/TwYR91Ng6
LQQ7uPY487xOJ6RpA/9CJ0IpxRqN3fM1Qq5yE1SMpYuEOoDaJ02Yr4HdVifNFgFK3bvf02hFwd/i
/EjZIOc1hKpEQV/obas18e3g3boupLJ53QPkExRXDq4PPoltmWKFDH7/9Yde+SSGTTddxWOHqzsr
SG3YMbn9eDTtxut4EbwOlbTY5nYBW3KpWFSTw3HKMMwgtYJA5bwAmTnAIlTvzRJNSf2wO/23PiVT
gexAwWf2da4H4il+P2/0woqM66vZomwm7tZMzxfQwyhaTCaEHA+nmzXhi8kKcus4wpbXHCOqZS0J
o5EvkbkBj9iHM042jexde4eZ6wBEL2mB6eJJdu5uqorKczmWKArdzcQICzq5O/+h0UrMGZCbh14A
KZNyvwrYvD4ZUKYpZYxEqC3aaTaARNMp55FWDqcVlO//X2TgPpSFn9qhvJL+80t2NXIMhXKOaVpE
47NQWdiZ0i/6m5/hhId6j9D52fEceRFmM96OLRq7ZSNxB3vHyNcgdnAM56xLsciwCNFShH6mJlvi
B2rhkLQknHr/lZPhHYL7ojTPsYPiwQSLyBZs2/dtrFHru3hwVpGtVw0d7eyTSIOgN45FJtgWlu9s
G/6rtoF/l0AqVbygftz42lRzZ9IZDAdc9S8VWy9kbmmXVjZV8vXeln6ARqMjWZcSR9N0bYcDEjzG
Qk0fAJItVbSir3peK5bGa2LEHUPt7DOjys5rBxQtzw40Q5hTYHYxqJalsPdt310LyrcpP2ipPbqA
e//zeapK+ZyPNTgLhQtAkEzqihNNIc3/AL9YpaIZ2TzgdM7/1/NTuNE6rANPKTxlQwA6AbS+jru6
1orOWPU+geFNK+DVB5qFx0zjz+zvM/BjF/GIL3O4vJOyq9U+/D2WYmJr0AAGZbIg7rqk/8rPlAgR
9lo38KFacf80Jmjk2J4XLuG4PTP1GQx/DlclcmZv7B5bVqLgquOPvFaNSgJwJWHSzMkzUrQYKn1G
7gD93rR+N15ERuh7AMKg2blm11FOWDnwEft87ylHFuWhizhO7MyHPlFqqm0lXXL5ScyfwiS2O4ky
/KXoF8gHsgd2Odd31+GQaz0sVMvW+JodmhlpCmcoBiQHTxPxwBH0U38Qp0DOdR0EpzBRZZfUiWIW
xjr8ctwjAyZB9QbvLsRyn/fRuNC9j0Lr8qlyb0Y+7edtwZ2iaQdBvQXTylMa/o3M6qMIyI4yMaQ9
miG4RCJ/ZId4q3+kVA5FcH0KUYrEFaR5vCo+7TsHzW8Ln21S+N+v6VcV9/DCBuBs1oig/mdiejz8
bsxLeNjmv67UA82df05JJ5DenoIbiMCXSSz4Nk4fBylWx0R361tdh0RoziwUSVCG+qDuij/6eVEN
CDTmQ4TjXfTCPbjGnfJSxDdvdRBQ0yIHKuQdRud/tzW0N6/ptKASB/Sw0Tcn2W6l4hn6okssDlr4
h8ZB87ivp3utFiNpnnVKZ9KMLWyu6+jDY2V6v+Wb+f2JhFpKDjGD2mug2BzT++J3N0aift2/9ivB
PDyPMwkggC44m6NInOZQswOCFFrM/sZCNKFUBSCQIM0Xd5eR2av3N9oMABaSOocWhqZCe9VrOGHR
Y/8ntgQJ8lH0WAR85p6VnddBUDbQL4cDGv5mHZuVVKBA7VYjaOA/X+H4fd3FPli8VbpNVd3WImJY
1lXbkSGrnDMW3BPq073EA8hy1+DF6YhuzYCnt45Vck6NCTx/qLrKgRy51ZqPFq2a6Ag28Cz70hLC
zHWCQee5KA2y17FgjSxyueuzEkAPcKO/f2hXiwgyoXJvknVPO4/9093q2htKzegaGCZC0qJayhYk
Y9bHTjEDszSb3tKNtXdrR6DRgv1MWBI2YqLtBRiYJkUYPCQuzvzcM2PQTgExCJhmjEtlGjoKpZpa
78o74K2V4P/VumeKLPiAkfhhOfdH/BFxM0ZPcBxjrbwbeRR1CjvYbcl5S+vPiXeZLoubTnKBDliZ
4CpCnkXJoaDJq+A6ozm+JghTUNSeziqnAFC6D04+7AE5AZok84Tq+2/lzBB7mDpC4ev4CkNTifk3
9xJmDc57cgCc+/Eud4bpZqimh4E6KrYOFC4WGfJRX2BrfKTb52uaIR2BzJ+Lp98tA8Lpz3HPjCiN
QGix1GOgwjBm7ZZBPIjrIoGFfnTW1oS01xmXLQfR1+a0N4tXdPurFmyfihGd2pTsHvbeUjnl5gbQ
3if25JjRVcWonZqX6heaNmoBLw1rkFKCAY5/Pv5aHNrf/Wv606GE15KJ9tcFHk0pz4pUCc4l/deP
/Feqt4V8KAVzcB6OGb6DJk7J4tziq8OMdBVQkjzo65qkvmSPVoeZCHCXRnjWI2ki7yceyKC1KygC
d2AwLBNH50c8VXBlAlx6G2NfUqoyahpSmOE6vtUcdgtAQlqsoFUUr+mAHf0UgN+iUHRPxH7CfX2h
28VwW2+Ewtca4jWqYdEMtvbpBo2L1qP22fu9SRnFcVctkQD16y0spIM+6Mx+bHSRPh64Z/+54eY0
+EtohgP6FBIslXvZ882tDuutHAu73sI7N/zrjOQijI+kWsmzk6CarEjkUzv2sIOFSbx2Jcj8v+Ml
tEpZS+a+diw0wdKH3XqEHqDhWYIbQE75dpA0hv4CTrPg3L51Iv9YRpJjkSZpGgE2Ut1rnX7ZIi4H
Bx1PyDY8N0ygD2ROJ27uspH9Nwykbd6MNG//hmDfzsHp73SS11eVENSjGxROvKhHsMLiU9b9qscj
dXSxArODFnnJLt+GRBRNrG8/Np0dPVxpaprtWrLnKpD0wHMPE/bpCWnydLVoO2rrsWCuTGe6VmPI
O+4IOr6452So+NAblJEgAiui0zo7LgEX3MCGG+dIc7zR2S/Y+N0AappuUUeiBaPJ65JjIxQ5knMJ
Y91i8ob08F7pFPDMAJGpy5sSW2gz2OOun0NmiLF1/G9waRNhoBnCQsgVLZrmWW7ZTX2LCq6Ayjrj
pup8LvfvUNgG07pVvTzyn4Cn9PceiehgPx7U4/tNKf/dzf9pjKVUKR9GTS85a/abaGreLv3tl5Li
46PDUIvtd+4avGzCexsc+PjzU9qWkm2/DdMSqnMqGFurwceIDdKYCGfYy/GG0MWZA4F6pP4TFgBh
G8czdzQ0hruVbMJdEFoasR7gjZg9oBkW/1NR4MyhZnsb/S9yPPNj9GhE/KeALXlj4pbz8PJpIwfR
51e8vkqF5Bs3k/+yt7JJcFvAk0+aWjbviCfrlf/7AfOumMW1Mzubffkx0Bg1L7tyoQcYIgGHUKL2
Qs8xA6Im8Bm7D6p2JC20j+QRIAiBApXWPdu/EwTr+6XjyvMEFIZKJCfo0kMr8djI5Bb91pZv5UTI
EHIoIIK/i9+Gk+7++KIZyrh39GOU8vsgJ9his62j4BYOrD1WlhQJwCPwJpeaUEZLQle+CLZHgJ64
zBiXSxtQ+zg+Tmkuk7pUIGo0wN/E/TYDJJ8VlE85lPxSTKutaf4GVKYHIk5cIXAjD5Bp3Tg9yFxc
YlzZl0v5+eegl6DlHN4KlNCtsA3kuPKyQkbAQylf6LuPF8gp8Cj5KNoUQVXyKM5W+aDItDYsbWkc
eTnxDNcoCKSQc0zpN2l8prRoO0VygWjk77LaGs5123Dq0Zff5KwTwfV6ANQvWp6sfDpa7F7XGBjU
qlXlSd5/nSK236S1zB06B3DqyTnGMYuW8PkDRcGHpjkDPDZx9qzVtYIQG99csM3tZ12IMIWTw1T/
X47H3ozVYmkRe3ScYd0JfmqcvkFRpw2ZYs05aS9SiwzFVOqcafU+MXYpNjPHcG/z7smcZfkqDQfm
Zkm3oufO3dHprBsiNHrwHjOpxoSjtw36nD/sXD+ejm6+OZq40OY0OG2tpVDTkFkIFvsXB0N7sht6
yrTW309aiizPbBufWw5bdoJW/1PgEmv12ITZY6wS7VrRQIuBReTfzzQZZ9OHT4XExNXIfp0lfgcB
zRE9pwBC019u9QWo2BqaoF9w83/j95fzuS2t4vRQmuBqoWgfvaT2E1EFELIpMIUUt9S/Y2P3W5zd
yAdVG5+8bzP7+Q330zdGAbwUQvfM7HtM9TXuWsMkKlgg+FLdxRzJQtuNrvyah3D0pngpkT+lT0zw
Xi2/iZVJe1FESxMYYWxgvNzW3bfFEk+wWJFDPazyfR0SJ/7Ql/uBMbV9V85m1QoQnkz86Vlx7T9p
NJdLN8sM/8OPlRTNXL2CIbcJt76Xibsqn9EaaE6QXvZuXd1BCiVAD758iEoGKQ4KsOrsVlQ2kqfI
0cLt3Y0FNNrSAD4HUOXiGcEzoV99SxzgWn00HeIZyBoomO9CNpmf5c4sPx3N5W5LZWXJ4zW6DJpq
Tp+QsrRD+VYTAUAlngvfv1+eTbRLfUSh6CpLlA3Pc8xJ8Fdp5e71LHyw7Hgl/uGQn7vamNjl6TnE
RAWuUkJzd4TjKIvSt3vUlzbttl8/MjTbXBoH5gDATOxuSgwlmzda3P4imgnMQZR4mHerDFZi2xq9
pp33hk2o8TU8An4IjwEp4ux5u5mhqPHp+Mu0bj6yrwOLT4q2EpAYGCXVITlZP/mEz3W4U8C3OfgG
MuqMF+0tjtqN1r1/W7dNRgQXIrVNDsGRMZ6GYtXPJEp5uId5KLbExdn2HxwoinRn5buEDOkFHYRy
/iN29AvDm154lxR6HLmxf+Dcg1185i3WTZVmnnvhxuDOjNlu94SiwzMl6i1rtJ3oe1JTaH9WqlAa
co771rvS1hCdwUxM1zL4J4xOR/dQD+TQsqjOp5XzY8Bc0JvVl7rCNwmzxDwHsE4qFAgeG9BvT+C6
jePp8ZCPkJpvn1ENnfV5rhBHYUaDGoby8S/x/IxjUrouvbFgOQMoyNy2hK9Y/dnIjLe8i7PYdR3J
5dD5DFnzPcrCSRdNds/2ZEBNXkNG6aytRmwdiqo5RBv9XV5hxfBGgpl5ZklXoQZT9txN10PEuXsh
7ekr2FACL7eJYnmfWbv3PFhQldZhK15xWcbEtLWGCxYvIWfUea1guxgk/Lk66pJIczyLBLznJz0D
ohovH0Ju5ebY1Zlg9ONZi9ruBvJJHuEWYmTJiRAnjlOn4FfzHHbOaysWQeicZ9Ll4QiK5o+kN8Kg
9Q4bSpRQJOjJrSwhacFBqMhGpgdcLQFyjwJXG9WH1JuxtdRVv5+PHPrK1eXEt0SHDJFqyEe/jm/M
Xn2unz14v4vJeJEA2TnWPvWdvFaPGgNm9UQOJuhv8fjmPuV6YJRc3YCt9At5G7iXrkfEPEFeGGd3
qy7UBnOEGgQ79fPGwA5h8KLcP8b1D1bYFKGq+e3efTTWBMgHuz/33+Y0HwC/N7KrkzETbK++/u1X
e7eM5awVXRSWo2bo/Uc4QVcuXBo48h4s6knU+Vzvlz4O/7cNsoVvPqvKtDJQ/Zutm4Rcg+5oBY6m
jBRU90448FO9ov1HmV7jDFTRxsW1tmefibGyL8D39JZcHaqniS4yLdMa6Mr9RGdJCRZb3SI3UGiP
TZY7LiwY/LMudGHCQpQQDN1i29t+lCNr9Xy1Ymvuxq/oA63uZjrIm51qRR6kaYX6w8eyZBqH2U32
uI8ON0v8NRO05b85hp+ALcGcY0ijrD9njHu25aeRZ6q6FJmMU5ZBWEzTL/bBRjZRMuxnGvL6TZdG
XdYClkStRJtQRl09sPcIx7J1FUVxv0QLSbsxa4IkU9PZacKI0eBOkV1Iwgm8eRjuTigKo1Dnxj3j
n7I35yBk2dXdGOYIi7s6PIyC9klHLNlBWo0Wdd1744A6sjBKaZGC84NyeLwVlyKYMGPyVsejT9+6
GCHM+j78+iGiYsC8jykCSxe4ZnCs4EM6mOMdEMtRgBi7TOxz3lVEDV0PLVWGMJ+mUAWwxN856Ute
S9sZ0BL7gxtjB/U5d1QxYrDtqT9i26cgaM8Lpi/e/gcHGYblYBjMskif9tUWOm2PWunaRCV9ji/Q
7DZarkWRNH0WNuO/u2n72vhiF3lZ3XlUxZG5wMa/zC2tkQm1pKHDRnMJjOkWqhP+HArqou4DZYNJ
m3jPRQADEYtCR+6hLdD76Lfg5MoV+Fg5ekf4h4RjUKhsPOhumZBpe4AFipei3wzYMup4vD9LCTlV
7oJxeO8xfhqqn2sY3Ja5aFA4DnbUzb1rMrzSsYlJRsqX9L5H7JdKbcTTHw7E/PIM77nzRK8FR6gk
RM0MRmmEvVVLFj15HLQpxD6oFD26fxBr+Ho5QM7hgwJ22aCrgq+CAnitpPuHz7KmsZabK0ewxiHR
zQZ9S5uqtFqHZPXD+qGeojLb676Id9Egufy3fpcxH41/JjkdbNGRf8TlZq+1faU2aloA0iQ79FIK
JhmnS729z5oiD0SmVIRJ2SEM6/rrvbPUAoE7O+Z+ahual9xXa5IfunbPqshCDAJU9CMMV1HKtcTT
Q82FqQdu0PnJyu+f681NcilXZ9ibeJm2JGnrO8YoQbnRZefmG6w2f4iyPumi+JbcvR/F0PFM4Xjl
b8SxiJIIeBP2ZC4FRtIdgK84h+i7raQ7GKBbYwHYlX7MrJ/lj24zC65mSMzfX4jKsZzV6I8v6iA4
hORdbg+hWw355ymmtPqfkZ/YOv6oZxpUO4c3wAJ6XA9mt6YTUDT1RIAumxczdusvvqdQ9e/DZjwN
8rVZlvptFt7yGCk1MZid8+Ur+cTfxDAU5OAvCEkqF/FX3Ol4Pbgdhyv6nWlwOK8oj7a2tsC2XaV0
dxHlWoI8bQVSrDHZkUH/pyE3ttgl15nIJsmNgkogQzBNgjEv1l4YlEdETHBZF8mIl6d+Fat515Du
VOjeIzClszwi1rgujUJN7/xTM2PtadbM8KqaCNzdTXGWIP6/+w/mp/bKoJBXyEVKi1tWm5DOEbgg
XpRT4hfgbBdvT2vFgZbnkxJxTNl/ScGFsUQa7hj7VaO84hTKhrtMEdTA4RChKAbaOr+fNVDwyJ3I
2lWDB7fWYzqZtSDmnma0+iZrMpoSWyo65w1iEwihKsizXHu5l9jfBjv+7ITHMAaDwFhxGc3rbGLb
41Tqb6g8so6clvZqzkQI4EwosjZtLQDwWYzoZgoPXCEasBu5BHDCEO0eLN7qs0jwQiBUwDz5gxwH
cy0ZSv7avHyTGjS56fYVzo0SriKBBphXmoTVt8uwym+MpB2ZAhwr8zvbi5JFkKlbF8Qd+HBa8/Is
a1uELw9Tirrwb2L5HtHmq1o5Ax70byUIxT+slfhVjQ7WtBxQmj5+tfCpHZ0gZJiQLCtJDa98NMky
mgkAx51YLFbEK4jGbwas+TI21zJs2B3LwmJ8tvmvuEMuDtvbw5HO8edj0DUQ1pQyaklsg7/fd6yk
dNATOOeO8JKvqcEq1XChhYXJljMoKxGfQz87Zztvxd01F8SbEzX8LwF3POOTyiRvORSA7pKeAQqP
DWFZOOFREEFSxMMQi8rZ1hORRp1a/bBEr2w5CPjHYu2kQ2RB5DfbPXckL958dAHY+Uv8rz1u8BLP
xQZhiMkw7NMOfWZcfsI+XYbW3PYuIG0SRnGWVF/0cTjlDng73v8iTXUk/pppoacMrvljE+i/ALhV
Oh/Be9m1TUHBCL6pntbBHyymw3EYgQKO5dlUQYmBWnEItyRXk0wrQSNq62kUNKE3SqvcC2HMy74L
PRMk8c8QQX/iRqehAUkMiPo3dRLR2XpLm4CAySLFhLpVeKSqx2TBNc5ioHTDLloc+9ka8KzTuP2N
9BNuBUuTjJ/aWtHBi9gJOvxK1iv5IxKUZcw/7i6DV+xkWV+BZnZTLDcjGVAndm/L79B+Js0C2Oop
GEaFDwxR07wmFR1Oh4V5ZWppt5yRsq8NNXjTPOyviV6fbiM8HyUiRXgCysaUjMxv8XO8UJE5sYvq
SpgkR/rRF5O+rDyxTPvehTGlFU3EgiAiVApqAr4QN5ndr2LlnBUjBjGXm0efoo/yDYSLSEJ4/eS/
PUcEki8tSXWGLZGm/ewa63EDdQ4JdIjeV6kW01hYVWQIzAd8G6sjXZoiajuP7/MuFJ2GJ/n5jIDd
SDJQwBPAU9gKBlaxNUbEQCQyDgYExcOc/u1yLVuJ2t9vYKY2bFpf8S2MrE7+c1FqpuDPMgymwmSW
35iJJDy+rk5NURrY4mJaLvuj/IVysqDb05sqt0+9iRVTFurOq6Fxzudy/nzXy7J9fEqoq+h4argd
f1HeSrvI5g/MjpLlYp8C/OO7AoQidK5qhAFsRgLHNh3dAqf0A2/Lx6SUcU9aF/MI3U4cUKUIDbSS
n9s+mrSYKA43KOT8yXbCgLITtE3bD+8pKSROm0xGnun7QYcAijaaM+cyEAPkm0SmUqJIphiaV4fx
YWUtuPtvDxTrsiJZAP4zE/XY+PkkbeDvsMTrIVoYJWaEN1rhAxXY+ikREYhWlo1dzp7wZt/0cuMp
W2p9KPwiVz45TTMBhx+S79S8qKgGEgTAZ02Xc/5HaoMyvjbECPFA7ba0Gss4SZ/uuDAnd4dcg9dO
aQvtIlM8NxVE+zL2G2W62CLGs4ADf8jF3UFA6jzFITdKxOQvZ1K7Sk3v6+XJ3ZgZjpOCQl2UN8Ge
Gft4L7NaYww4zySLJCeQHvaPNnqT/XFTFr1cajmdai84bJDTKrOhjivmoNCRn+rSYGJlejiSLZNf
/LAq8+Asgoxiu9LRQfYhnnYZzhsci88RpcduX08iY+Yr1r8D97NXCNI2rn9Q1PC3ipmnHhzZ0Rxq
fPKMtdKFBGWcvZyhtCugIihrxYXexb07mmug0LpXjFem855sxC6Ni+IYykQPF/B7DV8ww2/zphIo
JJlY5G2qBMDBGyAxqzG9geb+nhZX5gLrn7a5IESC+MDHZ3jLYXKiB40ZrwwUBIf73A/UPCQFMQJi
qXRj+WoHgzXuBSY7ZWygewVKmAA3oUaeR8y8L96b2yf/a3LumbCRxLEmsV1gWX/oBBtg/min60gU
2CgxEt5t1iT66N6x86RIe5xXyvEb6T2OH/otF/V5v8sq/dNbvmwmzp9oNrudH87tY3ry6Sw47Adm
kiyuKdLV4gxH8ERR1Wvcu+O1vfevGrPOvDq47yS3s+7Tt68TBH+JWUYBB1FMM20JlM8md3m7phNC
snRx6FOXBAb23QdUU2royzvp0awwu/+XCoP2CRjYVu62e492j/KCWVx/7ye+pS/lovSX8DRMB2Fh
seiL8MdtcSU8uzWjg5pDMcgzwkZckPTaBIJLiGAJ4OJRmeQzEWvtVL5QPQ5FnDgJghIog7w5TtXH
ypXofC4WnPs3fRQ/OKb4wmYpKmZv9d6MYFALvdPohrAY1q4RMReG7ZzoaZhGu6Ic74cl4i9NTzcM
1PPx/yzXRqajRuRTbX4R0xz+Py0mH+VOF4Xkl5d6kRHI8Yei2RkTH2bSKsuspeM0+AJSHU6IkHxV
u69JjBaguao4DdqkzrFTogz4Et2EZ34+QYm7WjyW76mJ5PF0mblxzv4fikhYVzxZnCQKVI/EJkxZ
BIaXKV+HBu9CzNnJP2T4P/eW2xIO92P3S5yJxPaxz2xxXCFp7DqXKuDdUzrfPkodea3cCWfZRcTB
xzbd7QTss6wk2e6qX9XOgp1wc4QPKX+mbvlYBchtdREEZTJJljqCWYhEhGEoDZeJ2fbCUcTLx2Xd
boPh/mpRzW2MN4WnL+6MTQsaTwMLroM6HsU/SMdHzt8J5xwRQwSidKRJIQIieUEr+rW+P2hsKLGm
dDlbggAn5G1kVBOjLfglqhlGPajpOB+K9EgB4+hsqTFwKt29xCwsQi66LcGYtj6Bx5kVEq+5IJ5b
tp604MaHqxFeSQLaPTzZvuzdud0mk0jNRmVA3VN2AoXTKE5QnRr2iHx9b+hB7U2D+gOqMfoXszay
o+wMSfGGqtEHF2tgWqfyRqd3K5x0NRX9m/n+uVbTXJ07d0SRSvCKZ0TYqhR+urXA2hhXcZmHjvRg
KPIuMA86DTQk9d0m25rSZWdwrXPRpbnqFlZUxb324iFNOzBnpWe73oqT5qTibIuc22QDA980Momy
3d6qp1ekg3goW0HKbgDXzJKSagZK7cCkOR08uyBx1tTtcsIlHFmA7Ps1j5zYJVwLmATEoHm/o0Cz
bUwUNIOKx3B2LGfyEzeW5KoCUaEV68dfHENot3YC8ArcrBciqqbbmZdz1APWR2fmd4a4XxlwL649
r8h+hAtNZx+LuzOt4UZ0QfORJfOKp4BLllm3dvPVanymQf2qC9YNnfZAvwLpfnFsJt14MXIUH+zg
Zgjb6eH8mtYKm6VolYhwLkKKZuYi6f6exeAXx8RFH1pK90j+1LCgMn5VcKaDQ3xvqQl7uGb3f41Y
et8jLBiO4ihgc8zyY1uOSCPj1xMPv5KiRsG9d+nW98i1Sr4Cd9QU/oYFpZJ4tA5CeLkou5/8VYtw
ftFJA8HpHryQKo/o9EQk52Ui0m8ADZ52kFAgJtqekLQlegkRQpeEPAcsnUsbhfqnCvWDdn9LCq4j
vNkvuWQcUoTLGZXzOSPTnqJKMQpqu1A9S9+SK2fJ0T0Bc2TwRrs0RC8hB7X84dTTnTC6IUyqsC60
/uRLm9foqCCNjLrCEuMhA4HNXNvtW5Z8Xg5dzN5BZw4zR7o/xmcS3L6+O+uXv7oV9wCgZOKQQGnR
7oRYepP8oxaqDXFgEhrqiae70cd62zVaL8ppwSHsAmqnf5Rf+C29f446oOeXLHScQCDoa8mVLJu6
l6wiO8qfomo04/Md9MFw69/GB5VlcGhSG4L3W10lAcScEGzGi61Yppaf17kYz/I88blXjlUwo0em
L6YM81aLj8IeemzDpI3WKvVKHC3339c9S0MjYijLXkXUkn8VgJC5ARtfTu8I4P5BT8p1Aq0MaA4C
etQKGwK3Ib4+4M8QMvYHOW0bR4rX/g/Eu+NapDM80ibDw7WOUbDgN3LHwCPq5XecIlXGRyadrpKW
2EjovNM9ZHv4snTsv1+orVavFl+MrT3yF3v6X1hYcerlG0KS6acCefmLfzYIGZZcPeUxmQ/d1qpb
OEiWWB/7y0fw5hMO2P9oifDpWPaCHOvjsdweiDeepub1pERJx3xK444BJtLIOSojFnFZzkL/BEdD
JruWM2Zoq0ia4mxy0i1YuN998PmZt8RJSVldkGDW4GnGitFS0guqPBKPRWnhtR339CASNwfCBNvk
LvvuC5V3EFASwEcjePhvaQ3aAGO6XKwLU+wXvEN+uxIkypsWflnlSrA/qO4m2qIkc0367lQAHLQd
vTwaXKpN8SjA4thos3ZegkKk3oaMegZEOLWhg3SVrgoxRDXR68i5kcxieJ9eswvheyhseo6woNF6
cWhK754vU9dSiKbmHMMfgD5blQtHjumWU/XJ69++svVi556/ELygO8jWHwtesWkbKPOZ2Zgn81LU
zNT+R4Re/CWW5VNCRE30Za9AL8l8W++tHL4z2YLOf2iDAV+FuN5TFxrj6exBRsADwu8SPpF6l4nK
4o3LAYLpE0dao4fLRcWfWBlFjcwzBZz3kFGVdUebcLCDbBxKxGO+ig5jSZEmTyrKeNVuo8WgYaAT
wfaAba8NvUVK7LhK0gSKlmqCPB9BtK0ZWziCIu9pNrGQiuUUjwMBwMpwlFWfCqNzVrg9SgaeeyGu
42Akc719zIjWXaL2E1jLp/6s3AFLGDOnJfiGPS2VY6z0K+jE+iENOyeBgMXJs3FtRRu6tAn+YFhw
56cazicBoVXHso7mUOdPPYib/6UuwMewaBGiQvNkmXXrWsTYso375dO32TZvMXtoGpLFd8BR9fk0
XQ7UM6qMf6YPIgyv6BQI4Kca6UY3ppSPruHnJaWPETOylGskjZ4nXJ9NXpn00klPbmgbPpLlwO34
NPv5LQyAn+xMcIl1vKL8ohrqZMsJYQ5PHmRq/l5imB5rC2EbW8Zuo43jhyYDxTJ4Jzyx4eiSDDOE
PsrXWVLLDiboTRRUiA6K/oBxGnaioUmPunrltXE5OfjCYRcM7Pu6pbKntkfK48lMByGMijyJaOb0
VEBgP2tftFS/xARL9RMHq9cKOyNqZR5QloQJ9EWJnAGRWse7vcWPzyJqjflXaL6Lzgs2ZBaIXkKc
4Apc9Udciyp3iAxDHizw8H9UpVsahGkHONRu9/bz94TE4AWF7SGKy5/76TfKUCjXck3QXvyponFG
PIahCQA8/avWY8NUitgJhf+1OVhMVNSb4U68kwd1UTLaxx4mUlVKEiQYkCrvNsZEZnW9XMy8p9md
1b7Ky24j8s1+jlEuMfB6FBHZuwOmDkEZC21tK/xSu9Rcvbkzzbu6Ahp9T8ynngFdEfGJQPmZE0SF
goTfBYJjWgHtcuAlNHQi/7FlNOsgDBdTJB2Glrj82ss1XbiVPBheigOARI0TwiPcC4KYafOfYNAf
g9v0GEwIkQeMGEojcV6c8lGRxFAiw1uMXZDTayLrAF/M2gu1S6cvGvcagxvsFqqnQDhW+tpcaWhY
KUIuXXEV0Sk6v+uMAQGhuIj73UrDPCE3TymuJe+auI0bNGkoSNcmiUeuwZgpyKOIZbGPHnJwgHpH
3UjGHlH/IK3KljJgur2V5zaCZD2Te87gCDCJbyN7xto9dEU9S0XIWiCpHHm97FRuaLR41JJKv8yR
fq4tcdGr1AMigUytvs+ElpBmAw6NRM3beZVql69gAfNPHdSbWER8cpRwgaljjqljkobxJBcDGjJl
O/dumIPNdbPZdcm0wJnRyptfluXvSvu4IR6GRLx4nvwRseAESUW93J3NQqYKHXQnmVmQT3dnYcAw
oODPmAbMB2XWjltPOHLhbWTj1HXFSaeTGi7n8sCKOX0QJoxWYDq/Opys/S7uFFOctUdl9uve6iXw
j0ZvLvhn2V8ujEK8kLXzl2dMp2a1JxNLSsbXZXhg3fe+JpGxqyMD8/K4aPk+jCIIT738lf9y6cHq
fbommeXiN3JPXtDes5pQP3TCitZ9HYj+ezYoyZH53wEpzDehC61ZNJ82QA0hpttUxeOpRbd1ALRj
O+rCRy8JH6oAk39NyeTXvjfIJ1dDoryA7tlXX5rOnpxZ5FCLSnxaloh3iJIbUP5Sg4cvbe6CMlJX
hqlpV4o/ONvoA1Xf20W5ivXdXM9p/y4QHXdbZEqQ854gVZMouXcPo5i7sTzJ5jJs3GMMCc14ENJ1
bkenM8bNcYQKB1QUCUfTAQRuJQ5d2NGIZ4xiGagNluiK7aTo7WTPQLUadMO6Ovt87rNoCJ8PWakA
T5NnyYdIVjLTDhd5hhEvybNrxe0wIqpgR+643A6n29z97ihkI5uGCUO3CY1pwj54ErRyzU3OeeZY
RM0bV33A65v76RbOoHQ61aZ2qFndHAWoBXBTpYNiY+bSQuAfIg5calXWkhVkQkY2VK0IphEz8edI
tOb3FgFVDXWDLbSxw86bG9tJk0EUaID+c52ORU+8bI744U1axJ7MR0iiiGz++4kVZZKpmwdgXOLJ
MTHw5F8GGI8IslqmjYZSghSjYBlcwo97HygGEGA08TzWLrNhEHlsf+bYaWY/iRe4C5KSROlu+WK1
rsqxdO/8IlTNF7kI088rRGKgzopb+Bu12iptBOhX3ptrqJdAkctwkztjpl50q/v0Ek04OB2qpil5
Z/aAwvETXXXVQKMxf9Zn0hpAoWIxjFAwKKtlLneEayFUvial68kplVYdhDqXXepH8RtPZRgjhdZb
29tWVbuAbQnz2QdwUTlFAUYQjGEExGJtGePZ739KwSVq0VrJ5qmoUU7U9MaFW59BF+gbCZ7nhcYk
VCVwgf4yFBtHU8JNYhtEy6P82laTjAqI+9YksZ/nUF68um8h6CMXLmec/fhDtcfed3a6/CK+yqBK
riKiZ85jlLnEGfZtQ0pig0Z5hsoWrUZxtVXDE4fztNWZ7qrmSM1gBdXTZnt87nSY+dCrEom4EqSj
+ezzHlKTUl6y7l1da2fD/YXzgX7NA620HvKKHuyaHLUZoO4HNdSSyfnhsktnD+ZAj5RmjN5O9RbW
a1WQqFgzOMiCiamYIiMTR2palzEemxhH7B/31HqNkdxyJ3YznOykjn3mkUIPsCfEEsU4LLrnmZvX
xakNZMLSsC0wc4NmYQ6Q75Wag7SOZBPQhXZsD5tVvKbkvKbuBwpsrfi1JGMdksWZHQmGqyaG3Tss
NI0/Zgw2WaM7Hk56r9NRkI62521Q8ob6cuGkjtDMUV1nuSWYYDjhhxNjVQRsKMu3pKYqTg5ESPdf
IIX2nfGCI0YYD2Iyx9sdz5piLsg9mvuTSy317DC9BQ81hkTfcAbzp3SuxuwYAR3fOxmpPGoQfblG
WZa3kLR9eFXmP6bw2BD5KPAs/2jG98coWdjZ8e99xqoZZYmqVEzo1hdTWfanj/0Uv2oPv4Kc/Fq8
I4TFN/P8yN1tPA2mmf7d+gUUG6yvk7YvP+sWzYW3Qn63PdwzYKWw/D9dCX1UJOOl6EwJjZFjgFwY
Km4khM9RO/6pMYFIirrmYUqh1PHVbSqCWJC3pJsG4KgohmSpHFPkuuZF2k9AedM/yZtIl6SM+A6Y
HQkLyvi81PyGSH8FmYPWpqV5ULa605bzUvdKjNqXOmXMEZjWosJmMHoxamLldOZSX0ET4ayS0sJG
a+VTVDpYa9dFB9cmdGghLM757B8d1oRf3rEJwGqVq2nXVPU2yRhRAKx3kNztqt9teEZ08SvSEp+Q
vqeE6TMMVWOxy0GQpJP2DXP+s9kC9d46rtDmnso9ZmJycidIdwCf+R62T3XDw6B++DEcxb6GSL6B
PnB1azYLLHQ4X2O3zYBhendjPhcB/qQoc6InxXmd1WDZg+8MVJjHfhzVXLtpAY1NYUZmqGuUC4lu
N8HxCq8zG4jTjVAQmFs2M1c9q4nummMd/gIHno9lfqPTMd+tx9U39ybqz7nQFVhsDSlzgqE5z+Go
qqDYMvQ5ByPgfZlxXWAFAWfr8SZsOg3X6wbICy8GADqysph2R3ejVQDkZ5L3IlM1aXeA8rnwDWxE
XHzS3UrV5H1SXxIns34N8NtUvu8TAZ4/dB8eOFRT2gEHryCB6lPTAI8QSpW/bcCY5Yq9aDoQhrfP
9xdCjmrramyW86Bjvw16R83wEDFwON4qc8puUvVrVlRQpVcaWkOOe+/SQ0hRh3USCNoHQt6d/Tg5
vsD5meWbkO97Q/BJ0hd87M26MibUfp40vPa9WKuACSDwVRvktHPC855Z9B8VJLGoA/8kJUxb96+G
GgzFOA7V/eQs2J7v16Fn/l5wFrJlJtCEm/dc0pW+i/+osMBWmxmWl7BD074aEyg1UZtzT30KydE2
aTgPtuxBcYV4P2+zHXGI1tOBMwM7EdhE676fpfLbGNY6QBgarfq+X2tI8Emc2FzaHN7W2ugHe2y1
68Qz8F8C1/IQL4hWm+ALJX1Ug0379gRLLVHb6Dgu/rqEIBciCvL/M/nBzn7+6LN91n1Nvnkya+Bv
sdXa2qjya0/gU4YAoP+dXAtVJjsjPvJHzA9ZImFmlidV/FRpI/Benr8OQsG6Mm6vGQfD9+mH9xcI
wpfoYcP4BnI5IGRWR4H0PxSbav/eQXWgl94pJvjjpzHPlrYTCgUeeOmMTEwig63j5h/XeJ7goqWg
tiMqeIvYSvpOdT06JVdIi+ApPhpLGzEiCCeNnjVIA2xIMxguDjeh8Lu3NfjFmWH9QcbM50bRfW67
AvWAwhhNNA/1tseXSyJHsxxiTMEZIqJFaiKEGG2pAE9quWEnco+Myyx70RGmS3nKoXQbMYn6wzPL
I1kogDhqAX5d6UbD6T8nOOV88TG8EK0N/sESX0q3jTGYT++KGDUY+dMh5AGeyro56dsboYyEWVUR
i7mjAd4ZywXr5IX1yj7ipoT0BtegU6kf0Ccx+OwaW3VdGMGbR+i2Mb76ClBO8qkokZnLO65KJjDM
reWNFj13OUPL0vTIbc/LeoeWOvpigbvMqScR8MvYF4C/zwSjT5mcGbOtmeKMxkO4GMKMZBILj4EN
PVRN5FnUUXSRqPitDFUQd32uCZ4qrK5tyaAFJA0NVzcS31LnPJKlPPCgwxBN397uyvh4REctkxHb
RVwCMWq8IbDB4xYK3dJGdgW3Exnd1WbzRzpqXXJ0nHyE5S6FJg/nXJ0JF0OsGsl86/oNcXhNvh2L
scT6jWc/EBXveXvDlDzDb83nH/eaGH64HfyPxDzZkunQz0owvmPzgawkQLEbTp62fEAkAiTdbEKe
7PXEKsr4tIJJ6NJ79ST04nv1TBileGURfSFtoHK2GK0l2pnoZZnWE/kXK3J4CesvzbxVtof2qw1B
nrmbGI7rL9/dp8Elkgfus861NIanQLQCM+FQTWnner1bU3ledjLHmhjxNmobkbEIE5StPqizhOhn
0Jh5XeWcT8tNTpMOBFk0NLA8ujp1dhiAARD6/x119WfgpqB4+CMKVqF1ueXfCDUqkLpQBYUGDiyx
FCpHfwag7Xs4TxRLa42wjhak9i5YDts9OqvXR2Bs2Oq6JfuMBxTTpyxE5LgwSkHR2KmOi35YjrcH
Sr//uhPCjhaEDzPVnyPss2v87O4Mu1nXhd/AH0NRsjCEb+pdC0KcQxOlMC469Zj5BTOkS57I562F
db79e+pFHR+VPe6xb1MtBDVnXN17+4+6Aaj19vCu08IF64ehhFZGGgIEc/OeRGrw9sLyKnvT7LyH
+BjgGpnAXldb+UH7j8za/zBDQ/HzcIU9weHWnj4W7qe2LCFU9GMICl3QRt1beuPA0Q/pnE1kVosJ
qlvzIXcw8jGNdqrNxKcmj1ddJh1aerCbe8sR8HkC6NvJeKS0fecY5ZpJf8Jx+jlU6fMtLZlGQsqX
xBErzpeXHiOv8LWM2hQJmwWwval620uzFBgoYfZ6fpaW8HzKAbO0kLhenM7Zgmoh/bvBENIuAM4N
hmcTN6YvLeQ8FVamf3vOriKG/DgrafLKQyzto0j1rKr+U/EaraEOHbn6K7iRmlKpa7ct0cXiOvUZ
iwxDUTQGab5046i4T7L8OszfUaQzQS0DNt270KnuB2YPcu+Ebjqkyo9aXUxQifJ1OTXNeMNAeFN6
unIw72D03MJwKbZbuRn8rXUMEorWYA+Q7yvwVJjYlWOpZK0GuHJYkU2mVQyprgbo/bAfFn7E58My
RT6j3detUMevQUmqkNwHsmUHKsWPf2ByBGlIZp/hdomUT4BSoCBJyWb0mbWpyKrWOOkw8B28O8M4
SXz7clj0Zx3ajJvy0AHlKBhDxBE6HYOUneOh2mGod/uK3gVRebm5VAhtI9AV0uRAQPGvuI1cJeVf
HhAi9G5qokCqCw97kFkNqShyagk1dPMb9chGTL5hQvV7KjWfO4FoQKGZJ0k4i7HsH+4Wz0F7E6h3
NWckHKjA/sV+Upw+EEOzXGgP5L085D/uuBYt7gPbPTILnibxyzh2Ccc66wXQzrnVOLyODnMJn0UL
CIckDf/VCeZDv13ydUs8c051/olvcK32RRgpVEg0YpmENCnmRcrAn9i9I4JVeV0g509YvF8l1Lk1
f5lU4UuV+t3e4t7bga3gYz6QFOK1Lxh6UzhhtlSH7/EtsYiOUTm9+eOqXo4Eswq+oeYrFIcaWG+r
SzZ/bAphpgW0Hmp8MdBf30PgN+++hy1S03u/u3FJ5XKNad2eJK/L90HnMebfB7N2W9p1QW85NkEe
RFBKwRaXI99D4NKmxZ1YSK/uPLQ2k5kZg8YkvXe/XsWVhEt1D5lL7lB8Xwa08gAJYrq/DMhb/5VG
aGJZpB26wMOo61DGlG9L/gA5Z+ChpuwKXnR64QdKJTDdqqQRRBSz7JXfnHeI5BAXJJ24PfbxyvFK
thyJlhoMUG+GJzoC9qWKr/p7UWTfMxNwzGth5cmPHh3QowX/p5lOvw3twc6eiFJfp9kjZFpye24G
UevxAnbc6ts1rbdzWIa64bl+ofSyS/foKJdaBrRtLUhzOK2ShnANKvXn6pGaZGaXP966VC4TC4Br
kf6BHbJ4i0CXwBxU3ap5ss5WyJe2rrkbcYf+zf/87WdPRzRQCPKCJhb5wiTL/Xuh+S8BLEmeUNDc
woiBTcna/lW+Y7mli8Cyhe3DrdWdSp1cjLhYsdq5HfrIZReZdLEbwCfib6LNlkXY414DxstY0fij
y8vXl0EbwDk4fw/h9+bke0FBAdgxXphMUuz8fK5i+8mdR4z4t2BOfngXEwuY73D13f+W81FBNYSM
1mV/kpMT+XkG7LGquUhgrfWRg8CRIRov1MkPOaiZOrQ0KOePvPCHkcM2pKjQ7luzb7CJBt6q/Gwi
FZbg5FFgaUxBnXrSgsF3uC+Tzrma76mfK6sOExSO+VXXXBksCOqdF5rH4WS6mkVMkpxgejPaY1Af
fOrxJDKW/W2KdhnPf94QMx+hnGckHJU+rYvo5R+4w/S/YwJ+nReUQ3i9dpW22y0PrTDWsPvBxpsb
hH4zrm5rvk0naBb9iU0ZVdH6uAUGr34RkhPrluMsv2HJ2KLMoliYb9TVjuWePSMLKGyHi5n7+rfT
zmtSXRanhvGR/S5H3DeyN7eSan8ecZZR3nTySmvSqAugAxDuM6dyVDYVKDX8xtDMEiN3gCTIyQt1
afJj3OK2lDi6FPJkx5MFpONSSoeayiyAuSbZy8DSRqpzdMK5Fpm4YQzc1WKyM/VGDVe5LnFdCEM6
YwqRM+Zwe/R/gdRIodmRkOpdhM1qVC96nCxOUJya1YbO1OFKpU79arOiH0qkHkFMiGeX51xQsTU+
cWb55pNAregZFbjV7CtrcC0VMavstAI8zoyrwzWb6EKzLlHykhD+leWGkxQ65clgiXYMYcgIBAYB
QvKF14nDlwhvVk4lzPB+nZeeKOShVPG05uS9Rl/V0Cy7pF4wX1C8F1bgEBgBGu38ezTiMo47ui5v
Ftw98mUtMP6i9qVkZA29IfzveZKAyfZ92xqVXx8o3QUYTgTXYPuMrcV6Zt9taSpe9mittz+CClsc
GcpSxRb5b8xeATMcuMFwrvR0SJNz3KnQ/mSzoHypK+IBJ9yjngoV2ksS2pivEsBBE3ei+k+sQEzz
njlar7pOLmbDynzTe38Mw0gqyA2e2xyMUh2iFRaVtrFaCPtDxYs5EnG23nDoiAB3/wV5HcmyTG/+
dbBhJv9ZZ4ji5EQDPM/UMkGlFiydGxtV8jE0B4iAmA+jRZ+/ec60nNh2y1pTi9W5zrY91d9SZY5o
eatrcHWHVhXLF5aQG4xen1yzMpjJ93faevpz+IWcyFPLGE8ZC35YHA/1s6b0LiGmwv6bOzdkwx4h
TFYF37n7qjzj/lK1pQ8lonlchhbi3Z1bdZziYRiCQNLJwxSQ50xm/Y8Xcuf2ULfPoUYwVmFlKmeg
KtdBtENAzairastKTL43t54+io+s5zVXXynWuy0kxr8XUvOk3SK5AyhCQCATpKJAoQTE3iZ0eeof
m7BMT8rRbT/1mUjrilTNSCf8b8okzr2jIrYBFTfJed/09+Lh8nAMXsV8wqpFEs3bw+WYTU39Z87X
oVBtetlIWCKmY5LytW+m1ZrCRGH9ovDCgxnrPsxkWMcKgyqDZVq8FDrsjQoEK1BReJ239v3H/6pf
fkN7wGxyEIM1/uJ6IOdPxlhX89GGy5dLNAAPAqbk4EOU4XdXVkN12ogZyORglJ5q6EyMe+3FmcLI
y3sfctGs+Zx7UnGU4mSZEoMfY6XupmZyNujIYUrMvIsxxGY9kkEcI0DyJG10d3nTOKZ9a2iswjoX
YK8gzwO5dfl8kLKEAcQGY8z8lEVKXYAHQ0u1PBk/v/8cnBukZKcy+k3WtXMrXtRPzp4PPHAwAsuu
XiFnx20xrWKk7bNpVANn24B426rPNobwrIF3HRfs2wEO4EC/xl1ok2bq3BvqsSqurzsLgbJ0I37U
sUriohB9YD2s6p1AbgrEGCmPC2KyQ1NIEQueQKrEIybN5kzgMBNwpgc3NUZ6dvwFnFPz1fWfm8Uz
sjkG1NDHBRDzLsm8eufLwqOLySPMpD8rC6aw0pLDtbY1++BRIjYu8fFvNcTKqawffA3U0dKAIMgI
qsoQoLHsTESe34EvplE1avX6iAQbmwaiwT1lk58QaVpUYE355uKjkaif421zY8nuk6wqkBIHYTF7
QiaZLvZ3j6eeFzT1w3H38ZxK/jqx3toUJIgTBPCQD68MdnmVE9/DE1TR1lTFonZ0Vht/nn6SHXGc
PPYCra0bDh+vhXV4L8GicmE7qmpp2W+gGBvffheOh83DuMvNL23Naj9xzqqhdV3BAl4QG1FlUIzy
r0JJdS5+zujVoFLefTcsCO1Nrc7AaubN48jeZvCXuwc4vqG5ez13hrLZMoZAfl6BcwEgfW07xVhJ
ybo7yxnhabqTeW5JQ+mRy2frYWzlDhgT3gSegCcbnw8/vMv4857krUJFNG3vuSF2A9yvC1ydhm6q
yQSxPMnLC5FoD9QzO6WnQu2JDkSwZLyRmPWjCDqsoaJfhQHZXDnXzqKrE2ELBAvUvD6Rat4+RvBQ
IGfljeaE5+Rs1Xh+q0NaS+wmM+LpHsadByCKD/XRYqs2P8pddzc9xwxOnupiRnalD7998HHywnwb
Y33aISN8okHbfRhzmf3iDG6x/QQmsj0cfN2cfGYW6v+RSC5eia9GTH6e/nZmiIW5xdN0TPBRzE/P
kDI1Yr+KdVc0ElqNfzuXmz2JKGTFUtE6yUJiIQ0XeE/iFM6BhR9Wzvglh6N/TN0YNcT+Z9T6dOLR
F8vgAWqfSNOmzpwjL7xr0dQpNN8GrpJD5RdJDSIf1MCBDdRu4yCo3C3N+rIW8IA+ydq3G0wjE5xY
qqh1dSHxCMA8fzw5WnrjPlPf5PT5QtoOSu7QQDQcyS7NFf8UWQ69N3SpZKT7bPmiY6PGPfQtOn+L
6XUb8t5MlCDdfW5ndFCm1tRid60dNo7qLoJFsYvp5Yyr/C4HQ6zrVNnuUM5j7Yz1kDT6Y9P9jgOR
yCia7m7DuDW3HMFl7f+hmR2ujZxLeP0cAOnA+UPmsTY2cQCyg5cvnaNQRk8/Vyi4sNGmQvaJRv30
yYBJ7wf2uegH1V5KpP2xBGiZHNNHXzFgBwflc/gJfAl0qb8j2aC3NZ+jOIgoSOgZ+4xZNtcFcp8+
Nt6jR6mYL6ZE2I68t2r7cfEqHLmIJ3ePEoehJ5kKbeVui5cw5pM1O2xHNZHfR5JBQKieLLfJ6NE1
G9Mm311HTqHWtJbJ47eKnV8scPaf/cc814Ju0Rda7Jq6L4dTvny5mQoNRARkqbP1aXHyPTj95EU1
yTDgCOJ2MJN4fIUuKk8jtkP2ILcMrLXuMJ12HTg+5e4rO3MPNc+vz6+OyOwJYwdcxOJwObC1kY7U
ZYQJBscrZidQf2fUk5VTaGIaRR33O5zGf/WhNcx+mpES2ZSz6YIjqurVb1RPgJYJhFmZAOPMCdPH
BC00q8a3fegNJAZ10+faOtEzQ/SHIb0edDMdMB+9O9On+4C9kIgGEbAHq/PHNWHJiPUL+tjZWY52
AfKR4w1fwZTmxFNr76+FBv57qH1Nu8Cnm56TfEcS1NEUcmtlhJWBAVGYq6dnj3flH7jgRFLOapuk
TNzSVNceVnmvDYvoFXmetLYYhvU5jkww/cSsEkcyKGRxdgt6eyZapY9QD8K/0T24K9NgYHxh0/A1
ihwTRiES4augs1dvhjhZTyVAJ8qr7ClTzewhhxGm5X7Ceml4Lgh0Q8gNx6C44I0o1ZhUmqZ2DZlP
0uYB1P81SLMPM5ZkdhOX2iVDhHvtVUKf5c+KdVNPC++0QTbYHm0XjUoSnNWYpX5oKcfcqjhfQJTa
woHA7MYrxWgbQdECD80TR+7ZLCsZMsaAt3hfPljfr0nqTFhWP0hIfxAyX2aG343x61nb1qyJoAzb
rtdnza6/JKzrzz/3aX8gLBvhgJMdie/af32j5Hoz2FnPk1UzdLbLnE7GYKB4in3sSleanhBFLw43
/vHV6AineN39fiZ4H5ixUFDHyb+PgRldtC0tT6q6c3k/EITZaYlLVCK708Gk1M3kZtE6qBCSs3h/
TLGS/elB5EZepnXfTAijg/TdsRR7UwY9AvIINH9T6woY0grTXUg9zdKsvRMkpAb8t4d0cktIUvP1
jdSTgV2Fk20XgXuQbJDgPm+HMVl3RhLNpC0I87CRBsfz7MVgvgmPFH6Yros3oU+hJmAaVrVrXKdR
rbsLh9cXAcFqfpD3RVu7uo5qpHKj/wLxH/Nabt7JHSfoF4pShC9+HHGpO1eSZU1b0MHc2LeiHo28
qCRbBv02zqsr6M4dWI+yEj29k9qEuS3UDtWY/6dXbwDWM7L6ZGqfT6PLWI4b9OWoIF1rEPu13/05
qkPDOQWNLYzp2LFy7HRnWX8udHbkmOzE1DMValuDXQuhLV6nBZ0435QoCcD34/Zw1A1NPqCPKaBH
9FqemvqTaPjI4+C9a96IfG0gvV4dWFifnd+HoSgtv5zopl02JipiDKsWkmD6QpB0vdd6HpZfMdtq
tPM40aHOAg/iPPzxyNxYcBaWq0CJzfotHv4mGJyw1aL8Y2rAdc+3RS4JO3dp6WxeXOE2+aA909LU
aSMjpkOwttevMmpYJZz3TYcz/zaiivuYx+w62x7BM0zHEFcN3l1/O/0nU1gK1xATIr6wsS5H5RdB
tEOpdNvOE5oahed2ImKchcelrZsYqn3Tc8Yy3g4iKF6YiljJM5p35LaWIfC1oXbhRE9w4LsmSVE4
4QdfmCC8HElZq6vDc1SPfpSWicDiyPV8zPyV/CIaSRnA5XPFhg3hS0mkNkb1CjRNuztCEZ4Huc4G
epCM+5y1FtPl+m14ArjZhfXIZlgRBvTy35qelaT8r1igDJstoYJspH30ChVMN/fn3DXQOmLoX957
pYQQTnGmlNwpoyVLSIhfPfGnRHEI5VJOk8tgsF4N2nOjjxMJOMVlLoURboUndjZ9qKATW0qq/NZU
UKufc7/l0jt7kiiwodh7cTdcFZJcYOeYydjbVjpZASl3zHtbe+Fz3SHsul9o/6UsUu3iIREfRrip
hWLu1NvGJGLtb6FG7SJpVKjfGlSFw9VBbf1733GTL5SX8s0AkbSihCKf0AcYSFdby+HOgJqel0kd
0ngfPk7L8FFKN4t0dju74KfaRDkPtYQl8/T4jK9drIjX8KrkEL/twUnJCGERKBQWRrl7uYdi9rhd
SsXQ+UlI3Vrp9zNo2XB7rld3PGA0bBF73RIsXzPYaPRVgExpxAiu6n4P2kd2jyB5pVyjj+BAeoVk
CK1yN8syAOLHaNxjpQZGl7BeOUVC0HgJiL2XZymQb1ojkKG9ulHWBboDRE7LT3e24ov3VvkTCKwI
TOMCZwe73AnFlOURfrE7dcRybK3Il7s+e6jyvDn6imFsnzJEjIwk4ajaP/rxtQvKclkHpsud4Cv+
VNSqi2PtMjqZGTPsS8OeyLGyUPJ5LYTHEkdXXQKGHmOr0njcYjOV+LT3ih3RalhJwk7oos8DixHv
iLot3owW4C/mOKXKAQFeYZZ/o6Lht7cMd/AjJVaovtnqaBnEnrHkEI9s3QG9IuYW+5BwiNg7UoIG
v0bnCFVCbulsw22gPvFHknh+G7p6B8qsZYEJFejqWR0shzYTAO5cLFtrnZuxE8CE5Jlu+m8zbq/2
w8b7VpDZFnscbNGVJbZjqFotk7M2SMaoUlZ4CPMldfKcZ2fb/OtFgkKQRVI8rQOUdVuf1rrgeYHt
FDGvk138nM54vvIvDi3/G7MDrhPNqHFhjYYImt1hL4+loY8WFDPX3PlZ960b5xV1DvwW9dYx8BXL
nor96zCDGIMGwW96gwxoj8CpmCr6AcBnT/sOtNy2WfIscR8Lgg3XsSKLtH5DWkV2mu9jpg06RpYU
bMussLrzKVGnI8ar4pRTwj8FlTmSwv5w5eeqz3jamrXpBXbZtjPDNrpqPIKbgHHxKscvkCmCvFQ7
A/NmN7UTV9k8Mbdhscs6xKAvwu7Wnvd9r9NxmLH8mh1Vms0oGHQYfpBqDFa45ocddy1e5JmtG0k3
fP97U2G1B4Pdz53XFMUGHAASRIRtdXTT8F+UgVQRK6+HxPpQVqHNs4s3RerDqA3qztdLSPqdFL+5
xmh2YKpTkh7g5V+nNp08rqpSQuzw/tzc0acrXYROATtUzETdPxRAXA7nXnMcXcrqVRX6QnX4WGC2
A4QY7fgmjQoyFN3TpNfl+dwxfkCXEPjdM27hIgRjCtqzVJYE0vpwBSfNk2PdBQ9qjApXvNxhwu6/
HsEEg47vHQR7Fyn5VSKIZlKXB8B/ZAxplzrtxj54wUFv6BON/5w2S5Qz/0919wegeBQg5wuuWXLN
FN3lfnHZzWrEyQtNqcUtXi9RDVnkDMmkuTBrdj25EdqAuWUihD4CcZ8wYNNzd+splO5224F8DVjV
EhGRrxn+JapWB/iYmUwjBetPX1Ar5qZTG6KYkAZ17JITRli2Be5QIOyCvWuq58JHZPSWjgxzEStE
P6N5kEIf/f87VKCzuBr2YSm2MCFQe+kQMqBrM0FA30mxA7qscZ2MmF3uIaAw+xGE9wKLkptbBfmL
XiIJCF1bE5uhLYgK086pRL0ik+EmNlWpWGs8SJbAJbyOJG0qbydQ0YPbxRd9vxTpgSH7Dw4G/9fU
jVY0Bhv2jDA3erzZOXMfDIi6VKVeNy6axlyfI4B7zgNWzJAD34Yl+i5xScuMqRXlXs0jumOiVCNJ
pgHtxjrMwiCMmvG38dZEoSLgNAMTXlNMSa9suLp+zYqMWNmJ8RVTXIa/A7ktMNPhZ1O66i/l+Svb
n7z6NNvI7eXng3we5HFCw2L99loX5DP3PysDivsKUVz0jM4eTSbdxNXYbfpl0HQxE6Ji5PoYishW
hRNMehwIo3OWf8Q3RC2f1Rnerj0XYecZ3LIqw9gLzXZknrmH7FrCc4EI52B9G1p9dzz4mLlUKmCf
4R28qMT5vdJjB3Fxg0qjJmkLZg74azaqXZAoAHpBx20cRWXcvz8qOSXaC93U5IizxiZ3HG+IMBAi
dKsnVmKQiN15QhjEA6KxssILyKKyyYtV7O933jd5bMxLWlWW2QcGL5s2nOqhVwtLF3LXvGl5okSB
10rMHboW9W/VbD1AngCTYDhZU5OvRHRiO8ZXpa9pTAOJqUKHR2XuLVMzIrRq0ayU4bNjJ0IKWW//
b1+Xy0NjflN+w+oOcoGH2iup8qGozHl868GQN03E7khIWVmqnjAN5rcfC/JsY0SYVPJjEmWF4+ZA
zQlLIumEX8moyvLxXWYNrRI+x5OYQhT9+mwDLKKNGBoVOPbMSES4+yEpy24E2XQ1NbRpHRtHfb3U
7RHe4OOjMOkGPG4LKo4HhhkHvqXEOX+KvZQ62n3usIw1e9GaqpVkCVMrp5LSZU2rAL9R6agxSOD8
h+0rhCN2NJBWZbWU6VG/qaO8ZWCu8FYgENZ80WrzOmY4PjKA56miImfoDqPLgv/MlVr79uvo7Mx6
QQvk1Cj8xWmUzRMhJMk7I5oUX/zkbJ5zBnGgOfep6MQv69NiTndo4S4w73feoy/AU9bYPDUnlf0Q
yc0fQ9JdK4on5B+cxX4TJkZw2nmVMJc7LS4HSA/JPel6cjwq2UJbxVPEWCARNU+QXzV4Df7Fa2nZ
Igv2mMucfUuBH1hxvncRRynB8IArjN8tMmB0f7dyugJr5cZ8MiJmYKkQISF2rBCvwhKt2NqQEZSR
b02wumHCLH91B3BbNzjBtk6DJihPKYTDBxbDyQXZ0hkj1waqmRqRQu/SeD6iEAD/hCntwDl/V4Sr
cLwZmPRuGOBIInmjc0ZRewz87mgniJozfFe8mzRkRtryTcSh6qBrFiMKR58C5HfUf6wvhsARpz8v
000uz0v9N6b/ly6R1supYBGG1pQhS3RippbAQqzKNG6omMrD0o/K3+nRTJFmdhgkJqvlyYlao766
9VF+aW9bj36jqFmJytoBPMoYMeAAPA4AezTRLUJ75xRUR5s1cLOd9wCkN9hNh2pLLczEC7ng8JKc
JC28R4HiKArN6/ptvhkq1to4V8ggkuzyD9Ch0bDmMwAerSZLRRXYwufyl7h3Qg/4cXfPeupnF40w
hq++4SDUSSVEra3aO02zRqV4DkZZRCMD9gToE/PRxkBC4U6HjSF/bUsLSywbg4QCCbAgX4UEqeP2
dgRiXG79keKGKllM6LTj1DBk5lDWE7mZxrWr7VEgViWAdmgKveRc442y0w0mulK3IuYMZrfYJGqs
2Kk6JpsUcKEE39S0fLmBRCDLYBZEIpjhxa1tGvq48bxF1Aj5Paxt0LZxKgXrwMvDftANpI+SLSkH
KFSoc30rnkABumSFlxRdFMvNnVI0eBiyz47xjSGLlpDW77DKefi4KwWo9pIb3cjpnoBZmUFtPKqc
aLUU07Vt2fB6KBqtBi7ks0NUJ8fhy82PlgDTEB16RDGZ6NTxXn+0PRJeH0sVmDyS/3fdwaZ7La41
bVujJzfWoIXkUXB+BE8BFIalH8JrXioLktBDcTKhnPuphEDDO97ygpdC0ZcuQbpoSTMNVCz9QIsD
fujnHh8tl2LwseNctyuLlFMyLTrnWV/9Kds+OzNGVFu6GLYSOrKrv0i7DrTq5ygf6VawfyO76yIB
e/ubn+omlH2Y/Z6nVXMrYUHG5TGA4txZfY6QNeLZANPjXUpDVxLCZ4FCHdN4G3U88kdL7umbLolp
6LancqnvZHeNyK0a4MIY22PVbG86Byvn1WpyzPlJ5NkeUnPnQFFvNPkO0t9EVRKEwafDFvzC7O+r
pvHXlvXGLDVBPAIOvvbR9hOnC4hQgJ3IqvrG2DZOnxYAIBtpFwv/ScCHRJQds98tqEPU6gLlh50B
lv2HOpddVwU05+Mx5kwmFU3dQih6e+wYYsXIawRxoJsxXWRzLUf7ude7TAHWS8Au8zOiQbgCYLhz
ZHLghRD9EMJv3AGIq0qGztjDyKYUuPhuTwpoREz9EajJgevoPlBCgokk56X88U00FS/NvCBtrJbj
EtZsyGzdSTHViPs8qHIOgefQM7AYkNaHEkaivWBOhMM6G3RrthvkVRhpI4hRTrLepwvAejn0m2fw
T8L/YLJX/gxBX0FbtrQ+bbuq8aPTQnxpjY2yKfbXNJZUDgkTNJcqFOrb8z4llmwcoDUlUcKhEtkR
LpV4ZH69DBlR6Z/kINpOHW2Vls8DDLhRXYgOGDr21wDIOoG2TsjXZ3gR7PnmBsDEcK9NFBKqvPmR
vp7U4+fdh2VJd/jl7fGxpr5gyDwsgd16WxK1tkwL3tf9qaxQ2im/YHoAhybN3h2TU0QjikyKWJ/L
QXyIC7bVL2Ac6zWEbaGdQ/sIV4kgixVg7EQ/CoN4jQIv3G64HDMV/frUDmxMRPBkYPjG477NBwiI
T6czopYtsthpGfZ7zrPUAX1nFBT6vsyvITr4vDXi66WZll1aKee/MJZGwfSboW23X21Ul2tnvlY4
yQtHD+tmNNeotdLYnvEkeZRVGZUeUqpoGV0cXq+lY55o8U/a0sKJWrogkcdDf9aiknwL36SLIROs
dKX5feA9Mx0rh08orxJRFlH3UkWIElmECGyjhiQrufitK2qNtCBifBuZPpyQdb12mFh8t2nemI9A
zNC0ZtVhFC2mXsf989IHvcE5j/cnj7vaQ4JqMaiN9Snk8wLbjoSwoLWLGn/L0AwmHF2CiP4TUq/2
AFmY2YUVL5IX9ceiwX/5ISiNpxj7CQw+PHeXZQ2aVFOI0lBLBASH/mTfu9DTcKqeB51W/kAkuTLQ
kEyM6651NT36qUymjJelAnZW0Y4EpveWjJMnk4q15oN9cxaaZ6jbsa00VuUVpX1BNLG1DUBANxny
HJlIlkN1k7VP3g8bEz2Hq4yDqhufIQDJx7bLsqmusnpAIPTeo/3ZqTzxmWYfxxkXBjdH4YsBMoTm
IuW4TX+c3my4hNHbnw96bIoTChKl8JTh/aEvCxjsS7libKvNQuGmOGGq9ZUh65jBeATPCTf72+DB
PVbVKdQWGJDkHIolasd2fMzp2HMU3vH0InIKsV/XoeaVGoNNd3Vn5Bz/chdAv/B/iSUgOf48Hcty
nKmVQidy64Y2uZLnQzZhPSBajIy91Hu8J2aWc6lNEpQHnMwts8dDOZQixT/C0DYfjCMxuzAANy2S
FwUjMZ0vpM7k9EmXo3faqGhwEoepm10pBiebt5CKBWbroTDYg5QNmDUDu+EQuzQnFo7xd931nQLW
sSWi6P2t5CQTcSkd0YQbLx/4VLB70dDzcphn7WgA17l30gR1w1cn0yI7iL3ZTiEkNpBRjLDJ+JCx
fSs+TZYn3JGL9rE+tF+ndcmR5pykvU+jwNQ8FFQWh0iSzySqMIJvOdzr4szi1ufaouHTY152iCcT
FCVzRVsPeEVUq+2Am+4ZeLoE9axAiTQfYxgoOZLd5w1mXRweDY8SRDCxc9hLtSQ1t5p+hlmYGxTC
4IDQhM+79Zpoa+wRFxQWrnQgwDKl9hI/244uS42G9VfrlgUcAGHZyQjIrlp/xkrnZL0R6TkkDhOc
/ongVepNV7ZX5QKiPyzhIjN6DQBimTHMUeuqSFKcEnYLxrwl5uYWT4GuRBed/8LEyZqpkAu5iwR5
vDwfhUbHFvt+M3W6NUVTVOtxoniEMtrRMUxucFqz4dxEDAYQJ4uc43s7W0UuPVqWtLu72COyNK23
UTp0dO8hinyLjPVRJJoKv+3REJmQJvLHiIwBoupkYltqvCb7CHDpWnHcHNld25714kTt4RmzFNWv
6/O9fZxu+oWFK1SkYCDwvy8PmbtBJSIbR03G4d1R2IEc/gIuyznlhW2OTAFYoyv0OtbIuCPPd5Qx
PAvbfNNV52MjoeEKtt8rfRIbtY8iEL+m5CTbmQk3WCeVMTSgRmmr6VLYiMazZ0ubQQkrky7DyWd/
Bfiy5Iz0XjLv75a0LAR+tZT41LJB85i8JZPeWxsFZkcAXtzN/Z7DjPJO6ePPXIVVvixWxrA+0X+e
kyMNRoVwNLbviUwWoQgQZlfg7Bow/kemXZQfYzPbatT+4cd0IAk022Gb+y93NS78LdmKJYGxdPcW
8TyJuhnsos78oUpxl/6D0NWiSyfxOoA54HJIbif2UUDdoB++MXjS6BY0BKNAIgglvHPNzmumcKIW
4wkeLck6+oqJtPp+CbxGAhhD8LQnCeKhnj5kmf7t1fm/NOdg99eAIsXV+B+vMmqWTxm+nOqMHxXs
agmmkA0bUD0RR1WJoSvSMDPs5HUYVvuyX2G+7uoG3eXHsOCan+TK2gXyQr54SLlIU7pEh755Q7/c
ogGCcDZvWy7ThSJVw2mFxerR55qgLK9JEIuh8vva1ezkf6ZMRt8Hbro3ZJagPO5N6ZFy1WuIHgmr
K5BKV1Fz0AFHeSlbmuTwlEOCNe+u4mzDBvVj7LCcbVzDrRV+JGf3g0FDiODzvZZc/DXhmx32BtXh
h0i0FYnSbNp9fknAPjDPgiIUsbLP8WKDqCcvs2wU8qubTKJy/gCxNuVUlom8lCJSG00DAhEdvf5I
6wYBS6PIe0fMMobAS6EEJ2/BzcqdJcgZf34PQImCJGR152Izcs4dmweZ+fuTwbvOFyunmIH2Hg2Z
q1F062/KyeAu+7QFR1Vo9i0s6pD3KtR1Gw4XfJZjt5PQ51scCy3p9UoUtRIKDANrN4v6DLMpsWF8
Fux1v/8m2W+q5FAx/3muLnroLnWCq7w0biKHuvqiyxjrFoVvscHazg4dSYG4gYmIcIRiMP8danYB
ITvuk46vUGIjKbLCqBft7ZvUGN+ah1k3zl57YtoXcppqPNUhO2ogPQ+37swkNc/GOwt22jvXfF9z
uoYaK6jP2A/D6zmh/rTO22obR8xrCHMFQnR2VDjtDsWfJ3N8iKQ+KLXJr9zYJoqTeRtoQKOtWag+
31J0yHBVC4fbKVPEG3LUcAPUMU5qAPDp10kFbHcp6Rp2RAfVzNHufy4mgQU3nQe9Om9pDHP3nqAX
pHsxn4QyHI3Q5vYOfUfJ8a07tcYEP7LvHEcsstEgBxdOilbokXrcNH+nxGe/Yku8Lwe0KXZ6JBKU
SaAORTfSVIfOzNapFs0uHqPiiL0iEegVkN8SGmOWhwSG6VigGH8C6rbQ1rOBFf0AK2nydviQYA5K
F/Oj/c/Z7Z5W1kvCG5tmA1l+4sMyD22jg30FNQ1yHmMBFExndpBLLlkxxNPQa1D3zXCxYObfvXOS
AtkJzS4jDSj/Ele4NIJIIB5Xc0prVLPwiQ9+3EKKNqzKhEuVo5wwknvIohJRGasvPUOebOymlLu7
2N9AdlIHyp+YqhxkGEMX1/nKK1fmIyIsCR0E3gy7ueUGbimntU1/5bibIoIxELRmP4gwUInFMXZF
MYkXIpkJ6vv6QIWmWo4hZOTpUNhJgpArYKWZOovaMNiU4sW6cbrRd0WwQ+5ll9IqJcpEDiL40M12
P68zAmGsv5CNXLmFFsOZLUvx5i5jqKLfO7v07oPSNGKNB7nB8J8L/vbS+dXg9+ilRsY/hg7qAp+l
u0FBgClMM5efZvytXaGd/gvmOQfyqp0pAFdLSlXGLl6+yw6rUf4N6zpl2nYOyeCTZS7XsKRcn7Qo
ibP7IsmE8ap5sBhH/pFJFiQbpBmsJ+nZ2bpmL9GWK57z5R7Ykz+hx2qnyopX33ePKKhe6x0FWNC5
2PfPWe/5k8rA959TvEBo++RO57XCE8NiOm67xis3teNw/ft+/Ox134N2TLWopdvu6FDGnoKRHfOP
ojRLh+3Ri5SKHsCd6AmQ4sCrTUs0QxreO0Ca2e+4znqSU4Hr6VrxwjwT2uCIEThsNNzkyRgpmivU
/QT98tjQCguh3nfIZKfbnBYoFn/lL3RHosIwMrfIzEirqOWucEoRv1UGc1EbjxoLjxmvQpdKMEX+
bcYoy61BshVAFlKa50ShCvxBj/D2N5hJF/1HrUrj/2HOz7F1pmyqXD0zSuAYRZYi7EYfTK33imSo
GY+VZK7gGy06K6GKlIIUBqOsq2HmPJWrQn2NT4/YqbiQhQOvYBzXHRWCQfgl2gFjgGjiSWdnGM5t
ZWlO2r7GvCFN252KEfn54NxbQf/wmoUfsE8yOEI/jN9j6R4KaaaGaTDbdbgJaiX0BBYQn9+RhkYY
wkdJXwlBz+SozkQgwyKNp0de+i8bG8PAyiGXALaFr9OCoTLyTIQRttcPgQFU2iTZk97ZT0oM2C8O
Hvx2XXmyx5dbZR63pjkU4dozl+vUPQNsuvvK/KTnGWhpfddRTYT7xOlQede7yOpahU5mxnHQez8D
fTTSzygLqnkh74p+O0w16wOMo5CZkb2WzwNYlLdYePV9O+G9XSIcXe55N4ZOuexEF07Va2F4/goB
MSwOTabV2LZEh6p6Z5wvV+GlYOX5vXjlOi2bE9wGb5ZKw0Pu4vY8VH+rqwTmmcptR9eF1bSzzv5Q
Gkz6yOhsYNYW0OH6b97m0xBhVolVKopQH/vwP03qvAerZAiFx5gAi97vqBM/LxFpCjFJQoJmg9Ty
AsdJHHnalPUL3rbdlNb6hHaIdRhs1gFdQcpH5UcnJVUnVQUl1VcI+oJyiSFG0tI25H1+Et8oWwZa
bhdkzA/dNaIZir3hbRQPMUzV/M/luO+oDAUowzCWq50fEE3VY/2U7QMzaIi7kX+RtHGm1EnmEFYx
dHyV/20Nl6DUm0b+0Pih46KNAZSBnQ5gRnCsmGoPDGiNyfQXZfKdG9fO8ZDFTU4ymA8rl1hrougV
Zqcx1AFEUtCqUIE+f4Frfs52C+n9kWa8G3HDpYUD/hock6Knoq6W8aTYG/MvOc98yObbnm6MKDAY
OELJbeE5DwH+yDzIG27HnwImn6Ze/05ju1hX0dZc+Ngd1BnmPtrGQ6AhN0XUCTaZpu8uQKBqCw8R
zw7MEJaabVuMcP6uvLNEJOqujcIYao417I5bELonD4FjRRRVRZFgNQy0AMV4JbM/v/XfyZyJndhW
809Fbxhe0a7mMqNCmKu6xzvDIkWxrNlH+U5Sq1YzTKuxzQICMN2UvCafPjrXg6VXXgLQajd5MwCU
MRomkugJEQ2UDkO8fMLY39QQma8qD7sQX6cBle2byWiH3PtWUW4jRfhrN+6ywbbtxAcAGi3U5Pon
9kGYD9eB+DuN8zf1NVOn7O60ymMrhGgsOOsNBeSKR6dK1aUR6O/FgTcEviz0t1OghYVSu2ymalqh
hceP1Up1mYs48/vuxUBTHt0REMKJem+YEmMH8twSDUS5LyJMhVUfEtn8gEKYo1FGIIkxAQkz8VPP
DuOo0BX5qCqbDYGNp3z5cKO8zj1R0liUdBI9t6ynqiSr2ef16lJ8yrc+q+9vnVimEvmYu/kv9KKM
6C4snq3V0/BQIhaozoq4UD3VUZoRMUixBaPUbFiV7oJAFUZoi1hi0CklTcYg2WMj7TjeH1ZeqhBP
7IVfTiPKLpR818LAMHQ8mSFNerb/Gon4yeDQqMc+4zBhRyLR6NsJ2SNHHupxcJuG6CGMrhtKy8MG
ytfiIKeimrWgH6Sl3ZI+SmKm3iHkz0057VWjUZpbDnpYuBC5+ID4vNMLO6wC6rT9nASPOU9NviA6
kSd67eZeRYImrUMXXqO7v/rbeSAsDGxTMq0fOjCCAPyCg3nkOlVk2jTMS/Vk+536MgX2x95lGcWe
Fnyj+2qt3drAqOI8gC9UvjWwTifOSGCqaQwJH0q7C/MAR9k21Pt7BhJ+1P30U4qyFIFbPZSr37s9
lqId/ypUxZ8X0hi+yjwDcgA7iKN5j9E/KtITXRbNYuCFNZxp9CqwD68T1ZHrC/DTWi7xEbET3bpr
kwabnWkDhzrP5UVCXWzGQ/hp2yB+b8xl+2spuOn0aDLcUoDA0rllKIgK1gbgOsKOeKX45l4xD4jC
olZdy1bgztnIse16coMw5NCbm3hG0AtqEESKiaqhevNey8XHZyfxp0im0Xdfr2qLrb3SHdFE6jbf
4xgMaulO3ODjO4GploSGzjD6bPqvYUPbPRAfccWCJmnvZmeYV/kwc1M8h7h6q2RRLxckRA0zfMzS
yWHew2PkUq7oi1UHtbtPTk4bO+wANx/25H9jG7ogau/jZ+pcX2WusB655OdUI4oG15t81rLMMVpb
asvVgr7miKl/xf4eUHZZSojXoNFFRpybF6NKIA6gEsLvS5Zx0NsbRIZz1iSTFW/mZASgS6Tma1UC
G8lID5hVFfB1Dzai2vwhMSz9ffFFITcks6RfRuX9oxd+G5MDHiWnLoPKQ8zPoAualnZ5grImkutp
ZdosKMeOvuESmmJIInw9nIQJeABjXwb5TErLr1SoVE8kSH2QqK6bOYqHYHUqCyLzQ9IrfiDIX8rn
biGwtVfyBmOhUpxLwvJgYdOBCsS30LegrExObAvi9mDebDiLYpR5UgCiKWSpIWoK9CHkc3/eLtf7
cGQfABjdtR3E/27SnZ/GgVTBxYhKBcmvwju1jYbuPOfS7KIcYHI+l5mqY63OHHZWNcR7Ci9ufsAV
NgubrIKJwcnAYM8fmYrLdQLigUaqqBxurK8bBONZ4cLVYGz+sMPFOmuyJ/UiBqIjkHH1BATXvS3t
Fv6chuUYlerHVvGaEylR14mm/3mKzgJ7VwDBU/mBM9nUJEoA/6sj40wknT/0h7Nl/NpEcupSlyhZ
/pvRpX/L0cJyW6ZGZRjvFSK7hlxVlN8Vmf0OTKI69a1a4eflogJ2xNhMflDGqdzu3COd1NPy6NO+
EnbXZm0Vu95qYtKcsDBFEmschQVMl3F2/yJc0UTWHnf603Ex9ZjtwLuPyMCywcNJDf/eMD4qol+5
UIYZhcgJlpTXKogdFwex3AavxvxTTM7Omx7PwsOuo1FaOx/l6WpA0or6LPhL9Lhhh95gx8tIXKO4
umcv7MRPi+eUADICYZJ15MgLxeoVCasO1v3AkCOLiOMsdCYZBCqxKnUrvVSDswFNwgs/8YA9HQy4
Sv5ycYONGdjQ1gvvohfRYglvE+px+sAhr3+d0HU9BSKTHgOX/yxZJQ+366uRCzIDoWE4E0G5lwBE
BMtSoTyQn/4F0V1pEd/kHKFVFXwMhEHexHXDwLCBOa/C7ichxKFeX4pwEeVnmCbDQryrRmK7nRk/
EmwR44Duuu8qbJ7iXjVMwnki1Bz0ya/5Ohet2aRt+D4UltTxOc9+IbndGU7gr6EidknmxRjLpK+c
PdMxaL52eC1j30Heji1P4zKJAVV36SkT+lu2eqkDNzRatJWFQCO6ocx5teLbXM6V8tsN+o9woUB0
Xv/WVBeizO95ndxYe1Fq3DwOyJq7b4wrxACKhi6zmM1MqfIsegvBq9FP+xa81sR7IGFNlseCoi6v
yZOFwHDjXu3kJV2duFRBUQL7ZVlrwdGtH/42lMyWglWf13bQ8DSRR+xLGsgrtRfVK/1872bjJSK1
UKj/5Jbsn0E+T2EYKRb2yyylH/vz3UkUjmhk49Wa8i8+gFKfzGn/rjfYTNB+/uhLGMfhidhFHXwY
fnfJ4gS1JyNqy+aJnmDG21o7tzGW2VGOxwPPoZInxkqXuyAbui7+RtZW+fj7qoFPRJfwk1qPGPQ+
EeR4ZBKkni/d8iNWd/liPLGhbkz5i1yGUJz+q43aDznbgRWVpdKlPppg1sEdUnUXYvUZtt2VcG6m
BPqHOqK293WQnnZfNVdi65O0IiM4MLEfhtSWts5zG/E5lOCgNuwQe7uuRfvhZPAyidmZxAVHNUvc
W0bQrjCaTH4GssUNTiDIjTRv1vEAAyqc9JAUA8rHMdiV1jVTVaYVasZ+YTHqROxhfgcdQaX3By7D
Ax9vmUyFnwzUqFptMcJzOlpkoLYuc/db7Elftu1tulo+TVjPcaeerHg41GySDI1CJoOGogDXhYyZ
kevAKsQNUYurEjCC3PT8greISDc+hqAlwG26vCe7Qz7yyKMkDu3BBSgMUHZpmd7gBsKkFMtIlO1l
o9L8M+9uVrpLsSf00V8QgAXtTS8gIogJmeBjVB88kC4MgzI+eJxGOLqaVtAV+b0LKKnY7XBsPtvx
Yau4tKzjaj3Rwc7Des8f/6V99RCxjd6PeYWF4DhJ/i9i3uBlid370JlWSM9PtSP7rJihVdmsgd4n
yfkiRgHdHpdSuGNOz45r69QwwyPIhOXWfAa560RsVSu6uZk6FQkQLYAmtTHWzNlhdImEx/Eeei2A
I6HIyJsaNJticVixPw+kO8Tw1nzDuxxKtRsT6fuAnP+MxI7TEhLRuXNZdvROqt14hIV/+PpxuzFW
6oAIO+02S+GS4u6J81WH4roCUyZ6OHoqDP+xEYZ7/O9UTEk9vUaSyG1jogf+g4/4lGvkEyJirK+6
axWIvjjbBlBp69pOjCMtF/UZvstF5YQhIihKoD6BtjdOfh/IG9av0VIs2Uw8JwZ04eDq6TWvbqI7
9N2gF+yBdmiTFCskVozJ3a1Lfoxdoc+wDg450uwn0hDqxtuXGnHVLydWa7X2oZV4FoGQEfSnbShT
1gzt2LvXKc5DGcq6/vI7oFdbKf2WNnCYQTu1U/sYwEpBi4l5hBC3zvNlHZ7KprOzq6TXv6YppsC8
+6J4JDufrjWxBdkCcEggMMUxYbReMitW4GLnoyVNUS4bVaK0TW5JUXeyceKCxEzhTl/DgdBGU3Uw
nkZF2zSzlS9Uf4TXWApborp8Afbp34SC0cYLqbLjTlhhZJ8C3jNdlHW4yJopqeM1VYTg0n89N0JA
AgogHb+PYSIS6Wt1ti66cho070pXIdN7hSiRzGDPAQWLhc0B8QYHd/Qx3Bnp1H/VBWA0rnU7TA1k
3P1wmLyKd8Sg7ZG2Q5zh51/nb8nTYmikWrKDDK1Ju8LVMIWVJcFGT1L3IasgdGnlhblb2PSnSNrW
wReYyRi8O3b1eneauSoorZ2mkMkYsEKZ76EDs6W1OGaeL938B06YUw2lKALzXrfg27xu3LDOBQdl
pZBWshkIPfimLSDz9BixyevtcNvovU095BtSlcWIXhG82BKPKlzp0k+qchbiSMTTXhEwZ/2hWbQq
S7ZD9lXoOKXgj5OmHJYiVzax1+gFfp0VqfbcAfd5jLD4CRG/FOWOn9wJrOrP7NMazf1NlQwXQ7B4
x8KXpAKHe/jBA4lnAvF9XMJee3gCGtsaozyiL7egfyQ8Xxpea6ygFR9Cl9pH/dXWWaGhfO51A75i
+c2ZWr3AeOEhGAkiQSD+wy8ktgMrYBPoo3iWPEDAEiKWvp1lQWyQSn2J9trEwCjskUA5TOOmp7Aq
nQqr7GYeq2q66eZzjFMcELM4CKJTGznyxmjx7yNDzEKh95AnyxJVR/s38v+/N2EaEanDl2YQnGNZ
7Nx3v6EW3xY+c1z8sQXsdalaiqIPfHqI0MLTURL83C4GG5hBk4uv2FTFeSKa5pztu246lyf+ox8F
Pg5qKgMUYyAFm8kKcJsmZhUx5P494IiW7thvWXO1qW0p9mdSm+vaS+fIvIAfzlXud75OIRTbdQKn
4s0eDnm37oTSgmzJGzv3OxhvV6f8fuLZIKomDKGgk6U9uvDF1NJj2rFgU6E+ouDzmhIgJDiB2N8f
UYp7tlnGlzTOD3ioo+aRGLUwHw38k9HXTZvUxnumAsXDWztYZk/1XXSnv3AtaGLNE3divWYNygy9
VB5LkI929pEXOthcvyz2JcGQu4YhwW7F6KiCNR5bXXBAY/n0nqv769Dg432mORm45zzh4EkgA09u
jKVjxZEUn5CUCi1UjkhBNKR68vuvc5HMdOgEm4ASVJFJIAnKhH3s6v7dyMC7eFReV6jP+5xBkqjV
TGymAeTBCjEIP7oqn4PN0miWiww8cKRXqSdCMn7+4P2wHenZVs/vOwLqaGwdkEP2P4wwM+xO7tFj
vR+JRFyx69wjo1xTcC7AA6lVrOKygPXJf7/6dUusrqZF+7Yh8+ng6zQhog4z5e0jRvPRduzEu4Tk
PtJmY7oCI7uWiskBLdoZapDEhRAIAjqOX6iT6iMLR/oarFBlnKNVRmkSBdUr8Pmw+Q9A5iE7yWa4
VxNrFWvf72mqa6Vu3j8V8Fb6L+ci2Rqjtezi0RYcIu7mtyXnCzkSs8d39UXuAWRcR0P5E0xx8SES
hVcZXysLTidlH9SSna8lEL3IWb/S02vuuoMsD4ErneGp+lKUz0xBqVcgjAmzY7Pddo2vFz8G7D2b
mNagwpKP78zhx6DPQNp36dX/PJPFAgXynRuy58mVqtxZyvjQX82z6HO/nGn0CJAM3xjPiFyXiZoy
EC9dl4UNA3/yQ5iYtdsiD+PaEjXJN9iFFmxtXRUHeuz+R3N2aVfeXvByGDQVghQkn9L2BVspCj4N
bnqO5VQDJ9qRRdrsslwLexpIu3aufhNuihbrnH7DzNa6OH6P1fcQrUdVq8K4jNpy4Xd3av5UY4Ks
J1DGmtR14mMJupDpbgh7j+vbHpbuo7JQY07srvCxmYGgMK/7N7POBI/39RwZ8M54WZaFJt+RHv9w
EGbW7kW2BmAjr02yeFBQMpw9H9beaTcZxvUvxWlUwnIIl4nmF0CSeZMwXnvA+bujbDLXMHZIcA6P
F8d/2XFvUBT0cLf2bYWqZzqmbY9gVB3TbkATdW78+LbKu/e012acqM0NTiAEsAqxPtMNEnVDEd6P
/rpw36K2kZ1P6h929t4n19AnlCSBrmVtn8bnLUZxM6T13rIfLxQSPkgRoR9GanvCe4DeVnkMZds2
jmkhoISXHpVGdnZ2yIRnxNVn636jqvYAreJ2LIwo3HVekQHbVBJzm/y5Yg1Ddj6B4+HDcojWhJt+
I+GWcJNrFXZGa9L4YpZT8uIRZCpWTGTJh6ZpL5DFnIUcQTSCaravKjvIO0B232fFCdhAo6n5Xk/f
2e6bzse01v4YXmWXkQ10BDjdwK5yV4dl/QcrbKvPFK71kslD4/2yf2Q10R48MAWlaTw3mkKc7BTA
9HoieP4bdfz8V0c6RWndc6KGX4UUY0YhKQxilKIkZ5OpYQIyQbL4amSUti9EhqLSiAbQ6WSNWA9v
G4QqA/F8Az0WWdPT+4yxMchYVTV9oFqQzs5N9jtXcykqXPZ22v2P/PkDi4HJNEHetd4ZQzm0kMPk
F3fVt36tFo52W+NeI+/ZG+zgFTH0d3tOTuiAWICKoQ4IcCMpN2N0AMEz+4gkJ2XOBgtZ+8j/oXU/
bjnWTYn2xtzrrqEWaI6QkwsFfPSuanhSqY4SaAHQLmYinXp5P9cYJFuqH+D0gOQAMX1mEpsvNyrN
7T0dzQi8mlaykaOhfXGDMmQL93aw19d63pA7kr5jmINii9CbUH1b5mQyMpPa2qP+/rEJKPCMioJH
+ENm2ko++aP+q3T0KbY+uPPNaZEj+Iy6er/gy+yKCOtSFAKdFW98CTYddQaktRWEO/TW9sDMCSbl
Jbqy2iOZtRk8qtc56DFcXZXzuQJBnOEMbiLQKs7x+DEFZwpe4HheLfQe2hn5aIxFD9Fy1/A2HcDT
YO4r8eMlYOgzWydMehuxyN7uOR1K6vP7spUa4i5ip+ZGZqDPKLrpB0yg4XNT86nrWhyRLugsHQSh
ZVsoOsHG0Ex/bFB/fxDuzhiqZq6rplYInHd4DomOYrSnDS7C+CM/wrQbisT7Y30Z9QE05xVCtPoV
5KuaY6h57P6Fg7yfUn6kqlZxCtRu84qcU4CdFnezf6F83HhEgFPD8USZX7kmezlKuU8uAzqEid1a
MiCW+zHP0wjLVaSsOCJLVHNbGHrZU77ZuUcLf+/nK3Ed3lTsTiQbUUy0z5X8quBNlfbO29X3es1y
DxJEAfqpps4YLLTFBj3DB/PYDgK4eG2NbCOtwdAf94LwlkLygDNL9ACMyua0MVof4KC9HfscyENa
BKFF1gAsgOxPNtX2rPXIWv04A04p1enVfCNI992I9CxtsOjJX3NTDn6sYn9os5gQSVr3YWqGJk+c
J54qO1rl3k7zq5cD6T7zRkohb5Z0UcY0hYhbseBFdxP4pNZ5sFYnU+7clBUWBwSquFgFwfPC6Iy/
Fo2qseMYttqlkA0sRkGWInzBbMUusCPsg/ZQYdVS3FK2+aOzl31WP8iKITxAeDJYWQ38MUOBhaNt
WsSbEuAdp5phfrD/1OeOx/3Zz3BSGEo4Dzs5For6COtaIBNyjjQUY5yAHtQuubPn9LU32SvicOb7
Vf40KHDxRaABGwiFyMTcJzuURCVSzmRam4SUd3YtisddDxXDLHEkAnr7ybt2lS2E+F/l6juS1ZAT
R//SRzmnY3t+KPGj+wnZXZU8GS6LhmtDbZF4ecod4KJ748gIG7FcjMyGspfBhbWfSodLuV17oLY/
P4pRCK0tNTSzTzXtQ7eFdoFiKFP87QdP27lbdlYXEEpuNCW8+V3Ak/lzsGvV5eKUoaOV0p2GGSng
HpIn/8w+7XxvVqkaVquWjxcV+UTmPS3cIFgoPuJHO3X/59UDFradP+qkU+Bon0QmzAfPFKPB1HOu
mgT8lzOhgkokOnNwZCYqOMnaT8cxQBRKxLU+/vO6IKUgwHu4wDprAir0VBaw0Jg4XtuGzoJhiccy
NekgrG647LpdBYL1bN57AYBuY7MayfZ3pDqKf6bK6cVtZZ4BWxSElSUKbE2CMLj5XDlTF6VxaGfF
SavGOAH5GS2isPZc/nZWswWHnbHCn9IGu4hL68EFieG4s7BGPjaEeb6cNZhRJmcZVRqeD+HLWsye
2tnkuQi2JvkWCKM5WdtM5i4kiwX2W//FPp0k7zHansvgDCqkQZwxCW/TgcpHSa8Z9xSBEZy/CLjU
gWCxsP96BqHIAmC/jYbOfyrR9XoAEK84EgzbsBrSN/R/b2de4s5tDJyZfovLNs5bXxS/OILIAAcR
w360ZihBdAw1zABLcaQYprTAk+CCQBdxnN6zC/00gdAVNRiamTtpjipyHVg25Em6WoYOvoVgHQWj
jk3d/S5Lb2ofFi8WcSO8j82FbGnSlFPm/rmR7KQDk1u5RZdEagGZy5Bz7LYoqwGFc4YVoobRTO0P
ERcD1Qud4anr/R0F8uuGyLbl5b8nq1g0P0qN7a+FtuftCqcnn5HWJ8hUQQBEQilAmCM0G841XAuI
XNd53HaieqrR0xaP9Zu2Y8J3rQ27ZfkwSFW7Fnx4Gp1MIww1oYfkLptXBg4VBLdKikxzWqjco8/3
RHrrBcpfqGp9reRfaFSDCteR5JDl3kbP18w9w/Sfnd/iobjhKcXgzcMvF0VzTf5tHLKlppVYWG4r
GVHW6XWJrUGJ5rjCxNt8NH0v777unSQSEmgXlnrJRpSFMMkwTlksvxOE4vjGz1q78SdO0iwY2J3u
4ziRqcStGq+OgDRTk7/uAMCkwd4gyeb2Y08U6kuvRwJbTp17DV98cBRSLkiuj1aA9AzUNg5tYDAZ
CKpNdghmcgoqfq0Y4U8sY7BnH98GbECF+byU31DnclQhCrhHrF9ERE0kVLLpkH/d14qw/6HnyxJW
JYhxBkJRchABuT8bERpwrxdcolqSx3JhAMX2GN9rASC+WwWHPMKhFxVl4IhoSASR8GcDlQloQUnB
blD5wXx+be4mXuv9uPKGQWZjArqh4OWOtcuJuSS1oVbFLbcvDUCSyQc9s/qIJ0/ZQlBWwH0SWeJE
IowME9VN0ffmOXqf2pYPsq0bRHhih3pcyI/Ejuxpz8UF9NMOpoifS1UdoAWooC2mG3URtlovrc7t
SkxeXGGsPDpx7Gn2lqqOjORTK/RaHxfzJxOWJIXmdMFA5QWHw7xZLZIonAo/IcejtpaWmqPA+waa
fmnD81DIV25JunhTrc4u22TnBprZ1HeKqJMe9poB96BfS1Kp1c880jpjqRDGfUvqOVXEmQ4y4PEH
Qwq05DIFV6XaQWFSWXnOi/eU1Qknnm1pbiGOfqZeu5/4H2iUlFJhaMb4yOwHAC+PuIizANamhACF
y3ieAw7LPBwZOJqMfSD8G9WbdNwWxetoPKYOiER8mfXlsvcrM1c2lplX7hbPdUa6xkTbkM5Ca2A5
2fq0epI2sEojXPXqk6p3+kcNFiVNnJAkgwyifWc2K9716NZdXPZU+SuQOjlTM6u/jNzNl/NOnanO
P6c2dB/PC9zZaer7BltsCN2wDrUNYXZWSpQaliEaM/yRYAb4szDcCFdkxZ3fiOUO2jbGMU1X3HQY
s4wNtgzSUJ7zuhaacke/Yn7y6xB4g2o4+Gy8P5rhHejALjGUwZORyAtGW9HTqyXsXg5VXKDYyDse
RQPxbp/VD5bo4iEEmlRaKfHvUzhcFwAVK4dI0WMXfMzh9XW3kVlBYL6gT42KG9x0Zk45IHcj8AJw
QPkzcofdhTVdW0nFNGWsZURi8IBlF4ctSI64eWEF+QeOe1lrC+MSux4gOYXN6My0j3zK0+pe/Eui
U7JwBmtG3C1rG9RhuC5BrmpC6XcyH2UGBewhdWjvPKFUyKsNu9EG3gN0n6n6n1XTx4ZKHUZJKAYm
YTm/ZwQDV+r402IPXHtfWlsI78iNxPjYGIV1yGa5IqjDs62g7TMy/CD3Z2mKRNCZqQcbPx4shfD/
Ujbb7pJ9i1Hr2eOtJUTRJXPeswTQAYawTZhLBOdiQbsHVQcAqOhmhVsyPIC+OEcMlKoZpqoPYi9M
j2C5PHN1X0TWqqmzk9AB8zFcbF4kRXzVqJw318rB1Hr16RLYtrhXMmsuQwli8Xp1aj7GrZ1sT+4U
Fwz4kMrk71EA5D7m95Iy8n+0qRcb/+KOVChQgee9MZUCaGu9DVGn657j900WDTZ4z2+0ASoAo7at
QDJqnTUQohpfbOs/cZTOSbq2VaSSguPwXTqtT3gUwAfob3cQVnKjnNqLLthEIZPLXzFq4AT/Kj4Y
2JFCIvaxHWglZdFGZnp1xpSJ9fpl5neUSLsvbKbGDm93Mut2culoM73pCNDwGxP9CA0pTGpqq6Rc
Rewf/BhfJTWKKLkEihxf1ZEaWUBOITDXBom31xu27NvDQk1WhQos1mcx+fiBhN1z86QFztlfb5kb
+vRPFgTA4jl9IDsuCJrrUOmZV2+hfZ2Kc/ej4VN1Yl9N4NbW/T1tCfDJDL+XxOUdgVT/0qwj4xc2
Ob+FYcM07TrxvXX/pBvc6YuXCdCO3BgTlB+bUSJ3IbrQcg8x3mEqJBZ5c/2DX8eDEW4ew4L19dCx
0lGIPNkkchnqWIY7CMzPRWa2vQKzXjKejxcDgC8CMknCRPjZIH9dPMeNdAKItVxt81eh3aiNXn/0
brNEIzKQ1P48fS8X8nZuzEOU39h9m4IbKiIqtu2Fg/dHJ9afOVXNSOYIYG8rcDX4h/nOqXNthw74
7teJGDxn8uKcwfrtzRhWaO9qY72EIHOWWUAe0+PMkuXtBTFUaMQsGYuYpLGt5euSFRUjltR0zdc0
xBEKN9+b0gvNUQEuQhhWrKM1t1pAqFHYZxyMgiyjLx4if45R3hP52pY1s/+0fKYDrAkQpmHMN11h
Fh0yIGSDLnWzjBsnaora5TQVqGo5DjoqrJnQEuYSRxoQ5Xkpcmo2HLsO7Hkij3O6kjYR8jiNZXzk
OQOOaaU7Z/R9lKIygRw8DE6OSfz5/TYEtmZcqSzBCdKlfJK4uZ1O5dc9n/JBZS2KflaS06SG5idy
VgwSGsZlQFU2QaCV8oRjiSqL92p5tcxOLKkXCEFTX0TFKur9ZpdURQL8hkMqN798U0qil/872Sdh
vzoXEGi5aTHxlakfi4RQa2ZweKL3M7S7jCkDTvPtiCztkLOu/N47TDfO2jXZYaztf+TIRleoj/fa
3BV/X+zLmR1bohb+wDU5ppKoQrIErVqpADMiUMqa7TAvlI1391KsXd6yMnzGWKwPtn3+BGJIuNLv
FCsW4u8u5zORrWnCZjJvUA0TmNJWqKqUFr3tUJuQdLovYo8ejkpxKvl85tYXSiBtt39PfqnqHihP
FGniLe/drNmyGhom3l+2aenzwtDEWCJ9cOp5dWm1LyZRC4FjZEBNuOcUgyKCbER/aiogt/vMdW6n
bfP2I4Tp9PVg/aa4OzKeefauygrG0ibtUGJnGdGNBoNEGOQGSCqZcmYzg3dhHaDQLrLMriaDsgk9
SUE9pl7gQKp70vgeuJuBmzfzZZm/7qjXlNgFyxvjKW0xxym0Aavwj9IeUpzLktGAB3W/K+mpMxL+
Y/DrQMqSg9QdL7P/wChun8X3CZY0/1OUkojcp2gpKCS88uoGqTZfpsQkbwMHpUhLMnyD4xt+MDHb
LsECOvcx8PJbPXpARx2urDhQvKbI/4gY7WMR7Wk6zOJ1cFie8QRXDbo1Wps4jTb6QKY5kaU0rm+/
xjQCfjjfzdbdlmGjZqqbZSTD9iDpEIic8khpu8KvrZwoOVOjU6ClbFak9RHHgD9ITW/T/fCF98TO
8aZfspgLNpyBO+b0arZkShw2eq8hS9WsvUGnUdZTOaao/aLRKzubEbaoq8FP7/djggSfbY2M70dw
DrabRmF6MDC2WAPCKHEJ6ckyQJEknVLjvLccwBy92DzlwhD8NUSBJKL2oo2AAt5AUjtKY4w3xKSE
bmQXcUTPMPCOaWmZLcjVLz907lola7V2DuMk7JM+fvp51LgI5vTzfgdY+N/h19ks+MB9ykrzzP+6
WxIpE0iCWMN3ySUXNLaGiO4bQrQAOB8kbrvDQ85UgdA9PMm08iyPDwBkfWUaOm7JzmyhpiQ7uqZr
rRXmGyRqXW6zlwggBUejxv2YzIw/kfWdOcG8MYiU0hqdc81w2sKgqPONUFu8MNQ43uDgJsim73U5
aYvlFLhO2vxByeAdvMvbLBwPEKpCGxdo5MfyaOg+tzNw/BC8TSWwPAFjpSyxyNP4fptlPe65X0LP
s2Oocs//Luz9Q8syMo3GWbNEnB8ThCjoDB+vkJfskZe0LWqiqLaP1xecX7eeiekRpwLQuya8Vmqt
impKKNaVox2jmPqrLSLV2xV2nXN0Id7mO+xzj+EMNWhB2yXdg8HnaXD21CSxkV7jC3isfW4hPWoX
2NBb8nc7JGIx3J4DLYYnhuSyi5fINGzDSxJnCvQmZcFqufv+o9E7j4y8YsPLi5ZbUtGTY4sbhAS6
JB89sIGpUNw+0oiqTH7vqV9UfQTW+DyVSE5lETbKe1nj40jKCBzqy8Ie9xlh+Ha2aD5m2I0Lo6rX
ZUkoPZzcwkW6Ef50HTu6II+QnyO+gcuhG86Yr6x3dC6KskgwdQo8m+DF7VbTPHz6yf2lEABFfCn1
AXaUzGTj9fJ8yvH5xr3SnSk6XYSJ4mTfbl+NHAJ9OxctId/iOjIgBfC9BIagnsSqhrBJ5d5vEvSz
24mGuzdsUE6b8c8IxF2+ajvre5dw1LAEx3nrngTfwobCdB24EUet2ukD965gCc+DLDlizQ1WRKkg
mchId4ubaq05B/hfo1k73Kxbw35K28qb+elFosQF1h+aHkC+jVerZ+AjFRCSj+0Qb+dikl+XRtiG
OG0odPMNw6jMb0eglGPdGyRTImV4jEoCdCA4zMaubdOi1w2C+HA4MSvR7D4MlhSIjMOOZcbNBhvT
P0LTsa0ZzHgIOl0ksDbPxNNkN4MZtsWCeyY0s/osRLOlFzIAgbN/6hato3VqjVWr/V5/V+T29jLh
69j/wmLQICJ9OPtf+xfpGdxBu5JBFrieisYfrlqwIejj16zA7QZlQesBGzD2lH3m/4fL6FhQNYsm
/wFbI1ilQOjnZWoZ/ZpRVnmx2FzgxuWta9f0BGkqYVg1ZHpY+1Ln8WLpa28lj7KEZ5RLhGqi/Uri
ZoV4mdqgyYJSw2siv/BQjuvDbaw0iXFnsVJO2DESIHWpliTrk0G17FSE49pyZt68Yu5zOIabDSlZ
TjOBGcsaIR2zo9ipiJKtoG449QULUbKelbRrOq8CqZzoMrmoN3lGa2A/SXt6ignmzyQCy0rqtyU9
4cGuIsISfvPSf4xsvJJFYjI8qjD3uONxSUydb54QZt+uhiQiei5pRQB+um7tULX2Azi04sCeKMK7
IcmYTlt9Gw8+E59kITsQPt7mkQ1lwlEfiy1FcXAp4Q61wP6wwdxsLJmSiAxaF/XxE13CNj0zHgwH
0g4BEOKeZkSeU/nsypRnLs5vKMh6aHMnODLSIYNeMg8HLF/Eh8HGddchiCwihhB8qJBLqr1AsHjF
WTMFHj7WpspiivElW5xrDVRuzT8D/QQUJCYmBoH+yQjsat3TZYtNOt8I6/tOc0RVo1fmhKnh78p4
WZHmV3PSzSSyB7GILPGTlJmSZ156I7yXXrCMuutldS+SSNeQp9PLip4xzVo7bOx72c5fRgBO5fv9
s8yCNyQ+XZFHf3deWQnOx6E2gr77I1G5mRAsLjUGOHoqLv7sZIAH34Gsf/zw5k8yBAI+qVgnn/5W
y+g+Nv432wzRsiyUqFDwOxz3J2dx0F8yEtPWG/5KyIiEip7Dodnf6JYtThxg4lINeKkClEym+1LE
KrtJOChgiJ/6bh7Jij9rvYHR28hcnHx/KF2eBn2MHAhp9X8m1b5wiar7Rye9IyhG4UFNFe/Er6qP
I9Ir0Mpm8ynkKRFuWvH8MKSFo8QX8wiFOLJC3Jeh9/OcrA3HOEDTu+AjTElznULN1VTTPex+VKsr
DrecC6fRoB9m6mhLbpbKkA2Mcnp+ugA339iUqAc/opyCKGOnalfO10VP217FliZg9F5gB37/Zl/r
0tYVTot+2S9Q+mq/kuVFXbc0F3c6t49uzkvlSWTncApDwRsEtrFNA7DNw5kI7Pjmc/8c3dq/CqvN
2xwsH4kkt/cH4zjwr2q4GvVyV9podGFf61bXO5dpz/f8+UkvSlPEKL18ReUkrvvmexYB/jB/G3ZB
X9babj+ieXGqQJpY4LeXwZnCP7eF/O85iFSSLXPnWOfVk/jEtC6d/WrgYt8Z7mIghlYD77LvjWXZ
aI91u+7BUnSHiAI82ISkC4SDbFVSDPvHAg5tWwRivzZV0kAI7/GJdGAmXpLXjyV+Z6fVOaFCyg3a
HSSxecFweplRbvZaQ2Asm3Uk3C/U1qHhmj32nsq/auGIN4DjvtJiV1Gx4T9xubMj5mzQal6U0RBQ
KhNpSpITZWqkpxIdPrtTcHRcK/Wh1Y4scIGHNBVORqB5yjpm0LcD2BM4TqUkfepHthaXknmH0Pdd
1nnvrIu0HDBED3gwPcGp0ZA5vjCSJ/kQUmOtdrP+cVBKr9ZL9g2A0Tjje7OeHQZAd24WmssnpqFU
tEOe6MXBF/VARrANX33dISz/BeY0G/uPzFVc4GjAeHmH34dYoFAmVCyHgHMCa8udY/H21we1rm6i
SO9HXY4fQU+HLnrLrbVwD9orD7ZAVWqJqmZLIj9DIeoShDosf/t8tG8+2xxYXTBJ+9rL22QWiXS/
VKOdGfw7LmSBNiyh6CIsI0I0VCS9wmFwzoV8mRQQVKBDLvHtr6ma8uj8CdZkV2/AUiovXNE50rZt
Mi1xZSrnngKeBptDjkiR8nO9URV/wdOgZY48MZlZGoVldOHFcrCfBGZKcwKkUM2eseslF42Q/bXA
sMM8D3IUfhtmL7VTP7XkeQxzByqnWgn/0x2nMS9ow6HsuQo48UpkUCLyyH1ByuRqzi1uArxFik4Q
+wfBaTlz99zq/AYi4k8Hnc9s1qu5F2xxjcDmTAmsoq1z1E3uU+hNHltfMZsYNhC/x3uXPBybzv2+
A8YUEasQteLyKZ3tjhk6xGDFN/PZ7xOh1uDrWzC9SaP6acLynnWEHAPUNRveK6G+Dq9LqIwkHXQK
l7LDL5sCq0UV6M9iwcN+C8FSyIGcB+Kzk7ZjibxFa6UG2zfi3Hvnbeex6H31f5byBzYICn4gqAfS
ASGDR9PSJIkGdsF1hq/ZjSlmrwqe1JxdTHYmFQzAalb67CcwfNjd21/fJs9KDEqNACISs/8UUJoT
8KSht6RwJmAwnHoWVpD+UbWyjUXLWb3p60VGoy/UkMB6/23XkKmvYDi4Lo+vuKymrEDazY4lJ1BV
sogU8AY6qEBcjjF/+NSySjuSD7TxeAAl/PL/mcKUhdc1y/HEslCtRX4zOfc+D+446gqzEUOjZaWz
ioY5xhf1dm/AmTpfP2ROcU/uNVDWw2JUPm64TY1KEvaqxl9QRXrYPogrRT4WllwnmCR7gQFmKgcL
vFWHeGoEuogbk16Xg6tLYwluW9ZpYaMg8jq+exF+ELuBoZVssdK6VsxqEDlCRs+S+IdrN1IpS6vy
lH+46lJ4I1p0at1j2LjII96MDVAUGavuLcm7pnBl8VovBdirkI3ZWq+j5Si3K1HuYj3JKC/KSI+I
1ld2/2wrCWL5RSMd9zxpxWeHIF+PLJctH1SZfmPR1dh8wFHT5Gd44rsokm6op6e8UWljK+m8oy6e
IsXL5zTpBvyd7mB6OgPIxHk+5A/pi6HK37i08st703eSOLSWXxMS3euYJYAf3MbZs3L6tM0AMV+j
mlaU1i7d0F9wq0GJF2WYsDkmzxEmE0QL0DIeRtBIcKp1AQ08aqTSLwJN5ScGeD8B7iJYmOM1dATC
nijvPZPkci3T8eHfLxGZ6mOjQKBWyP53QfN+BqeVWYq3RCIuxCaRyUPw3kBu89OkL9lDsUwNNnb+
ZBUksk/BHVYtJ+qNs02cakpmEFKfv4F89XuFZHlVF219z/LRRCE8WM89LDvuYYShL5ImMt7qisQT
V2VyX7mRP4Xb6Al41ZpybfcFUIul+w4J8/q7TlUyZ3QZlzYj3VaBmFJ8l9UQ7iIoC6Ygfuemom2Q
ifamYwdouF3Jm5snRLyUBmRvApMe4RpPeEcHmTxOHe532mIJZLPdU1xKGSQZsLBA0+RE666U1hgG
BtHtHhLX/UVAFyizi1Z7BA0IbYJkIAGnZR/gY1rHcRzZOhF54fWS2iXhXXj5dt2kKaDjrPen3Ta2
zY+zXqsooQ0srJQKOHpbT/BiqR9iG6VRd4z8q+DuWZI/qYXqmAVL84TWwnoBHKdDsLHH5yT/vU7i
RjKTmq3SROqFKSSu9E2hyOJjcUKafe7pDyyfIhwBY4Ys+cxn9H/p+fZRdRuQ7b1zOReGqs1yR9fQ
MZYkhiXoogIUOocGc+GxFYUFkhuG7EkVrfCqseTtuy5dMjaaD0jtkp/akulxy85/ZhJcakuL3Lva
RS8FRteJIvReaVBK7BP6iZsxQnkg5Nf1ujbtefH4pbpd+FohK61oZCjmlDQi0s+c0UP48Eh2r0f9
oH3HT5elpCgWKkYBZvx2BwmbCq998QaveAEAQLkul8wuBSF0h1CZY9ReQltIzL6YW9EjeNtT9gQ6
xmnEixBw8wBe9vRquKqjL6Ooy/+KFNkl5Lm8KEXJWf2fu7jZh3jwGSF0btU6Y/mzvYurew/lAK09
qu3mWm+ZC8XufVB2gZ+YgbIVYUKKGxREPbA6VTWaFnddtj5k6jl44DR0zl5fGqiqyfOyDfgQTlPy
8ITTpdgw2wvMSW8z8oVwy9viuFFt6FOcXQI928rhFGfXJUK9B8TjOf6m1mqDp70clsdoy42sK01o
gbz/RmJTFyzM49apj+vBCLxJpp8fY2UxDRm4/sJOhEMP3toFc3hqqKjyPvN3zYqutz3prBOkDlf4
8u1SpK//8Bu57z+IxdDSyvVmbuTWtNhejFK9onTXUqYINXbxKKRDH1gXhUjYOa5OisneNK0a0VGh
zkYLWsX8Y6hD6sU7pEDeOgLsy+6bRJr6ISsSWl/RhZyMrnVQb0aU0w6ABER4+nh6o1Tp0z2mn65e
X2z1xSEouPlmuNxvgaK/PYZtNpUoB2h5Ok8wR7j2gxah5t4tE4F6Y1GWEGBFh31WBJRslB0FOtGD
0RJ57fW5fdZ+TwE5Ag5mqJk542ORCmJ6DM9gnhZPWDSr+iGoZRlA9lCYIw6bI+oudu+xyKeNuJVg
/exDWKG0j9OkOwezci/4T/17CDdatqm4/2xbDmPdIkRnIge4vkvU2Cn+XJ6VV053xocP5LQYMJ53
CfNxTN0tbB1LAHBofgWW5cDZBM4byWNTbFSnqbeL26k5Ae1HsyYjL1WCYzGf80oCjBVHKkXH0e0g
jd3cABv++ZBaVZQfBVD6A3zAFqMy78JAWXDWAgxQEVsUjrfXFYx7/GNRTX549t/sxrmA6jM/pf9z
O84ZKRkXLUxGDjSNrOeYZPZxhAynO7KCp/Rhc4RnB/POxQVKGDThgAgxsAj/cmt1tKPYSQx0ZCvv
hCNZ4OwVs1eyKEiUhJgj9fminitZMB2w9l6pJKm/ucsPKKQXEGGa3DuJbkCayBf2yfV1pi/EaxI7
TWsPNzBI/DeqEXC6IIrOV1nwo2ovcx0Q91iVM5kZVrWMRPp/LUNusSHo1unjtLcagHgA2DXEOCVw
pbGqDmHrswz+Z0HlGh9nKqbQQUrNZl++6Aswe3E6XrUVprUoUW8uCRybE39tZHl190uqyWTvyvr1
+drBwUhR7oIXlZQQcn4iPzyatiEyr8Tr30u3jUICMvd9HY7t5qSZX8tvgOegRRCnXSG+zk2x1XvC
ipSuUEUmvVqy79Qt6ZSezMIFu6O6/kNJvlH4As6C7O3aMjWtH+obXXaW1vP1kdhzUurzfowCeVAA
nxJxrCYUegyzFYzKCZHhiSay5qHQAZLjgnuRXqSQPhPabiC+tsaNT5bgqG1tB1R8j2yPpBWeT5ku
vutjZ5hpA+uLHOm1L1ii6JiVQxrhoVF4iNsMzbV7Wqn5AU1kS0YQE6KE999gOuJrU5GGEK/q0AOh
gLn+/zadH+cS4ngIGNWNeu3IphASpcVmkPUQQyG0ePJ4bqVYwJqBTQywU6Fv7rrIEQpP/lV/YF55
lMMQdWLFTngPv2WDOeSQF3UGZ99jdsbQINWrLlq0M+YI4FMHaKIXLsBI9B7pZ4qsd1f1+fou2zSb
O7u5+EbGtzK3eQO+BGoa7QtZ2exaR3JqewVr6itEDBJIQhuFofTud1Uoc26OQhlsJoJr0NmL73QN
1EVINK0Pzd9H4dhdfK7IYw9T4Y1nPU7yf1a+9SifANTWcmaZj2VcOkHNkxuvdzAo3GHVs6w9lp43
AlPcjOsSgeRCr6wITL63h7OMHT0NQYBpnvA+fxSnrFRzHg0hGiJYyY1DKucsuQjIBQ+w+ibSQXhh
oAuFMLCQ04Qf+4SzHM9cvVJJ3dnM7u1SqsYcKqW1Cv3HcaybmG2euxUXxGxeCdz2kjbzzbuITCIq
ePfSK6tmDGqVwl1EJuOIpxsGYjfNjj6ZlpX+Jc4goOIvskRKMcPkdzyfJtPIZG27prj9+D3s7EK5
+9xjhbSh5uj124WHVtZLV/0IaQFCKtVEWLUf8Z6DbXyIqyT5aVzQgxtBc7aUdQwpabU9U/jTNita
kA66lFC6MSamXHcm3r6Sg8q/Zkwe1cVnD0kjDTxeVPVcxf/82r7z7ONvmIoEfJ7ZL1Ul+6mUkoUE
gqZdjmjPOZgI9XcB2NsuG8TWnjLu+5MwZIZ1XSs7dxIuS846LYww2B+zI3E/d3rYeyckOinBP6v7
IuyN+i8PqY/X/Zpq0QXxVMATmlcxbhvbWW0S0P53jIHa4u+YadSq5lGIln8uCVyniOuexpUNWUmQ
XbI1qLjTjEaFVJnBooRbRNQ87Cc2I8ta60ju5SZYro5/UamA7+IVm0+6EQCe7TEZuQ8TEBKILkz7
Gipj3XsTln7jh/G6TmB3VOZNX1MhI49+N17eX0o/y9MDBjO+e4cb4OVmuXUS1vcYfTTWm9WAUGgy
w93J2ncMG6e6+MBmKdEjhn3Am+RUku+tYTUAfP8GhzraqHf3I92OUIKGBSRtqBMC2UXWdTtLrL+Y
m4yzUyTU3E5VWnODhW4DqjRCrItkT1zJcWcyokLf6aWezKJNnKeUnBGlHNiqr7l0ZAlNJrwLKA4f
wPxLCgsOe8Y/RUYM6JleDVHuxx+E4s914Cxs/xLgs81Qqj1AO2nm0tPhl2VRyVAj7S4od6q2di95
0yjNzYqEWIQPDzcL1fOZh58mMb1W8wP/zChOO0WW7v9XrEgJBySV/slQzU377qNuzQ+bVRpBm4uG
9yD8Dj04dH8VepkGEWNVtw7KLQIC8je1RqaHnRDEAXyxNbjVzpM1yDYWslfbqMxps6tbG29DOq7z
URNMvfxBo5IHTdEkN5EdoiOURHsLLHVZrpWwPhGvaFmhkIMJAwfMfryVQL30uvyD0BtQKjebvdkZ
0jxnQiazenZfr8NJ7FH356RokyIr24WB7KmxxD7ozWoAWaX6oeXTYTNhrOPXopMAgV4DJL8moIa1
K2oieiQKXi5QhRPhEcf2bH512qnssWtmEzvPpAecctkKWusvo+x92I2QboDelCFZPOxfM+Nkx/eD
hL++NLvrH3sP07X/nXrhSXSKxfSU5p9Xh665X/Jw9Uz5RavXwmPZlsUzPQOdqtFZa0gagvMHjgW0
f+l/9qxIFKlTtqNpmKO5u5ET2c0OdxHIaBw1lhFfQDJuadZmAaUCuPi66IvyWZXSwNyeShrGuTYt
YY4U/VKWWIZFJAnTtUAeuU/kD8KXUGdvn09i94fILjajDJr/pm2rPN3ht7nsQr89JUgoKbCyZGMp
nbU5bEKidsGZrlBhJ6VgxmKy2/8byK5sPfBAfX12qDtPLiFcb+/QjlDSKAo4pyf0Orpj8G38wq9l
RUD3xt1+O6r1R9s+/yvfsX7L3q9WtUiAF9T5akHwjkCl41jPxS4RFfj0LHJQnpk6uHB3uNmpvbWb
KFWgwFrbd5YDqPbmYQk5fvqkANqoMmSkgZoDKVU8iSX/uIXugZUbW5SoV90Y7XFy17YYVpr1yO5n
nZfWxgAtfB+DSibFFAw3SLRy1QS5XBCmasaY2uZJxKJNkqvxzLwRX1pX6T7s3WCKCb9FoGylkcc9
odE3SDmO1pC9h6yYrT0NzVlL2C2UVUAeb+bnoEZjLcYRzsEbix0N9k1ACSM9CrTMQLF/gxe2C7QO
RwwMkEjlji5O2LbwM54mIcn/bVYSyk4aWUyluv1Ga/bxhHm3SPTtqFAyEfyzO/9rzGksr/46kBQG
+Ii4ebGpiQglbFdVbXfdcvOmoF/yrHU51p/VD4EPAYakvcKKXCLH74z69KlBdus38oZHjuolC06M
s2siiIMW9oR2PPwc7w9cPbfiZEU6TjF0SswfiSOyIi0AHta/FCzsMFX47MdKbLCorOIXLynI4gPh
2TzyiYLABkx3CpPa80jlmA9V3vJ/mblq5bH/jqMlE7eG8Am57b8FH0rV3lu3B4gH4w0ETqUJpI4n
1ZuWLrOmKtvj+H7eisII6j5IwDMlCwbSQzjIcM8m82oSelHA7t47pDsMho93Me5gFQQnhUFQ0T3v
MRu/rOmzANRBZ8oKEOFgUhl4vm0eN+JWFOCjNnDthwRtyVsrr+9HujzvqDl6t3+aSh0hFDAnbL3b
+GyJMLX62siAwFnBTYADRFY61E2QyMl/6ErEjm4OPnLkBA/bSCQctUjbOlBwVThCNg9203zFiEuf
HOKuWVAW0SaoSQ+oE24Yv6p7j4DRYQbDenAE2iUO5LFoybpe33ayg5hBJKDUJRVZhyOOSWZkDj8+
OVoJyDnkdrz28tdGBE/TKOGo47Hi5SGgWGUrmHorMqcNtK7bVYx3uWjD82qNT3TcFpVuj28qp2Dc
IdwgAkKDx3UgkbaCaumpbvTxV/TWXL0zQzEsorvcj6zq+LNsKJNGk/rwpgdb1QiLSUC2BSUHNzLj
vhKC3AYAeSOiT0Ot9LelvHvBMVjCr/TtrUvXVksyLrODtWlPHAhosYWt633IsjNNXY+XN8N0mok6
Sg6jILQFiuuxn33E8LsuNtYkXh2g04KFvb53hdnrgPPNMcu5ZCdCZnFDWZ1UNMMVEQy3v5M9cXum
9Ao8sQsWqpaOyI2Fq33FQUjanVKMLfkNzxZMVDb2WiSqnwBICadzP/JAKU5AnC6ITYLBZAGn8SpN
ruDPxBpLpsEGlfaHrZdEAKs9DPVvLoNmN5qrEEgnCvm2+5zItw12NGLDIt6JNZT0bQM73aIroNXB
qmJDtCeoJFCFPWTZZuJuJnD+H7wfhU9fi0SBJCph9nvNz6OJfUmAU7cn6xQ57RD3755FNyw86DIa
dT0h6eqHGjPjXkJ0leXDFcrHrz7NDS0/XQyagWEqJ5gCtIjjH9HDiVGliRZD2tVhHAfTEHMFYMyK
NfZEq5vGKtTL+RJM4eDvMFB7sKcA1cHNaeNXpkMe8gQCi5ulLdQcStutdkmcB/qljIqGoce6gG0F
lw2if1Vo6tCXGWfWqPXJRaoM8oPEwoOzZ0tgT8suHap1qpvmXVw9kbFnHQWYOgOS9RNHKXkqRmIL
1b1+6GpE6Rdbx9yxs1QQoCMLYMjQuRLamujqyugrnn+AReQkmINte53ywTgk3XjRx/KK4cfZcUoM
ilvZgrWF0vMV5KzdhaM85dZnE7ZLBjjx9mL7IMKkALWYdMPqcugQ+XUsEBLtjeNYJA9kkWs+DhXJ
cTKrrRiI7aEnIdENO13ERXYDDAaMdAFsDSvSvXMACKrRee8wigD3cMGfkws6GOeqRDtyUJsyRP2q
sGY6yphh6ACd0xU/yd6tqf7Jt7N4FYsFPDzwm+UiQ5KtTZuyN15hZCvBGV0Xa1rf1+1xuFrJ9Imj
6y2vog/HCc5xpnXK7ZPwJjKgmV1SY3PTz8knzAIgV+XUegPshIwl/gbxPARAiiVBTnWe+lFJgzW4
lTGpKpdk9Lq0Kkpc3B2s208t0GzriMx4abSSOn0tH+s3ff65eHe5785/Ct9Xqmm0Y6r/NwMTmUOB
r1JqpX6tkG2FC0pkrGWBAPUdpALp3ONUslIPyqfe7rTpmUTnA2becYhuSbef/SvQix9O7AGJ9bVZ
7ov5c0F6KPM/0mZShRmHCa7Ps7u3Xx8/PZT5lUaGnc/SYXV9+8qC+29A+wMtG47Epv3usJB2t2xd
Z9Ziex4K6iSgWtRt6r+ixfYvkJRArT0j1YH3p2tQBWWz2T2NFG9gMqNn0fyO5uubcdqhEEAREYpy
degZFTJFXoAiWe1f6Nofm5CLUPiI2weriEBEa4dFVf45UaCiBsPMxT/Rc9POeZrIC6z0dVqA0pwN
8R+3fVg7kfgQ7hh8XgqbmVlqpmJrKzLZp51ltSFf9uW5XT20c8DZp/bp0OVG5ZiirphDRxXhlV4O
saCe1rBUT+TFFvHHsloVYGlYTDwPr/MvEQWZ4hOiSJDNUPc4BDWHeUoInQmeW5oc6IuboIjMAd1C
20yDwFfiOaNTwV7+WTLnvPtXeqWyUr+v6kWD8kNpVupPNSZbpeKdLjhubzM6r503d983onVtQQ1q
iV5nALrfaMfWxvF5mIBLNatgGtgRDvnrTb2R9VaLOEwpZWzKuwqufcd8KFMOsCbakz6Ae/EGrIxT
k2zMbVfBzudNXp+RxFgwaXVzBWnhIViQXFTu7SW9qstRkKvDfGJs4Hqv762vJIRkw0jwBvpSgc5M
2L5iWhKvFb8n8knvZIeemKsDBkJKRai06jZ91J09lFnoYkgiPVBehxeMpjHV+scVEPxpQlTtYQ+m
OJmm17oyk7ONEsVjsWgRHI+pMsHmb1q7DsajzbdV9UZZnkmV9L0y+xgZcmSxiWWLI3r7QiRcL8+a
NZgk+TfiT3qOLtctKgwvsR+CvThJNLNlRA9+VXIEh/nsdKVJvGQDC/Sv7AYMR8A5ZyRFr7vkVns6
qThRVbdRocDUgByQ5vsWM9vI4Rz2fzj5dVI/O6pLvk5B72tIbLjbZRicXNgbLwQ/vSG0K85WZPVu
Kk8GKnadO4vAE7NFXg5/cjroODktQktS2u6GzFufU23KyQ1mf1kbHqQ1tlbGJdTNBabI8DHE1vtM
cnwreW+UuEkN5/rpNuMsPoYLEWuxLzyAH9hkoNJ35bF9Z2INta6N/Za5M/nWYuVmkWrgOhZwTdwr
5DlHQFIth1XuJLHLzWyWTl8liGTtX0YgD1Dzg2E7rv8cgsKFm2BGgwaReY8h0KTIuk4I4jzJcI/p
25UvFDufAwDgMPw2jsrhTEU4l3dFq97TPoF+GEFoPbeLx6s5/tcC+T9+QlOjNVT7b5HPLII93NO0
mYpwfrXeD4/pCL9UlliSFelL0z5Z16yQkGZ6YMHowcFczqAmCn0NL95v2Xpi7gTeoQ+/K78Z3NhL
XD8dHheMu7MUvqdjb8oNplT0yeplAAFtXIF/ebeMfdXf4LzbamdEgk7KhgL6YBUJfPbKG2btHQew
zuw1g3eF5g8g2j0lTOL++XrWmPmu589sbgGrwYrShve2f9cPMQVdu4LwvhyMEqVK1z0TCtCvd1+K
Gonn8vKiNeWLTbW5bXxK56UsWj3X422mDKV8zSqgDHcQHZFfi1llTcccwXdNeDx3ibhw+ZGXyulc
hJLcKvZrTRYofbziQqEElXa96xtC5wDxEtWFkspfnKBlbwj59ECFuzKt1H7PeUKh/5W2tTQa4wgZ
wCV/KUM3yZmMSRAQAjvuD1nWBthGQBQXa/T1az6TYz9DubxlW+mOFSx5iuRA47W6FzFSGAWJUUT3
1wg+gpdVQmva+qs/7i3OcSjjOgB0LLc/wrr3pZ6vv6xzQwiBU12R0Y7PMaUPByWwjdqkQsEPd/Ga
nvBf0kP1EXJfjsQO3wPmRlhRsk47q6zJm6E3bKR5VwVtddD4hT9CW6S0b88IfnfeIlkbUHdjAezo
UY3g4IYzoObQLRuIBTBcoMLSF1QXmW+EaWwqrJWIDIDqBShdTcM9QeFpogL7xXNtIX6nqliFwiOU
np85kk5YsRhskKS2Br/8lmI7AVGu2edmDV2l9xXQQliwcL3BbIf1wsfn0tV8addZKc3qdaP8XJUQ
HVvRZauFLS4gYCh9tGbILow/8TZHU6czF21G9alnjqDF6NSvH1iFyGquOnL0kTb9RXckbnNuTDTp
n7EuQNDnIaXxLW90OJE4nmXq/e8aabfjMm4tYypNArHlLbA6KaRCeYLvQyqOfUIpAe0SKj3k8rNZ
XnQv48pH3ef8nxSrPz2NA8uZia35Zv2sr25YRVmx8D1YtvDvojw/VIZKJp3OHaa/8vXJ5k/bFMAE
FmpqpA92zHWuNI5ytiKe2OyDcqWWCFHSARpXBlfI41KnGWndM4cueCLnyjA5AXqupTQ8tRyG3+Xz
l2xb3Q7uwqCrjacrjxB+EOONf8iDqWF+IXyEkf8TBrWpF7TXhPk5fTRqXFt5tCeCdacYJJFDfvRG
PG/pGtWCnIA1eL4p+LSlAH5vnc3ByFX6sweQ0XQavwPqMSuBEwes5MMCP5fliAcS66hESU72BAV4
BVvouS2lLbHq2wQwPS3NAYE+OzXX6mAXyKOC5FlKf8qgmfq/juLVtYhIYikhinP88qN3yVrPyxGQ
t+aG1NF7RyYXESzCQRPQCQ3U5yI7DiB8sd04gRTpeZDqtLVHT8vGq0FtUOrhBUY/l1kjpie2Qd1I
loiClrdAaV/Ngo4cdZs+B5bd68/uKsUHCk77mdy5puOs9c7xvJv0GL/R50GrlRVJt9XO2QUPToCY
8WoPDYVDzpyQakSvJJ+Mchex3U94poZfEToj0Pe/hMtpEneLCtvWM6XLMr7LHokRYrC3uYTBrVW9
pmm6rursP7Dv9595Zkvznr0yO/IuxQq/LiSyITmEPY4VZ1nK30dj/2TOwoWNt7ZH/07Hf0r30Wxh
9V96ReEs/hf26aEJYYPzBZnWMMqmyvlgdQJVxz1Rj0RI8mEUbaGjAk66o9okg3DHMjRKnZ9ua3OT
LIvdtpBVOGrLPw0D1xriv3YHHyVQOIxeSmEC+z0jeWA1V1xf6DrwDbwdxbiZXcs3vFeVQPv8S4Xb
BQ1vrDMPf41ppqJnh9pGp0jfjG6enxSdGG6vIlDk4bsMiaOLScxVy8q1rdRwrNoS6+MS2YKMmP+c
G+jVRWwySSn4x1wOAioH0VltVTx3YKOF/c+q2qqm5GSY2rf2BW65M8TEp8XEwbI0Bqr043QzGjs0
qtmSdNmHiTlP21M2sElP8tqElVInNyCsN427QR43IVH7anVW5wWIA3cZEBoB/I1+dXz1rU1ecTf1
T0l/hzIFYdizevNNW0e9S5mCC9tMN/DHocJvEwBuqUQeqIhTqWPP5sdHSNAHpBeAxEpvVBK58BZE
47CUlqCRtDa+7wKYw8GxwFdyUtvknSOtI7aTj407Xf68MGFqyDQ6mLMq3hlUnfytPUqZ7zmNHaPI
fcyygsRlJ2LSyTl/gAUHci+PbAt0LchHExNqBuTyzEz8gqs22cZz1WXqG0Kd85p1sx9Du8TZIAxk
bUYr7WfEes98GhJoPhxvndWi0i80fcA4bk4Bf004LhAL/K8SIftGBOg/ZRk9wU36CDzLmYZlQEx2
7RBTrKUlDw/nfjU4EruL+9+BKD14ZbvgJT/T28AzJCKHzm1vqyvknymVFJEp+iAyx5O29awh6nWc
ZhLlekUfRSzzhY48upk93I7hYUIogMsOdzlzHl4VwiguT8WhanbUqNL3OMh4Yj0CnsiT4J7BTpbH
Vktkh2qwKUxCHyh1+GKJmW8nGHlQp6R0SCro31DR5uwM4yFcIBFTjHYlwZgAQlkmN4k0w+W9ZBJk
udFzLwLexzsFoHe68U8/wo+kuR6+yWViUlhABBdesO7MS8gs7XsX8Ii9PIL/eC8ezm4EkXhuK0W2
xIHzwOWq6HoOtdF5z7DjpFO6DI1Ur7M2U/Lyicuyz9q+/E7FCz4hFQfA9GVwe588Lp0kJWSmoEzY
6/cXU2HksUw0wEDYLGCImEZfYRRaQFVW1InJUt58P+WcfAiX45e6/T8RkA63V9T+rXGBLDu7itPW
2Dfypx0bF/a942Zt7EfHnsbJTNoyhaoWlqX+Ai/MS58nvfTUEIti8Ltne6AYqppkqot1XOdMd8uL
DcecPQahs4xESqmLMQytdTxU8+wSEiwPZBHFU5WjYE8rQChHgyR/U5d6qwxopIA3SAoXgu9kx0bX
lP80/+u7rGUF3cEpothJT5R6GnKgI4+1TOvbleJishXg
`protect end_protected
