`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
czlLbtW1hECJxXUk+MbFhO0XmjyFReXWlaNesdaA5W7AQJjWu3VVNuQw+r2Yei21+9kWRANs0u1t
bN8TNj7Vmg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fKBxfr+pstTIKLVc6oqTFGlWBji+1dw+fTUJQwAQ4bWm5UhTQ5ZyXGdVQTmpf+8pdpKu94WLVtXg
7wHsPx14555KfmRSUBa5IWgcmVCNAszrolmizjcpbqWEy2Il/2AtaMpULwWIdFABf3+AjA5ZobNG
2UBdUb7k77cDJl1moO8=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mWMPW2uj1seG339t81enaLUYEJmXNqjJQ7vgYDCwd/S1rGKlPn0amsUxT/3JCqhVIyD2uQR8+6V6
n4nPJ+fiEGupVp4sT5h6+A1+kDI7ltiXABf/WTZEu5N1DawyFDvSLQ1/sGJtXwTkEl4k+bXWMyvi
SAnTH8k0+zbkcALT2L8=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h58tDs6G1Q2JLvR6Ac1lCW/zAjvlvJiRNPLpqZ/Z5afVhHWNud3Vl8SnyIuFgFuc88R33wUa2NEW
LdbTFeLVpa40uw4fbSeTffuD3kJVKjvlCsyJ9NO32QrBX69J3hg6v2EIZvhOyqFsPRKpyzeK8jWa
P/5UBEEgsHyJYCvwi8tFGhOddDUfBiRmRPttEpYFLL6Tic4wJLeEOxXQHospRH8BJWQR/bLW0qzV
rmef3eo1rCmMSZ7h+KtU92T/OkElYmuY3GP+OAmEHBvvxlxGcGIM3Hrz1H3yDTo7v6XNhFk4o7W+
w6HrD1L5mNIKX3d0XQ1vzrapkmaWyzxUjXuylw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FE76BlH7KqvO5fNON9ddJDc0D2G+kNV03jL6C8TUm8hYgAASN26g6OqLtMjQflkgugb1kyeAfrqK
SCdmFnwQUmGP94bHHnQz90J5H7JqMpc7qFo/z6P9uHzYjvPE7sh1Vxuj9VvOeMSDvEZcC1tTQBCO
YCbfOHLQhomKn63IgwguxMaYJG9wZ/Ln16fgjjVa2kIKoNE1TH2+GG2gz5ejn34qcHFF5bDgMUgR
1gBP4Xb8sReX5gV25ZFbpaDLhO/XMV3qIiEex87YMQEU51gdhbEmogLkUXTrlVFgbVtFApoqKwDd
EClhGg4k4kSGMwKU+yyVfzr88VSPG7PaDBduIQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GukkEP/mm98jNTg6/bE3+HAZO374v8zE+196eVMdmR7FZoqv7xAVYRl4N4DRi56agbpSAmbguq9E
Vmj30HyI5oesX/fJR3apiPbueh1hW1DYS55xFBYRD5HtJsQsafH+8VBKBTgxn8NTQQKZmfWGRfxh
GrZ6glszDQOAUYGEobLtCFt+cAmwswi4mPnwYF6Jkd+n2RMS1jmCDJzA5c3eEu3+fZ51tciPMTTx
PqFCX43YC6hnVOQ5FQGieljLdAZNI0ZyciKp1XzRF38dJlFNxQDpuf0ib6kfWKfMnfBH6a3qMJ7C
jzWoOzki1gPA7orOG4xrGp+CfY3TEQfBos5yag==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
rMaLfNizD07KYvaclaU/ywa7nl0IkgMSMxE5ciZGJDpQYlcdrJ5sd29IvEUe4pbb1v5kWBbuShxN
jgjKBARKXj0YgHl0oduf5Q6uxU3oodYk1vZzMJvjlPdBgUF/WKhVVcETrk0dcrWke2nkojK0/T7x
unzPnEDvqckZSw8LBGiGluVmWTry5DptbqAspCEB93tgZB7ABAOOqXYBgGcMSHLLUnpIOFHMNhPR
sCwdTONA36jAHsg3B76Z5GHIYDZuD6LomoGrq2YXdLbbYttIO0ENtnSZ5cN0AmM77EV+JalFzKiN
Ruc0Ydiut5QzfKyA45AZ2FAwC+R1fvrAA9urnrpaoqAfucyfCp7GND4Lt0N9ZetLlsiRPk6wcz2p
Hp600FjASLgJD9rvuvRCe2Ir1wemeA5/VHx6kRQF9FUnvIt+3TQlcYgLRgz2DTnW5LjAOQphvSLF
IzQVpD2zsgY/QLPhKpRlz6fq9MG+mGOdEkbuHaUcnO4sbSFj0yfcdC5c5UloGY85q1y1rFZKzsMD
Hnne5bnBPW073OGzUuxQwuB9SnSDUQAteYCvp5HUqPyUi5mMUdSoAM7H3/Of9I7dJcDsU5FZ23U+
bHjTvKg1d1vYCo1Jk7HCjvgD9aF54F2AorTkkn1I8M2KZR9rVSvyjrXfpuaOwdk012NGEry43ZAq
sqGtpopfYbypJpXehnSCCTek3yZi/+kdL7szDpvIG5xkktlqvRfDPlk/ViRlgseDaLQSrnAzEK+N
8K06eFTeoXQUq9mTE8YFq4gWhKtI1XlTWhFSIj70XZYxO9Z0et2kV4hNQfFD6FjGopUamARI1eTS
vLMDgy7Zuo65hYLPAIRKwIopBX6TdupGcTkm7aPouKJ8BGOfVaCR3MPAivde2meYT6/AO8cQwORY
X4yppIkdBBkr61JUo4XJ6andYVt8na6Nj3hTy+nM77PLCkEy/fShTyzdU2QhZeuNCyYu3HzlEYIU
kmsV5eThU9qz02Jz0qjmgrGy4Wj0djWFwnwdM4rtRFMIA9eEiWOOcKN2wEIHqQ5z0ggM0wpRcX2t
Ik7Pu4aWBs35476whJq58I9Rtyqiro6bEGVXcDge8jyahEHZQegZYp15V51qwEZUW6syOmqAoD5n
78soBWUDRdghrpNCfRIglBVNpqkDO3AVm+zE3nKmXqZADyU4ZcG93OxSiSBjILCooHJaH6+tYPNG
shA3SbmDohOJ4CPBKr5Tl1O49yhYG9YDJlsYmm4dKphtXIKkZgMUAmKUjZfAkJ/Zo0EDsMF6qdWy
Rg774NXwgLEAkRV23q6EbC8QxFn+P2XlB3gVNwG2xhPXTXVbRcel/H+7iKTDxqtT1QTOFazYhSAX
6Gfvk5Y0+lSmW85gj1uUc1WNqu0IEfHKOiCNv7t7tmjf56hmUTOTzS/9CgNmMgYAAeRnQ9zrcMAg
QhqSmQZ+1Xx06v4r6OX7BizGSXnEtGOm2TUnR6orj0OU3TPtR4Ll9g6HkYH87XADaZuhs8dTk7ob
EPr8NChlcLslHAVZsKtGDQuGT1Khq9WUUzcDiAGPMhD0rxczmQbfnB+vWYWGpBlHF/SBuWs+kbS6
d8+xziZ31XLjhkdpZ7fMAYrywrWdVItnujyZskk/C26pTRR0yE0kAXVG7kg6qE++yL5OJaE5jagF
8zpO9vKM5ym8p86DpQLfN9iTeR0u0WaYftZwWOgB6XyNkaL8cppgosC5NSAC5qxVNpvujx8hgm8I
l9ZJuWU+tA1VBymGpke5ztUOu4V41YAaVXnQqtyfob8jYsj2XVVJyWRNk6a7bEzAe0o2D83Z06D3
J7NAiUsZirm3FgvrZrqRWvtfQtLolL1+MaT4raswr+jfp+1ahbXeniFFFxcKB83OzGwcO6RsgnT4
mt0UVX5WZt2FmEE9ABOntaBFciLBIF7B8DComkWvPhOjNlbsOkm0REfJFd5+P2aKig+4VlNP0MFO
iptr3ctB8Ig7aCPg0lDJMZNeYiN1RbJ/WxIPhrDp5bWzWkOHTNNpp6kX7gekU8i5V/MbnX6EvuiF
ow+W+gDQYh3r1iaTMRJ0Uxg8+umWp0Hm7uQjAbdxR3OLWl/XhHWeyroGNQmoc/llc6ylSV36bXLW
7ivlFqRCO4zBqmxtsh44PzLhHiq7z0rViDzpBFa4Ozy1PYAx3thfFFBP/PFktuEP8ROENOV8LgfZ
ol4J5gyvCna0XgptbS4XRhygKnIxBN2BZkfr6SsDwLhN8F6kGehgZKPoa+F5uEizcWQECeiAdii9
Q/KK0qC9KfEzcm8l2FpBBTWRE2eVOgq5m7qClYItud+dIaqHLZ7QhEfZvAOUjkD3uPvh9UrdFf48
KCP739ck8HCl0BD/9JnXP3dKRWykn4qUDamEAYKrTd0N/qZY7ue4PofVNlGJgXZVA6CJNRH6kt7h
BKTIc8RwIDC0f0U+WXnCauWOPEZz5V8uvHvIrvEicjDnyvFGpHQQ+GURYb1K3GI1X6Sew5xvBADN
hbEjuvfbtp4tDoSomBSOB36jg/0IuHtHh947FprNQ39DoNYe7wCrjpk/c3OzKiHGT8itIzqJ2rcj
JvgtgrxuU5Kmq3uoncm8jJjxFgiO+CPL7JjQHhdd9+O6zTcxNwLiIs8oflT2djr6fS0np7Jj3B3l
La5H5KFFZRS6uHMFO35SMOHzyk77VHYa86EjNMsmKQJEqzExI2+g68WOIAG8uRftwDvwiuwT81pw
yKgHYPZ6qDYHtWlEDdZqwSUZsOH45z4Q+E5GWj7RU0wey/yho+fOrSV1N+yydYT56KCxWIBCHN8R
IwUtlKh0hl0P1BV37rKD76PkR4y2DSdSzSkGG/j4wG6neKdZq2q7mjhYAA1KfO1oXD1J5RtUqBef
CRx2stsjLhpRp2kAZg2vGMLsdgsLjXnmIIvdDFJOgLmUlk1GcMolb/nvVI89Ao3psylTIF4daNMA
cmdpku8Da5Cn+G3K7mKSkoNKeyySi6NWKVPcW2b5JBkv6BDonay44A4dKekvzEsBzhV92N8E76dy
aW5e7wb3NdUH23gM3G2dUFYY+EGdPZl4cf40WrT21zFVCHKKVtUB2cJUPKmfaNGnxoVwLoVMaZw+
RHXXlNCaQ/QL/nR50JPUDO4HMA3f3hcG57w0R8P5ut1K46yMrAQk7XdMhWcMoZjfib/UccG6Kd0C
I3t/zUO/HzAEkMZdoeVjy14myQPJ3aDVrDmQaWPjihCZz2xvSI1x1ujvmIFFEjivADuHSPXxZcRB
sXxLWKSWus7Pri64vkfuoLze2t6fy1UWEolHGKt4QU5kT1ZIYSUldVJiRbrLXM3axBlu9uMPf1rk
aM6K4di5khUtJXk8+rYFdSFeAG9vZtlkpTTdhyCOezUu9jOPYuUFW2BkuRUG4V8G0pKEujQ9PsU9
Udwn5OOJvDWvJ861FkZeoorcSOuI4nttDSDzg2mKDyrCna0Cf7IMCEwAUz3rO6WDMBG0v91MCmwS
pRCPf1FbHB+Fs7Bdf9mL+PycmwJwrOn1R0JBFSK0zMttFg4n+q7IWd06TScsW2YTEKKYRLdU4UI/
ofbKSeChk8KVnyx3cujlWkJHInls8fyTGWShSfX3uzhLoyeAOf4Jfai8U1isO3QddR8xfGvklAra
Fl07XV2onrotUHcAC1Yk2BMNIe8n0eyMN/DJDb2dvK6Ly2h6n7tmgjWM+6+Kn6/a2abyNVILl5IB
2d0xDGYa89xAZ+hl4iFDOEsCqYiAxGrgW7D683I4A3zg5xMQao1SpkXUTCBmKCQJD/OwV2Dalllt
AVYhQfEH8VcLmYyWMB2R73xPidEZSCGA9BvxNaxIsu8j0tj9JaFKM/d7E3fbU5i7EHgmkoGNO0B3
VprJ9NloHCkkl2OHdnHTp8E+1jod7eBjHyJpG4H5gwOiZdIw65+Ojs6yktQUZE0khAPuoEICqfL4
OyvmdqkG9eec0OncBp8VJxC9L2YkJCWAtz0ucMGcWE8a+sU1ZgjgaqOF2S70JkicErj9cfsUD99u
gRVtV0ABdKHkb+2eEXfgRQqFTE2/tGNY1oT8Sf1iS/K3nsyfMAvHFGcFchWCZ/Oob/Zeko0kOWnJ
UtXYGjTq0Ac4/jDqkbE5jlgBBEQbHrL5ZA4VpyMC6QXprPNEB5XTUo6dUSOPGr3ZOFq01PJO1FPa
+mN8tlslVK5jWQOe7alG7ZM0VDXFkYGFZpxAy3ZLwUFxnt5pQEQcxRZqZ7cq/K5BpAPtK5ipbjTR
FiAIOGZrYqZpa2vyDHlAueaOF2SLqXViHLDQ3YcffZGfLXVqiQ4UZsJ3muQNmRBRZeGgkvUkWQS9
B9jJyjJWnEMe3XRXvs7ifpjyIu6IdzfQyl8/PD8IQogBey0XYcj1kIMOdd/uhxYTYEO5edZSmd+R
ACH8S0AVStCAoebf0vv52QhPzN99Q8/rUGLR35RMK1DRvz+t6/wpWeSC6It/YrZx4rnDB8uSA/6T
b0v+S9ibEwsvnVqgvb8KPxuqhlbmtVWw0BCrDyVAKOi0HQaDpB982U7AKFW6Mt2BowFbwSuUERPH
1KIklu/6e6S3K93nJ5L3hq5awxoxtd86NFOxkpvoL1i6x+OmRX6GL/f/LCru3BcAOzyGZkB6mRr2
RyoWmUUZBkXHW5cF5eW1RjlDZOVKIUKgunBresFJ2YZwPLo7A9IpcFxAoYdUvrJnr1RZYRp73fPd
o4u6fPV5n7KFfphX0zJGLoSh7haAqHkpEY0TAsNLFfNEiMK+rBzWSlFmQQvQsC+eZMU0gk5ntymQ
Oqwf7ZZCxggofQ/1XhWYLJBMi0mXnl8RGMrS14T+umblF4btiUVqWlQ8fJavhz45/5gQNnXpBMP/
bIcNWg/egaHWMmYPlT7dWojtrNeto7VbafE/NGPulq4u+FjEb3JGWDu/svvUqWv1Wy39XaO3d74Z
b+7n/uMC7y2pSbKVEM6d9vJR7Wdrav7iGAbPRg4b9OJz140L5HantwrYAgEksDLP/NP42UOjlIab
8LiJvg5ultCRoU+wv8sj5Q/hpHoG5l1b0NUpM6OYMBCyWOzLGNH5iL6o+GQfDheH+f5X+M09HjVI
TAlg09bBT/3k0MdNF63OkG+hj+UPjaiSs42zcefH+leypID02X/pz5jbJjWZuTATtw0e0WRHJKT/
576HSUQbhTRs1f98z77JdjezEkW/+AZxaIlc7n5K2G8JC/HN0UAZOWD8TVyeUBvawF1/MWGYoaWB
ViMlY5gxuK0/gZL2R5NJlbEh0dQ+AS9JiXthEpeKt6vc+33WKFTZAgbZ4oIveux6nIKXYe9SqrSZ
3FKR0WW3QQjsHFlHRf/TeCcUpSyuQaIZvCSi8FQW/H1cCWFap0g58TqiwDldYOzGc6NQwyKvAqii
5KlJGejnlcwmIYUAbmJ20wdNq8QwZe9LfI2WPYCRuZuzXm2HMZbTWThC0vOwdOXfDrYZeGi/fBAT
KerB7BNBS2XtnVyY9vS9O3XTT+SoZtSJ6VVvV9610Fvg9+M5DMTs4KMt7KwnV21x57cK6PHTvrLZ
bFRns9O94s5mOs5gLNyroo/WjTO/ZvpzKH6iu2K6T4V4rctITyraMsgB2gSb9U9G1LCRxDhXH2aO
GF3WK/ut+m+oR4WO4X9a6h2r87Zxz0zaBfLIrm7wWHxk7cKxt4+H8oRrsIXrAE9YL+KiSr3DLXo5
KJxxIbKrCtQ1zprCi1JLe1jNMt7oh46OZJXFmd8feK9BAZdMwuZhkFFledkHTRrHlyjIy/6Tz30G
3mth+l4EFleG8rhawLkx1ZewLvctYZbp6qVpmxD9eviLdvjWOdkCNMjmfiMzjmaR0CusZxLzeDmF
J+nMsMa2pLcOOYoEYHU5z72wX9oODBf7/n1wbJGK6BY3e4jL44EXKNA3cLcqv0lCMwO0r1QO8oMD
x4Lxumsxl5isfCEZ2LFB78+/kBsM3/YxIjulEDSB3hmWwCeDT3W7Q5uOHiGUCb36h9p7ZSXKKPcX
Fffy89MaTAFM1y0kMbHl5UrZmgaoohuOy1mocc0Qg3x19W7GfCvlEa/1nut1qof4mroTX/jKfwia
MAoLGWT9Tfq9W4MD5fYT0m0w65RSqxUAC6Ib76MzUhldGtGfGWJpKbX4gEMM9up4oWFX/v56Vzms
zZw+OAfX3HGxT+t9L62NWFt7cDONVDxk3KLf1/kbCkyC7/AMfBy7N9pJV3MPH/7bqq9a6zxzduX8
niTFvyEHtf2mqhfRXdEAVs+PPx5JTPMpE8bvFRxQLd0Kj84iYNKiS0TULirmcjohtstdjFRJxruD
drE9t84hnMNhamn+4rgbs2zWiAX+d48KbREWlYFlolqXGU2okU/TyRCQmeI6fr8mVzUCM61HHxup
AZfr+O/anwPSeX0q04GMh3blZs8vGJhmzqWdiTEzx5KJvQ4Ol03MQiyw7DEoM/t6JSjHSspw2179
v9jq1/OcUe7YXHMcssvGaK/Uefm7pt3kIrESrkAmqNsGOkaVIJH4a4KOjsV9XHqzo261+XoYPCxa
NXw6kWBpbOwtHfc4uwdgSMaM/mjTqVLoxVE3dj1gtjoeIkMAS0IXe3gfsjAH3KjTDbv6ENPJvl46
AV52U4ZiP+zXgz9XUmCTpJhy/DjHZFzjp4EWeeCpMTgJOtDHiFKU+d7yq07HrR35W0DCb+o0RQP/
H+itKUPctm7q1OG6LGeoiJid09L+HmOIyI33fHb/7Vvk1LTiCivFBCpNnDPzMhIDODNwfz9/GZaz
dvV88qnqhfL/G9fMxNVwUFLeNqhaK/GmXT5yAZu4mvrpg6pWK5fNAon5UmkJR65L0n5EfohV5Eg+
RPa0qFje9STWk9Bp/Obxn8B1TiW+MqV2HTgTuB6F2Zhbkev14trnWGu6a0/8BFZo4PaloBF3TbWU
zJ4QeF3zWGIdaBCLuVjdJtS2x9jgCIRbThEdyGRRId3vZIzmqXU0tCUMsrgCnI14Mrj5LtFP9G1Z
6U/mM53vWopoZJJ/gxUaaHm4gXTOqfq/skEbfV+Szlca6z8t3GHeHeLZtDpz8WB02w1CSecfNPh8
bR2Kk7c09687xaK5q04xESUGHENcTsxNpKOyEu6EGX0Urp+VYx4of06EJ/I2rzRF131wagFC6iwL
+oY7uicy3lxwoysxoGMDFBnbrxg6ehL7SYwFY6uvbH2ufIW5IBpGswp6ZeW05X+6gHo6XlgF+H6+
33B/Xo2MIoBFICm9jhSjMvS2BuVNIBvuXFOiQycG5/gRvPXASr6XWf5eQVMa/CeL0OQbawJ69ASw
HH2m6gzxHYz0IQZbm+YCOuOvDAhHENskFIGG+P2Xh+BNIX1GXbPp6FEoldED3x0bL+JXC6wY5yCs
DKPv/QVTDYzEzrLGOpqfQshppryl3Pu6zZBsgOZ1PGAB/QtTSL38DTed61Cy1gMaIz5vggTXZnRk
teaKiNytRzZjM7lmKuy1l5Qq7zehs9+gr4tEnOfggYhJEkgicLbik0Mmo32fwC6L9aedM4jthTUj
aeujN+ooVh4YJ6d2Tof3AF9adaYKbVUMz5rEDPDVG6Isj6rRWTtlesR68XhxyiUAkdk3i7YScpZB
PREPC3T8+G2o3FXtqbj4fXlFInYFgjcH909lCvUWwbytSDBusGrwF3Qd6hvQOzJ84UQWJK42nKV2
7n1caM6O7aIQWbYAYCN5EHwSbNZFPt309TFmmmGazZJ9uAHQsc+TAMK80sfmEudTnowaNFuiQmRl
IB2QPzcGm/ORCV7EwIvtXL09aT08SUbRz5VxgWBm0UbujErhOJssvnucwmlvItG7PKtlMb6ODy3t
kZ4P12ClGVdaGINE6zu6UqtRK0uNWFEg4TCNJBN48dVBo31vAiX3Ft3XMItUEvKNUygW/XsAFgMz
Yl+DcgCdZf+3to5jZDb8yGdlgreKa+7mDE8Ej0iZmng157t4gS52HqiXQ4ZWh0PEAZdwNhDB4Zfa
KnqiW3AiShHcx87O5zkfmmKGAJfP8XbpvCw/Z4ohXGG+Y8zklVM+90lKgFC9h1gN1g5ABsWtvvQi
YjOWk2jJ2Nu/kuS3TZADlbRlixUl40+vr8XHwwdh5OCdeBhUlJGTQCcpAWGxHfu1LHD9EsMiAD7/
NqrHVKgqzFclYua1f2psOkeCvzFBS56gR9nvnPuEqq24T1QK2sxPeLjnnLHuuZDvajLyvk0AR9hG
HwRAavZdo4FXOWaVJBbVsHO7Jewvyyu2TJ93Ro/RrsjbM0jFLrW3Qb9HmI9ksqs9f2vS2o3sMX3y
CKig1TfxSKAhf16ZUdoz0RQk9spj457JilIMT5zPAqOJvhm4V3URsdhEhtoH2RO1GYpSMzlvHjXO
UsUhUItnUAn2PRIefJfm/lvRFR/XG65xUgCmNZ/HuK2MH0bz2tc5rFwmeIQPKNI/NYKr086B+4pd
f4nKc58lcSekRujztUcNGB3El7iPrw3T/yFpe+JBGt+sL4LEtkCSVErF9oCDCRDLd/jf8NKLNoue
rlqIBqf+akMjO9YOAkNLMrbAN9fWPVcb5I1igJTOOKMr2rQowaNkLWsrEW4LC2voH0/i1h21XMiW
sD7lHgnJmwacDlnFXGNjw+qBBl80Iaatj7qm9S4XxoxgeMbcZynNdp/hnOUC6YqGRvCrdZXqXXmq
f/q+CxWIHqpqnnEsn8LUmYHwcc/uQZSpUVhUDFDfBUaUMo0kjHbEujsTTiuVj1hIItq3nOANUI9D
FIe5+2OQNRE6FlqpOYG/F2u0OKv5ieGSlsL3Yc7npsfvHrXHgRAYU+2Uq5QY8zkSLO4xb6nz/lK/
CoLJgAH2W0rgAeFyOOfQGnx8HLvssYPBQVqm7h4MYfGcnZ9bLcDlLkwEpERBgYQvLuKZWpfyZf6d
xksyHSyHx9FaJ2XoToslz+tFzpysbbFZc6VNJnA2UWFeyJBChOZMDpEEMTs9SEtkGv8iyO2d2cm+
9xDwgjdXQtZnPE5BJEtfz+ZqqFzCqsMgf7vXlRce1zSB73PcNO+Uh0S7Eh00Z/a/vPAqBByMP6mf
tJg0CfNO2c7OfQGQhq2/IHtR0Y+O+rmxjeYhZXBzQY4zIJq579C7N+x4UbM0V50fBxagxxr+tDjw
lNQn7sXxqcRv1eqAftRWI4k9YYnVNZZsP5bpTnmR9XXqAqlWrNmpERfjNh9gMP3GkDT+pTN9dNmL
kfu5K9Qfy3TKcs4WRRVYcu7o+XQyUJgH7rYK/qibmxQvyuy/e5V7s/A660PnEkAoJRcKSJ7Zb+CY
nQCTfQcpW96wuN0Uc0ndHWEOo3BPzbZGjoVWGTxv2CXIzS5TW1Uc5l0Aw0HwoXef+nm9qyEqETym
xyh/E/HjRWQSEL2xOHDnnZpC0M8YOKhVXdmc+BBCWzHnY+CDdc1FJxfXkuKVD12y5BJEZNnC/UBn
CO/ywZUucPdcJ3kwxbso7P02+3K9c5DSeLj795CaBVIvk8sOgxLonA5/+2Fb9rJe3FfgYiDi6i/Q
1wFN5YInSMTGPXT2xZAYbiqDKQsPGZcD/3DNecVyJONCHb2CXUuAAvGwwr3F+kyiRT1sEEUgJT4V
et+gCYWNquOYjsK8Y1abOndWZcWyf0NLmmMRGBRu2tg8BpWeloulN2bMM44dXjf0Rs8Mi4XDAZ6q
ZgQ0DCC4KV7j1Y/fDh3p2F/gwZPsOQqNsBVxrR3I0E4/KwV3sEC5R5nln+PbAeXdcc94QpD70EA6
+lkb/A0PtDqpNSMgnAgITq7UV4tx8S56wvDZ26ASl8Tlsz6uTSCgXURS4aXW1vfODVZDdy/t39IH
zMHSqt556Z7YP1FYTVlQtmKWt6slQbR5Lo/NFE3AHbQrHyceWc3NVz5GJgeZtt/5T/J3pq1bIhIF
nAMntxITPUU3ZE5uVgx3ZIsV/Xf7b/6tcOdH6BZ+EmtK8HiVvTa6Ao0d1Fjz8pWCW77ufCrh2i6p
GfIhFRQf5ScsbRNSYHOfLYIcAIro/bQ2dKcw1sHnm3/cLVP9pwwCPtDaka9Jene8T/sQcjSxCx8e
icjx5vG5sATFBY4DuLDVu6K639hUgrt2BRSJKcyg9qT2f4gQKrEaLQ3uchcbYZU0p+vvFXYbCj/9
i07CUbPd1/SwRWllXtjqSyQ8dP9r64TcOVuSM4C4hyVPp1+oeNFMGbTylf8SGzPXtCrFttuLgvNy
cAP/fCS1P8fJzMPUcFR8dvOvieh01eh54XLS0j0quSC5gJQ2gb9H/ISavTKr2IKjgfCtynlrHYp4
nhfzEprVUyVHiJbIRGHi0F1fCJQA12vrb3Lxx0hvffTvldzuh4pmIHso94Y6pRO9qI33Gja73ZF7
wh/nrGPpa88/FUSYoQi8bfa13t2HLhKBeSaYvq48de0s5kSdr/i5xs8+AMdp4Hpw1RhQ2Iq86yfF
jJZCTzunRuFFfWCFd3+KiumajvarWNz4O9ii0AG1SEaJOh1FbCe2VRM60wNXtmn+ZjvH0csqiBSz
C52UfLTsMIDw+TPAhFUvbf8dvG5UUw9iBdvmynJcU8zHyGhbbZ5i4eAlNq6gkGuAi/sT/4UP1qLr
MkE83KgpMaxFNp4unvxWIySEmnA0/jdbpy8H04e9hL4d95oBxiJ/+NaqRJC6XLM8AMIXGggJ16Ox
E2VekZnb9F8fFderbBAnOYHzuxlV5Vd9Meud8P7V0eR/gE6omADqEoxzsBVgDXzD3xg9JRb4LfEE
bMFB49y7WqkSwSvW5rGgtoEp52vsIsHZDDo9cDU6Lg0N9FchkAC27NaoboGb+FJemCq0T8ij1iia
lIrxBHU9lijBfYjPxrLVPZ1LYdHe8RP4Mdvt1SbHX4HbietyQJU0Hr/9JHPteQOg9dkOKSZefuz7
eRzsAsvsDi04o/OAHVjDzPfrEi/kxa74F24LhmG0lwtkpBDvvAJMZBpdBWzrUODR0qv+LJ5CWqJs
0Xe5xcmfEwEong8aU4/QRqxQjPdP3uyNr17j6+R5CPIBl+NfN/kfVv2rnfltDMAOuKAaW7jF5hd5
u/FtAR3SVs9sT4hWRT893s8BUQhCPTI0EyBROI0L35mV9kURMeEZuS+ewllRbgF37qCHRdQRAP7R
DutojJR50O8kzu1WciNXEPCklfhOJMobkCd3/1fFzEQEFu82fQudMVjiwL4qgNytJp+5X/YQ+XIK
lYRbARkyujk1yXj9SDCuDrqZAVNdPoFUgw3FTi4k/2mFQC/xY6NWTuVWsJn3b4beGwQj+SoKgWNE
Bya04v9HlYki4dVGA++eohOUBs6D1QQ2cffWQXE38dr4QuPJMdROrqrTy02/Tjel61JamYJKMGTG
LW3QVl1O0LwYltZKnICkSgrHBddWf60T9zG2YJhJwnZFWFW5Omj1gdesYjdnPTAA/i5XPH1hwH/e
YA64F+CKETkCzwsEAf/+xRVvM4/A/2Rmd54mAIzLzqqdJbb9/TmR0EcoBkVzVv9RSSM8NdTrl5mc
d20b81PeISsug1NJHMtsI5z/fJiQCNZlQQIDKsCzGpFsLfXQ3XcUo2LmSjGr6sEfaIyDZ27XAyub
6ARit2JdtcmQiiyIGfO+4ivi20VcMylBmVCoef4UcYjc9R3en9URmBC0FTjn/ylEGMgSDeaGPQb1
j2KrcM6vzceUmMxCO69QTd4fdXzT/aXjo/+4wHZ2pwyPc3kpCgqK9dTJhgg9OH6PevXRnu7QkB7p
AHpArr/hj2uXZ1AH/EkjhIpnYGxnodObvP8HND3QDh+OObniTYJTlDUvpF3jpqw7aFJAh4GyrAEf
QrpZBpmXJuTfeEwrhu2r7vjIejZ0jp6YpeRHTJ1P79vsiK29pSLiDrSggtf8Un2O4YuhKuqge8/L
zMJlHMv6Z1PxEzW1hkIrh8W5PczSfbMDM3bd/3Hs/Pum9D+deFqUchcAgPcszdswDp/zPqa3Zexp
aTOY9EJq47hnBWuKMvNSI1h0+PLSLDYHEh3JSwr5q0f2YKNfV9+Kzk2e9XZ07bAIQtQog57j/7+o
bwU0ToEnpnq3lNQ1IZgq2jLL8aZvETHyo2PkqTS4OfUq8vPImwX96X7vXG5ltI9YczoJTNekFxnU
EyG26GS/vlPpuBkbfoO/digS+cWVaiLG1MR6ajhj7QCMiRJAQfX2/Hj6umywlJbDwsvhtbuAd0Q8
Aq2RbCAvWiRwQ9L5GpUYcEZc4ZnJbm/gx6rBhCuO+3MVPdMSBtHurH34m7crEMKvscFKcMQUdwdQ
dUG3iXmbwDm/NKVCwLpSKa8QVHoHjrQlKGs7rJQ5lAnczKPXY8rvqx+wL2svNsFdd8zlZu2cKkdi
kLcqJvWF/MbuHPnanw4C33K1Rt5A4PzwbaqVtThj8FiX0xRNaAgw/dY5UXGGbmzdbpcB6SUfTVuS
Wosaj93tjnEOlJ4TGT3TN6rBQyW/HRDuZibEwi/4FvYkyMHbNwdLNh31G5exFIMcLTs5KONkExje
CML2QyTFhtMhO9sy7AVInAHRrOG/UmlZADAjXHKSJrlM0k2ZWnzdpeLh8xLkDcmD1d8sV06W0Hjj
zTvzYeg9GmTuLxQFrTqBCekd/+W0c66k2zpBaTTCR0oYPTmvplFSsZKKPcoUfP73VHozXzpCrwpx
HohZrQqN9qP3+rBjhDEGWKyPMDgnCc9AUpJVjWvsgaEiIES2WaBlCUPszwQrADr1TJPHs+JpG1bF
Cs1KUFjASEvCtSaRNxK8NvldFnNnUy8N49PFPIrZ8uEwnSQwbnU/oSSShDIIjBf6z893Qwu7lJ51
9qLHWqtVUliZMfkgGI5YPWvCNFpym7pEuM4yYCnnDTkYI8alUz7vPhkFaOHQG3rxBtESuPLwRAi8
Gt4uA/tRVGgf1xtwZsG7xllFgdSB+f7D7JKRUw6hppsV5p1c2UcsjGhKiHNIfQzBCaSYcVdOGct+
PsMnqZcji2aWhBYpfDEfAYCjqz+05qkm3M8eC61Q3PSBseMbMkKINJTZAzvJ9jGcs5L0I1PRvhcr
vcJEt/5pA9X9cFt5GPknKIzy1aIvFZXSyxjVhow+Cnj5Dpjok6vIMu+yvNKfYGZYb3zDrNn537li
Xxrui9gfhCWJ5NTyzRd/Tg86H3WL8UAg1lrjeZxd/iBVyuxki6HHwaJhNAAID8wWlk87o6hNF51/
NAchH6oV3zDVfwPUjA5i/oSPTw+jtaK67anEskD3FjG6eW6a0mIQGNbJjow40rSFlBUbxLiiCnWj
PgelQ7fwfmgJETVlkylc28zt/DcbjuOyJrgRZEd6SkLnXYUyteQSE7BgiQtPGbV+EMVc93F0NX+A
2Rjk3kTEH0e9f//Qpgl04VICiaGGVorpCas1Mfp3A2AujmEAwoW7kqY5i0PBLqOULUIiH6MOmYwP
uZFiGeBcGpsGs+TZNBb8pvH36XeUfMwNuCNJuV5mA1LBrjIx/xmddFJNhfn9pJFxS6IKluylR64j
iwbbiLLFKGIcgxwRsv+NZ34aHVBCxAvrpvj4/CMpXfJbuhNelJ+htDNTCCDFvizSP8eqOgmivzve
kIM/YQHtrztG1DwCCMzayiaNONNCI18S9VM5oPyTg/KZQaqIqMN6GkcF/dnft/Tqz+i9vbMUvpiw
10xBsqTXdXoAobU0tgx0NzHu2VKHyvyskz1X9jsjWVOXBCuaxUfbtDDC6V0aacFNRUJ4dhxTVSpy
X8aqkED1v7gYyP9YDu0bdKvB53q0rbEbUdVgLOlpAnG5nQQFafJ20nZSqOrX+jCvUmip9JYkN30j
/DuMW1T9TdNRJL1ws28rRv37Y0WCEnfvvOVF5wXByaa1yMUxi0l49iw/K2XTvrq08XmNNCcfvija
edVnksgxjJwdp1D851DEjMJyXvQrsXEiaOW8wDuyHd68hW3zbzboMMKmpKE2G4R9ImmIiSaWoOK9
av5eiKKo8sc3wWCHmg/gc81XObyZB9ir0Cj3poCbJiUjOKbhxSr7GYSqkPYb3VZqKXS+R2oimYMy
CyNXg+/71xA9wEALtIcUqOUhhH4FbYW26whV8TExqSRkwLyFQjAO78Au9qb9zXJrM1gPotFARlhK
0trYB4kwVgDSvjtraUXEdeKRww2cJXzEwUS150ZWv1vFLdSOHTfimdFharAtx9p0zZscYULrod8N
DLuwSlKYyM6S/5Y3PuO19iphvSE/5XotXos5ylmrlFL6xmK79u8YVtdQ6hyL1ewjypNoJUzEZZ7I
R+JzlWF8IlAacBEHsOBHxbRyh6s+hag6cE8u2ACj3XZDYmOphsnssDneN7aAiMhzMhiKOx1f1qhU
MDmcxO0qTc4iE525Xa+C2pOA8pIlAH7phHkcZIi/G57whGjBUXCqkh5wwnX7YGoCL2calpcMymO6
LnySUtlSFzdfLUugUB5sFEz3r6WmUGAEiMaUnoBtCH0WefyuqRij5vaVflOFNwqe3JPRzdFJ1MoX
ffyRn5SFgn0LoL777J/d0UMf+pzInrvmCwKYlOoKODDzeyJPO4Hs9t8LAH8tBQ4jEJ8OEOHYSgnU
VJq5JQBVmsqeJlo78e0qLl0qTVswbGAsS3XVlWh6TkT7slqfAkcUYdBMbHbDjt3TX5VTaa9mDTbe
zBgstiWg005KZknjTiCUMHw0sPNpS39qUMWFbN8GwXQeq7T84bXy9AK3hXYrF8bYySQf5g4+kbwA
vo/9sTAY0qd/fVd76uV5/RElS9pzocvHmrDhDZAHxLczBqDD1qCGQJ09rxFbLU3Cu2XhIGmXkg/i
uc17IoxerC48aoBSxO9VoDAoeRfLwa6/y54NKUOcqrURM0/eFKUc4hWloU+HGYIfaIKa2pL56tJl
9fg+uh75m8U72fl1BpsL+RdyvCY+P77EHBNtI8qD5+oH0ZI9PcDoTHyq2+cjke4ngTHXmotHk4uX
b8d1JtaSBs8iIaOMH+SKHtpxcVnaqSTxb+PBGIWhNjQ7cUTKCxENQGl/8zZP/KL/C6aF4L18bUKV
ClAZ5Ue6dtX+USnUT2uZY7TvWwP3dzvAgCwpVUotxdsRMPfM3tDNo9znQ/LrAqwD0eGFDiKEIbFo
bGNdI7m11OaUv4FgM7YB3+mvhFwbQC6YG/PAGl5hebFZ8voEobEFhoRVc1TH2oHCHCtpo0c0ifBv
GW4I6OqGAVSTYQ1Zb+3gd722XhAoL6ebToCioURKxiohZ2/1uhjJPL+sN3VMffxrVc3AsadvEtPe
JfMSqN1JyWwICk3ouK467lPoPen+dkkt/y/MtqAJ1vrpHCvC6xHveWkJ7POUY9sp6vvJrLcbVbUS
ICvA/MHeix+tv8NsdzoU9yRqKOPTaSrUoFPIDq1ShcuUkECNAhWCq3sVGTNxIinL1L26q3yoHqEu
YlBiuJJAV02EiT9wwuVVK4BFiXnLkp6IkTfcvBx/SjIKGh2rtyrVdDAsfjP3N7v+aETQyDGQKxPa
9k8zHDq0aUpPWkzY+w3Dl/QReubLr8gWqy5glTRVZ50UdIl7EgqGD87ikqpCrAhHAO0rBYOfg7Jy
i5fCTeTDsi5ENmXU0cF5X17ukNKY7hEx58DdAzNx0cU08D2eU3QPrjkblUNs6RmdRFdFLxXGLsXz
xPldDs/lDL4R8YzNHutdIPbOW53mv2btsoQWbG7vwucGw8T+D+KO7O+7Mv+VdJtn3nG0JVCWhjMz
Rw5Cv+eQH3HKWAFQX8rVyr2ea+A25GN2lVbFMh19AWa0jd1w0XqoZCnIG4nZk26FFVYw03GVZU8V
ra/pDHtfJoUmgaJZMtzyPFJWWeM9gdzhvGc+gkFOCO0s3Je3oWOJPByYZMjB3r5rPSIOzgp0zuHY
tN2cdLDnDRCJGyGkgkWOkVcl+PL1Ul9YeYXV8ZssoxgRi4/ydkbqjOkDGfc2pFKHDF2/S2DsB8tw
TzK5yJCxGLbl1XU05d3KeUFmpCL2297mhMpg5QsYvL4ynv0iddBGfPOb505ve/1v0ZuCv/82JzG8
9hRmoQMCnIXw/0/0ZKAgcdGv7BR8GKBrv4PSrzp5r4SMeMXiKLzLDaxOyeNdIMtnMIAtdU3DMfEC
4FS4f0txHUF/Tnl8D6zD3TumCRJiws+hzPdhO/yNlS5gS1s1JKqVtvfmSkM2D8Bmlu73FziftWN9
69Xg5D4DNtmND/eJ+RjJJ0oNdqSPvYeNGpv5l+3U1/CbpaiABQlL9Jtu+jfZG2INJDRGu8oFtPYn
1h6dS83yvRnX7r9Xmy+z40cAGtzGkdSp5+ie5dwhjEc3VcoPUQxFtEImENjdXgXXlStPqYnHPSlQ
p2wX7kdB2GX3MwYJmgamfpWoSQT2SqNRG1tdgr00Zl3LWjNqGKBFUsKhirsaoj94XYJeDEukNBN4
a04IrS5ZUq2xM+3zxBNd7nSdOhuIKpsbjNQ8Y7h3iJLsqSkphRmer2oWbsbCfkjOKEcT4RiqMH3i
6Z/qVeb0qZj9dKuoFpi1eEHHAo6+WPtRG/d4/PlZdmbwBMN4bKfF/gXzK9l7xc68rOpkaKSfy/+C
0puyHujlxDBKKz7gsfXyuA0ZWGf5jnOKh6ypkzTsQarOTx3wARgyyMvbfjbilho2PysJJ+KlpYr/
jDtgS+NZRL6wucbkx7BA5fZZDE9iong+mLfH1NOPLp0MmaBKWdru97QVx/iS968IqjkGnjT6mMzs
MnWJ1PZ0yKaWUH/9nF1vm09fvx4agrJRU6/YlzZ5CS8sR/BAb7qzcvaICu/jxk407i0weC5AonsS
7mfyksFGtokaVx62BnT5QwxC/BRyU4AtgpbsHf14YayPKI1oiPj4QxjAmteVXlYK2sTk4OoGgNAA
4LMYP6CCIf/AGHc51usf4o2GgLoP3ADpmXPLFpepwDltVfEaSoQYacGvWtV1m2w8MguXmhxxfEqL
t4WVZ1ZneBEnHaolPibR8WdgeezGRhxCb7NZA2dBD4IkvL/3JJTie99ckm4E/1eNwve4mF91N+X4
bLme/luplpbJ4iI0hKSaTQnSgJcjZfpa3rQmhRluPUPUl2XysnrOCyn+O38XY14BXToWVh8GlJsr
XA3zAknnXvWFPVfJlfVmJe/TY+JIdL9v/W3IUwpOOol+XK9Fl/kEpqu+mc88C/5M80X2Qf0eeLG8
XHU+Eg97Aa++VNyoMfCgEYJbN7jyg0vHQdEZUazo/RhkRS/mGfo9zvD+hH+8MbOgv7BPBGRVVncq
pvRK/AejRNPQUnnJLgPeOafPiZp7wDPbcqMiL8ZMXvb5M0mM/r2Dk5nK2+diaNwJFv3/pn3H0v/d
sKVJfqD/7zoH6u2Pb1+CNCX9SrHw6P94uzxCJ3wTdHgdS/jVtul5KtoADyhe/TILo31R/eIhL9k1
DeNgDdNUcw8VVNkHVbOw63j0IuKzGjqtB/8ga4wuQjSppVzLg6u4G9Ovq/AVB1RnosLDmMVK7k8I
R1kNihBKuHp8Y8tVBWbN2WKQcyfN33xcrenk9NJeH/olQH6ci6g5zgqHCzcKNbeyOLQfTTIqiXxu
tuv827zmhSkNni1pp/3sLW7P6ni5eUa9pOWPh25XtKYFMuVPfyBzYxZQHxhavUmotTN7pMWcRjpi
Y1zAUNIZN+DcBMpiu9oJOtUnQY1CGNwE1C1OcdSq4awYYlXTo+5zirPGd7ckNkKHr8e1R4/RpQVl
V3wSao7oSZ8RdeL4gCQHqinI34weNBhRN43ue0XgOhhbs5XK3ybRY1H7ljj37og4bEWa4ZzKtmXi
ah5wePFGR2w0PLbzHKGX2tAl4Yqd6fuqYQg3q6DrsardZkuJbuad0aUqJyemax6wY8D/F80DuSVO
0hotqN5JOlXdLrBzx9WniBR5F2pq3bvVBQ5dDeKwK9KUyQso93m66hOZ2megwtC9t7ZgPfWY4OS+
wB5pqevMpZogzB+jFt0H44W8CnW0QIdGCw4jV1DoneAFkr9GwODfNPtVlurst7cgI1BeVOtKByad
dQ/rxcNTT5gL+dJRnlOR7kAxaSwbZ/BhdaAtxbXTFXW9DC7pFITmT/1L/BmlafQeRr40Jm3X4P8e
a+3zzl3uTpwkkbuvDSmYRqTjBT3FoEkeVgVZv19yX7RCFFeSvI2RLRIOrM74oytJMnmBYOxilqYY
vActGxbTYnqbn3gO0gYkmjfr09XP9E+sKe5XFRP7aA4UadI/jVCQe6VX0cJONnOlASmBGjGNJq9J
48KCaPrUlrRL/62GQAVJNZF4DwKsl9BomT+cX4zlVMo6G2OxTAvwNJx5rOVEBThW53MQoWJtJDnk
VGfVfs5AU5izyK+8+oXRP1yMrZW6bR8PzMnnGgcFy+VpwMiWWQC8efbjKqgd1l/kB2FO/C++RJFU
YzGAX1x6+G8s04thAQ6VNfSY/v5ugsN6aCg5NylwqpCna4XCACO2TFbg3Kwxu/bo+Zib1Nbv3chQ
daZMo2ZKPM+17wzwwhVEBC9dOWCy+6Ci/wzjmdrxi3HaHSylbQvlnbctqaRHzAIpfLHTaaO1tl7V
muxoBQOcolF3JsyflLeOCHP+0NhuDJQ9tuN4AzIRpiwYn9haR1unyPORKpqG2XxRHsvdVS7BJLE/
A841MCpDaKuOcB9NzOHPXfT8Tcvxj9gL5KSWUV7sIbXN+923Dtt1LWfjbYssycoKt36PYMEy9p2v
JVusOGiiAhNq2r0D2Rjcz/dJb1tq75/IhtPzNVcfRqDGU3Iy7zgsEAuMq9q83rF6iMV08N/ZzcB1
CHubbGf16Yhes0Ycg+d33asXde2Ah5Ws/1H8miL3yMOUOILFeki21EdEm5lUDJ/ahBCfdQmQKMDY
pIh2t+0TClYMiHdWdtBo/FW11OGMHGTg1JICZoC603MTbVQdZd/XfDklIune3lxRf3NjptIEshah
Dyb9iUhc4OiDelZGmATLG607VvKTY0g+PWyliq9jb2Tgk2GXwOMjX0+b/2kSQwebZ6SHn2FrbySn
ejQRCNJeT9pZHrEwl7Ob4n+RN45UsgRSn9ypTrMC2WS1Z/GGFN//lm2vtqoqcA096ARrDJQiNZ+e
nR651qwLRqlh0UOsCEdiDaAkrzJ8MD/lsXciLjIaUV4HWPcqGTe5icycr7/9HIDUFh+onTd2h01J
k8uB8Cp6vAJqL7e6CSzcqQ6fpcZ2cIDJzvZeBFI3EiJvmGTvAkh4SrZgysME35CnsLLVu1rX700Y
+/9twYJHBFUKgyd7L8ggWS4G2t3nC2yVrCopwHwv76cc+J2W139bF2HpArr3kzNB9DQwpG1u7jlz
zCOqf4LTnm5Ybaej+L1R0csBR7Vkep1nZBxpjC46HUY0jbhBD0fTaCr5TKr9cj5Qo6urityVb/C1
IHahyd51iriSKCFVw1opboi3SRqIvqieEMLOMBBLclaLCvQnfiPQhB2LKHMMOYMJaiVlLNpmlWha
FK+92h/4SOSlzQbyvLKht2CPFen+b4V3G+ePD9//xKjTdqNshGD2Ol+ZYczty83W5iIInW/bA5cu
lq9M27/nEO1yMbAugtXA/khSAXQGapErZyd5zyHPzszSXLJ77YBoI+2RR0SF1ac2lGYT22AjiHeH
mOwqQtKDb9ec/Ks5rtBwD3HhVfcO10Fp4BlCS8Nv+M1m4cgXKTuppPJn3pplQF/zVUJfiyk7Wc7K
PZzjcc409UNquy2mc3f3oPEr0uw4M+eEyC/Grt8+JkzXhCE4lOLkQ7/o36dHC8GkAS8TDXosQKz2
CYomB+DRGxWG2HxMGK+nFHeXrMW+l3T0FmpC3MtsU5t9K15ZbdhbNE8DCbPkGljhTnaHvPPqaS8W
8dq2+1rowg01TvZw634jNNKdjeymkodC24gbR1ywk9UjUKAK20SZptIpATfR4RB3fUXF9jlr33im
VWprB9yRIpoePssYi8dklkXL38lzlUr/VMxr15mQt7sku0bTaUlwXDi4azBHRv6GZUWy5irEokVq
FdSmseyXsoOXd8U2B/xp3qX4UVDMg4vo4Ind5qOmS8Wg6M1ouhl8sYS9T+sVMX/lNa78+m7w1dB+
XB6M6v0kwwPYt+IiJjufld5F04fTFXlbhEegBUO80yfQJDBUkHPhIlXXRK/Gey+h6+9X0+8KU8sh
lMgtoWq1FdNYcbWyiKym9lK6/21U6tFhHQKgsrgjvtA2CfIZqy/h/L6Y8JqSUqA5AkoMAVWY/ql9
UCNHbRGeJNH1ZOGeX3hmz7YMo0ZJdbiGScYglJTxZipZbqmW9qpFus/yS+2jN69LETgOla7M9SBD
WGU3ceAp4bJLQU+g2WI737Tdv1zZeQKRmLv4C5oFNUsv1aZcqSasGS951rixxfrQp+pXJsHXLJWE
OXILZRzYwJYeWyiS6AnZPIYusetT8P+wSODlC4WKS80Ml3Xormpte+ubFj5hEosfBaDxYZc+abPD
LDGZCSOzuygIX8E79akJ8Bx5LPXc6K7LGz+eZtJVzh1hHIeImxbiztFVqqJHK4UJUBlSiY6o8y13
kjG1zEpAnCRh80Wo2/pZlgqStSZ9ZZb/DVneyFRNxbzL+TwsORK7xFGgt+LqWsG2iDaBDGkaq4fd
dofqxeNW7/8/1PbgA6aVqIyW49GdLA/qWhGMb1ESU4plQ+hPbdW9wHsfxF4bzWsQNgrjTt/vGzFl
3taEhKC7xkeJB68miJoV5Jblf3e9cB7lBYwHJNKILihDXesmda+U3Ms/we7IAwkHGa+6ZpHcJq+S
frGhuvjyMOIMzHdrtEvg+zgwMLj1bXXVfqusgPaey+1NBLoOmr8Go47F5G3jjibliybpVqBBb1hB
NrwYc7NgFNQU3ZheMfbzvbfyGRzfxeIu0cPeey5DjEwkx4mPmTkhvGk8F5vbmZY0hsnKBvNaY9ay
skHv5tNFE8XmlNeO0ioQysT2jxUsDJpNgjG+rEQsaO3nPjocjFe3/M5AjdP5PLAp616VZMAOxBvn
NgEsLhZP+J7HC80xLEu5LGNwa+c3Q2qT4ys/6bkhRr7ELuPOmMur/lULHmFSO/n/8QtagYipuFJH
V1tMPqhYehpJY2EMDna2N+85Rt+k5GiaB8Etc+2bZ0nSNHyWT5JmNl6UmsYvpvpSwv4cQeM75iNN
cO/uXVMgEyIqh24yyClz4IkUNGfRtCXeig5YnLCklQl7z7DJi0tfMgnED9OB5n2m0uDrcjCljaxY
kslKkZfhGXSmcnG7MdH4EdcMC2HtVp5uGmn4hXOL/VIzpHOhqs0BnQPIYLeZb0k92wZpBB0J/0ii
5IbQPmPF/zuHwWoRjPtA7CLIDW0S4448RnLTPswboJuj5b24huDF6Nu3ub0+dV7oQ/Z98AAqYkOm
cRNcp342lAX0GNz8ZXkX0OeOUNGxrGI/WGQuFlf7CUnZJOlzY8f8B1c8urY0NoXBNBi8D89Y/XNd
6s2mEyv853zJRBREWL31MlgPl3VKeE237gpVxBhAI9VrxylkXffpEtNDLG+wRrEjWCExtL0k8cNA
RZQxV/7KAY46efa0wSUdeJbws5Ih8o7orCh+MAjW17OR6EXhDfbXJ9RnVxLZYpKXCVocGoI8mK7f
gT7NU1bealYrF3Pw5SzxaH3zUB0uRkZT9k+/9R6Q0fvxYzLU1DjMc+YEkQENLO1duFU05UsTTjn3
Qapm5mKg/xyFNZZlcnQrIlUTFNVmOG1ggSJpjKRSyh6PstEp8AjzFqMSWJWNbjDAl/ay6yo3bOxT
ggBQ7MRQKm7hDdQlgVOrvYO6aJ9uyBAXqALc/Rt/G42WH6vHcV0dMQQS7xGyD/qwoj8/uApV/g8f
pIJaaI5ddE3Cf6HraDbapJ54aw1ZCuL+S9xgn4z33w9xJ++s/8FeSiCA3T7VqQKcFzmnayjxP+qb
itqDaOvlaOTRVfWu5my07dV7Jn2txckVDmgAhoSZq8QMvPfOmraWPtWa6il9/gwZOM/mmGTtFWu2
hufFbSZu38z3eJJVzxzlwWcK0fDtzm2HYDhm8HWs/wkaQsg1xaY25RqL5Ni9AGDdH9sjuzwptIQK
cCbWxYZh5cX4uzU6pjt9lnX4paH/bIn6FtFW9L11XR4j1gHCq0XDMMhyHOzZRJ2pEghSOZwhMd8s
QHVhwXcQSHJojualy476CiXF9LX3546xGH/BvOiGHS8Mm8D6LTkLVHWaKz+5nHQ9/xiqvcQV/KKS
sRRvvUHmhjV97GdyB9qe/XPAYhc27uIhRh+XEF3SEEllYzZlsB1iIvkAwLYt/a5qG6aqaV2W7Djl
RdbZINhGiq3j/xh+qfMu5mujJhR3/0kNF3KeKRcha8OPJtiK4iVyqIhBEzW3H4QdFMMWEZV3+99J
LZtGGcNom18+kCSVj4HD0Cgwv19vUIesG6CjPf3/D4v1Z+KtwVsL0Rb0EAWJrpmXQtOllMXxHXhZ
KewVMo6wnfIMtxXm8jdx5WyfcZ1rThQMlie9z3mh66J1GzwbCmPm4lrZ7zYLB4K59DkyE3b9rQUD
EaDJBF4p64JMbEd8XP5DGha+o4xb/8UZ2wz6z0cdkpk5/hBWItTgJXIYvFrE9TWoHzngwLuuLUtX
+IOaSZgzwuLN/xk0s6o1+o+MUaWQiuXWeVr3KgIcrPZ4WujcCjfqRsOKOcyVLmExdE/uGkkFIQYP
vNLojMvztteFR+3rRZnj0Cg9PWMfVHpuTVjEKvwXdfNAKatcHtAt5QFDacb6dEjHxIF4PAxXjakH
cPAqN1sdDRIm1vhmSlqcxD5IRlRPuSuO7YVRtMK6ioMwoFj6mxmQWe46sEP7SsLeyz7fxCQFmeGC
cNOztyUZguwxk7Rj50VegeM2faAwKE1cmamVImXo5d5CuDjqJFuriDmKPHIEivO+Ukoc+CVc+moB
rqzsS4IqvBLC8dg5Dp2ZvvAOUTVZyyOLAnTUAu/Od2dGK2JgCZfoTUFhcMd8FdglrFycvqpalr1W
4eAQWY49PY6lPgYm6bLLIUIud1OxApKAcFN6JtyqHSd3qKzCYlsHhoslAdIYSL1FF5yxPn4J5JFx
i0UblRBI0K2yzkTCo2RbxhsrYcE8clXtsZ25KpUozbmvPnem34HffD8nV1UYYO1LbFadQUxsF06U
0sImUk4CjvDC7++XSGrVYxSpBikFP8LOabiRRSpGx0hSTHf0QfVF9ino9dG6522ytG2YqBQ1S+Gf
1FAJA1qW5LT+6zOjXH2NxisBRHE2cPl/o5fgJT5OD193D9iZIv2dMUC5IQanwtDTT4veq3+L2oCo
D/pTKesQTSngFqUMa5q2wFqppBgPgjjSXAayytAUTNEg6q7RLFWXNiOhIBRR1RpVYSWZCKpyQxa9
61aU72qvvTpPHqDeB28lwQwosQcOfKrASbFbvQrk2h8ku7118L1DNQ6/h71UOtDO2o4tHyFmRZ6U
QatSBd8j0xf6RaZtOMPPWcWEtZYMFUJKAL4NXAOcucHVYSZsfpGLDft/mMjpDnVuvxX5Ts890H23
kg5ZmbSkCv3+/Nhe35l9Nou1xt3Oj7qQKV0G41EnvbSwSWXzmohHoiVO28pwokAD70UWcL4B5zGE
ljKLV4yS+CWwpdxEbc/qbEkcOvw9jFWlypbHyj647PgGs83v9ctZgAYh6KPp0dK+9wlfqTqlwEuT
Z/niE5brNjCnFLtrJctRT5zAYMH24voZkbL1G/Xgqs3N4P9QSwhkMdaIkcoTwn8byWzwTlu8HqsJ
6ajUUOerX3HtNwo3I3GBNVLnpegALjkwdOZmnZRSL9wkGo5HF8p9nmHpPgvuoVKaxjX6X+AVUe7p
ME7W5UnUX+T83xJXXYqyVHMmsF7gfbceiJ4FLElac09v/AqjXkrBezkZt7t2PiKyQLYU7KBHwhi1
lyPxfmph2zKeCt/C4IP6ft8MihGzhemz7W887gbkozZi/AI4bDcAmlZH2Ei5zTDx3bQa9a3fHbbm
or57YmrFmGpxQkv4cvbO7QGPSk9Qnsk5H9RAnfY4j9eRb1clJrYYAZFyB9njzoZW07LMPsfcgK3X
dqE7oHgtWtof0lRPIBf2lrrUuhnuBHwImuNjgCchs2ZqOBXioDEBrckrM4KtEp/xy9uvLv4262sT
Vg9TS9Kzv2wFX3pSjfdyZSAIqnfvPCfuUMwekIqEOy37+V9q1MZW2s89ohmAJWpI/kkxEg9dNqJt
DDdrd0a/4ynuy2w/d5X/rboJQ3pBZ4uIuHJW52QGX1BU4NeyGCalohwDBhoY10fNXFFjncOcV2lW
QhWVpY/q+8dzBquqKin8MRYzXb9A96LVBz/O1lvlKYYTtKfD2iWZI1UD9C27safmPPNQeaCGNtEk
U6Ifw2aC8RhqoBLON5rK2/z5IzfpvNEBLEOCWjKwxRV0eHuLzC5ONUIUOWUv4hEGuQHUiBXCAxc9
n3OVVVanGVjGkI+ETJfITgXnZwRLlSgEUNrL9wm7Ss6XdBykW/fby3hGzMkiqOx/BEDDjZt3Q6DW
q1LWHeF2cBB911y3jh1/epS7Fcet4O30rdW3FcltfBp3mVJZQGvisbCjPkyBzvD3h/U1K6+w4q6A
HN3kh0J8zqqpxLd5WyD88s49yQvhc5CXg4J0a67k7GeuGLkq4NcP8wKtCzE3H8WV48f3xMI4HXMU
iiHT5Si1LcTaMjvhzg4fvun/7zYaHgZ1YDF6BwGwW9DT6m5Q6+UfglirvR6b+4m5m0Fau5VkK6dA
h9B1JfGakPQHiFwzBr/BwFMyfcK3YNqT9krhESyFur6nWWjfDae54QBAMSAJLieQ4wyDKbv63MK/
R9pHvsSmauIQfv6C/LhFk5oH+dxarBa035iiLGtqmvreBxFGLAuIu5ja2BEXvOeuGe7tm2i69mIn
fo0vJ66bYlvQgj7ZwqEnegKAFrzE88G7VMnSzXxKEt0DDSV3U65Xx0notkix0HA2gQfFobAG2Lsm
K5LmDGReuV8uOJOHGLbEzn9g1XJzUA0ccKwdwTb4kcONAQp/WnA+Q75jtubEhtzyY0iFB6XIn6q9
KAR22TpQ/YGBdDF/cPWRaSQwpyHaPRfeE3vkqaeWWzPXeUpI74T6mb4YmrfxItEkFGt85aPUQS4M
+u0XEkMrockSa017FK5QbjZn2bjagGH5fItqW4aU+WC8NWSTOOMpwKrCvbEEKeJr24NDcEoYbBF9
YCPSYy61UVD6ZcgoWeQgKTNyr1dFbOrnbmiHOSAY2M2n/HGT9JYt4FImV0OskRDCLzaQVEqaI4yb
LY3cEBW//j+a/1glzsoifgrOBEwVls8NqAoB+sHlQtT3A0M7zadMK6TB0PEqFSEcByWN6OMd/84p
tUKLWILe4W98xusa2feQ+9kvVS34udlV/5BSn/ogL0EbHudijd4HFr8gIZGQ8DXLEsweNlK1apVd
32xXzJgTcnT76tkFWCKfIr0/GwiSXIGT9/TKg29El3StF5e6wgTZ3ZNRLAgDkMraaAMXOYvGpZAj
I3ZqTxRFhd9rYJUoUDypmeP1jT2QNweSb8iDxsKzGI9jPUbYIzODVqHfaQ2DqmUjOV+afREQdiXY
J0oDbeSOADg6GCwIKQntZ0vOMp+e3tM9qT69l2O46y/+3SeduvVStbSRIAKBaY0Qbb/IqJ4+1Tuh
LS++oWve6Ff3N434XlE08HsRjTl0aaZXVWnb4Vuof2NN1Dl0aqodOMqU2INWl0Vf77WRbJEFB9Rs
P69HfkN0uhSFr4ANXEUaY6n3Rjjtid1KgHcVwFBSER8oklPZLJQ+Io1+2bH6sOPn+fjHNQNCmTv8
AxCyQcC42W9xGpJFBwElIx8RWh2pPBdgubazmyD5l/3UzgrpIaWj0bbidIuIbvIRfsyJNqCCm+K4
eAkvkUugFtWKETY16G8kE4qFVyGxL786r0OkcW1ZaEJa0zdc6knYWpC7v25z+WYo9N0SFlw+I1AU
ErS5OYESRqCHNsSytQotvJLom0IAP/jlUlJgiqHRN0LVe498AcYGX8MBffZ5WcRKkbNuiJE8LmXY
PagUZh6SRf9mkb+TWFHOl0iLeYhofaYCffoUsIK6Ml+Bd8DUoahFql5t+9wUPEfhGB6dbGoJOq57
V8YTpL6uTujRLRGxPog+4g77ZTsrN6GPJ2kEDxeUqk8IUIg6suwk5yys5pzn+sVhFPPxYBDVxKUD
x3pBv+j6ZOwiI3EdnA5Y4TjKuOwDNCzKmn6Q2Po/GYvt1YujPHh5zdUuT0W1K3LTcS9SvlekZSl1
yZYYN3CnAZfep4uGpRkdVwXN+ykDVST14fjiAFL9/nkK/qn2kTCcYEcTwAy9BFB7Qhtkqh8yCfYk
xdKXY+ThcBrIGveibsGsL/tO28LAsOAqCL852VN88TA5BH8d9mWi5C2KVshgzgpngFIMPNeRUBcd
9rr1BJqx7sgJqa21dsChs+gQHL9PPdXovZy0F/7y2DcdADs5Ba6qpMJMWuFTEMJCwM98TcQlB5kj
S9H6sYBntGIX7E/Qbpfpl3vpnFbMoa9d2qK9AbzAd3F7ZBUag+tnUQBxj9S0jzPOjyFYob2c9Ndt
74IEqSVQbXG40e6DzfrSHobUiUcL60vKm3WQxxfeYpgLqZVifI4IxqjH56F9drDjj84lnV1aQc32
VF+UkA06UbJ7m5yaHw65Tt10wcNJZGaDD/NAAPep6a8KbtfmuFB3Fy0fPK93vW1V6vWvniRLJsVx
03yu4NPtFZIk8KTdk5fKPBF35PeS7fLrThShLjApSmxE8+ebucc16BrJKP/6iLpPF0+gKkxt2Gf9
wLWFbUTwbn0JrOrH8l3X8zpBHZD8LBMNzpPow9DlXlwNVSGCixSWkg4Xyar2l3tIcxEulvIojXNV
XzlgD5qcU66K9ULg97g9sS/Gi+YvgLlsBmEIbRtjNfEO3AYkbZKmQUbp9G4xSlCmhM+rQQSXermB
naZPbSbcx+u3ahrcGpcDhXi7HnxFv0N28khFvELxg5CYT2IZ0W9xfpSPYdY3Ng0MutsUyg3JhUK+
dEmVJq+UOcMsFcvrytxJSecZ6MDW4mv5RSD7K3BUNIr4Fq9uARNPEg7az2C+HpQTqRV6oYbWGfFH
Xd4RYY38bhW8lZ0tkK0P7TpUuAlRpsK1ADqm3NO88j56sS1Szs2vG5eNdovEBfYmFBw8U9qREBJ9
pv45i4gl0Hm4ccObG055C7BhHy5KKixF7UAh/o71iaX2Q5rHtGGPuNLKpwhSznxIQ7HTl+FCnfxW
5MgLteWRJqeTm21kRaQhfc5vZ7NRcHntTniMe4mioz/zqPXnvaBvfZdDvGPKrzDC5pCjNilHi+pm
bZxpcIbI4w5ia3z5MB2o84/YEuJWIsnbBfc6KQLjiF5w0smFK3WXJul63eXvRcpq4c0s6l+XPE86
fkLfY5xpLxGntThMFDyht5kNTe0PbNFj/H8dDV2bFqKC86IvRnUTottzp6rR0Td1qhrT3HEvTZXs
EHro81Wv42Q2eAon0tsEhyr2hXeEqwWWsegE91+RQ62XkPOVjEsqlbpBv8T9VXJacZdjG1ZCucXd
B7eat3ElVp1HkpsFlAKVEDjW0516GoSaDZKxXoJK6I4jDWRuDnBlrckHC3ysah7pycHf7FdX78F3
Rf1JvAHqV0TfZaVEXdKP4jY8D0PYx5/YCOi386NBYj0fXRg7z2TXMoX663HWLJpQ1eIydgsQSZEy
LnbLM59Qs+tuZ9b3FCn809GFiHfayx5YVdrGKFpYilFq71oAcQL+IaHZDPt2+eDNLOq6CFR5hpRB
jxRDsVzvQP88kLIp7sKLyCZ77C6gDTrJb+19TEeqB/3va5PCugafW/CsZhvqmjYxeNAuepuUc9Hm
WJeuyOTyVLdvxuOMQ5AkP1JziYuMtibUpLdWO6oC1ein3sA/KOgqZ1VPOSTZEMNT00eXp7CnR92t
gSz4fRFSfol4wKPvCVBOefUtTjUpXwcvKjRQKF0YfbSVY7RY38CgvpKfAgnQi772y/GzTSdEnkz8
FjYJHyj4ao3ThS+VqLNa17rtMvpSCXd5zm/tPy9xLiVDpdlNNSNQe17SlSPHyIZm0Op4Un3UvRk9
vqMdJHXsYgXEN0rOUXZYY65L8iWDPPQv/TKCPzknjpfqOeoUhUUP/lk2amOZ2LaHnYk+ObgdqyfQ
V6Y73THcHQFB/498ZDACJ8v/fmhHVM/vKidGOPwXTE0/Su2D34Jbhy03ld3DxU9QNq3T4VexqeY5
ynihFdQx1U28jMRa1smjuozsw6T7W27mOIjSQ1B6uRdGtRyvxaFU5QtpJwsviEGqN2uErExZ7Lpp
ytswxMUecZunHV1d86p4DxMcZ/9OFBODnTG4DLZdFD+ZPs41Ijp6qbW6h9AhPBtG1nyLdeWxH7j1
tMCbIwPLAQpmekJ8viBD4ejy7mjbGmKqf2diyZrgeCxVwWztN//17cM2U6wwJRbZd/msbi6+492d
cErpjLHPzbyfxoTPvBxw8RICulqNhWQ21pHMT3A3120Kc6mtUizSm4uwexVXjjLVWg431tXrBDQk
84IkMZ2f6YSdhe/tZ9Jl3Q8iIBZkuP0+owbYb/BwKHZc3YqtIVzcH+jB9wnYW8dhfcJhOXyFOjQF
KNdbGvx1OoDYstlwV7qn1aeWVPkqT+GyO6eTWaaByNeUE/Pf+eCQnCh/MttsNziq/+nJoRfQicRB
bzYsdQ/J8PK50/TMiMkPK4HLGxp7P9Kz+xdWoKutCetUQYjioeGgu1nSTMEeqVslAM2NFg3orbsE
xwriV95OS25wro7QYNmrpdnFNbfe2ekForhR6fB5NpPRbR4V3OY94vvaIfHFOnhNPTrkRh5wZc29
Ds5R6AZ15AnfW4oC1mD4Yb1a+Np+9NWN9IMczYKFedAb3mu/Tuz+jbqodjanOBxnDz/J1UHzsGb9
b6vsE1+XhPHQL0q1bPw60e+gY1xtian8GJpgm6cgO1lSuQbMp/dk6ciiJT8RAwAw3Bd39mVXz9uw
vQXzE1jce4cirRNWYfXB+nMvCPlUfcB35Xw0DD4sSlOYTHSGFN3vVpDPg+08Vikz03bOhXt0AvjE
P0tUADZSmgOmwRbsaf/e8sZ/icv4pmcdf84sfK2C/crLkP0MrIP28+dEz7F04Z8PmS7I7Yv5d5Ed
a9Mr46m/a6NEvcm71tVXw7ZRHsV2Y0u4tuQM19xNLdloSxDEksSCiacFJ5I02LNCqagikSbjZ2iP
sTPCgUhaKvJoMPSi4Qes3OMrcOcwC8kdgngcgwnpwjX4U2ccYJosWjZRuRwtrJuikJdUq1AjK+UY
jINQpaaZcgqrvZCTRDrE2u9xdR38PiOaZoaVYS1ch97dD58WABJWlYWdiyME4N3OP4eno2ubklWy
ctxJm4+1wh4HTE0uAMRyqw0+3acmtuXhGrKyru8DTqKHKzpEVbvzBw4ofw8IjrnYHfa7gJgUQWRe
D4YDldS9FgJVxHM30Sl9hFsxEGTVqW5hCAQb9xVWpZbBOyE98XMDA2S6AO2PZjykyPOSf2yVi5PG
SZRMNdmc+5uQug3EO1vXiQK5mNZYgKRIgUB6Tm208QMZYULHHE3lgDkI2jouYCdgzx+tRgRy6ft+
U/kIXMfw4su8GLGvuqYAD7BEtvJWcSxB+VW8UNCVPov1oS8iO7rKkGbyDhIT79iFaMVqylhAHK+D
2B5Qm4hae1qyINXYsLSXY2coyU3DNa7rbvsq0DVcdMKHA1USjPL67TZrAx3usO5QZmxhCtISpk/r
tbelU7aGzGS3XsgsxIqrkrv+tyokVrq2tRBYyxsJkBuqaZ/q2CsPno/znLoNgevjjKLjhgms/6nN
67K7e0Gwx/lT4P3v2/h9X/juosIlirHpbhAuZTc9o8ws7MhnJovRaMXVW11PMeRWJOruCVMDx98G
wCwVxYMhPyiDJaVSfqVV3D6WSONXW9y6WsEI2JDf4jDkh33UiUo3zvuad/QB+DSXKWsRO3Cds2dd
6NGLQcIavAAzZ54CXYuJVA4FxMbNdqj4CbdV7w7owGSxZi3PtbsSpNwQhc4Hct7UeP4MMaNtNO1D
lQ2ewMxMRPSgTs/ipIaJ3wsZU089BZOvU/m9LG7c+wtcnmYM3R8J2o0g0F4Yy+RCzptG2/GpD7Mw
GJfCkwoCdhLMKHkZ7VJ6IhnfRr9HnQdC4XFNgGZvp44QWjXedmf9gU8NmlWmXm8ihiXsru4KrjnV
bnhNvJxpyt/V4wx00WnRLI4cD2wbQSsaProNHdR0qG8psM3x0d7v71AEwUm6EWTrrPTjL24lLKyd
C6s68VzBZ2wW4v/T10D3MOPQWnYSYPb9DDn5hLzshUgN7+PuzZa2jJylsaJjENnuJfiDlFYh+/6c
jbgeWQG2zeRfpi87P8oAoaSRJRYjkUL/LcjNDhTqkyb4dXZ9lFdKR/MfIoUNeiwcJTllqUqthr69
og5mwZeSW0GLElsVB2pqz8Xyss7XZ8M77UuR7sq45u5GQ7TA7iafD0F/RupJNnSHxGNr6Mo7Tquq
o3d70snuDuh571mGN+CJ4/g+PA+8wpcuBXiyX8Sqn6fa/MUw8N07/yWPeXAi8y8JZdsdhBOCLpzW
Mx+DEN2u8vlMo+S0MxHjt2qjQ50X9mR0Eyezf0gUNutu4vuY7d8eQq19nuzdg0ZvusIWDravLj3o
IkTT3vpFIi+vaMykZ1XHSYBgRgzurMi9geafsCQq1Yrhs1vLOSOcb5ABtyILLJCgkHzHBrxLYNf5
6bxx+O84NMwJJJaWjgnsJXl6Jb/mJBBv8Sx+fA7YGSJVwiZarNC1/myK8irFEsFEPSPtbQK5eiMx
9Bcj09cbfHnr9+szENqKCYPuvDKM+Xy+jK2et/0X3eknodYQOopkEHiLU88qzydmDRValFp+B2aF
C/jdfmYPCoBq8sWQGXQ3XuGP2Ouz4b6YXN3gR+U+vWRc0/w1RYKCQJ2SB7spgolgsm0OozjlPYHr
ytaxbSvceI2U6E3TdwWNMY9bUsLxQ9aOqROJ6gQyNaomsNz2bcD2oha9V2kuujD0WD9u5t+z2U3D
Z7WJDyoopGKMqg24hnj80lkdV2k9iuEBfXTAF76V9kwDEClakwfPXs3OaArDmUhqYuzlAY97EOnc
0PQjCWu6pDzqHinqBGRkH6GoZqoT3aKM5F/YpZY765HovuidiP1FUBqVwrm3fKeSNPgyUi4RfI8Q
rXSqPaXYScEd8hhC1zvoI6Y3jJnLdbS4KaToIFpR7eac4NEmAX7i16Zow3z0BGi/26bhkQmQEyLG
FtZ+AiyZXJu7DKaY1mO/AIIRWrdswJU7mgbJDtPHcjyMI5kXTF0q7ZQgblyJxLXW9U7izTN6HI4i
MRPPhVZR0RwbhVYaMnt8EGvYHpFjHoFh5jOuGfKxelVB4U2wLl7UHTxA9ZSPXmWog8lfkWwDBb0x
cZxNJaArpddWPysnl6yGpAkQnBwp9Y+UbiX7YkQ5MJN4xR4iyp5adTXf8AOC+cvdGDuEEak9tpsw
N4n/7gCI89hV+T7HFotLbdmq1PIA0wsl5KICI7ijsPB5w8pSM/UJSAZt2yXQPN2Mq0uz1zb0YCY8
HFi2WCrL1skf5LF5/1g4ppiHffOh0e0k+UecV0JDraIj1MnPnFNLs9zjqECwsMwz2r1cr7Dn294n
h1etSQTPgAx1JpeiZqSNbJKKL1s0KSDcLycZWAi9lfR6Utc1rtzRV2bO+eJjpwxbRscrk3kSbSwY
I83xkExv4yoyj+wmB+b5j8pE/8PzTGwY5BOag2rtDTEj+XHhByQ4iaHjDiXAj3HYsd0AnBMa5jo2
8CzmpDKGU/jidqAuuuB+HaSMrvwKpdHPFCzA9AKyAUOTB5KtwuU0DZR9Up5AOQ44sVDUUkFgdZMM
Cv36jgxY9WJnngsSBckqFa2x+SahBCrNSapAiBn7u0odQiths84p8NbSMPr00xh8243uW22X+Ba7
3aVfD9R5I8b+WPReeAzddTAHsvgNE/4pZ1RWFSFzJN4Bg3IQiJ4pZmsOb4Pjpfysqn/gDxPj0+H2
hwM4eO51KXV7v0cEC7BdNik58RLRTRCXO14r8s1GkpJTg+UhAuACAPC5oEme3CvcRaWqGNG3h8L7
T1DrgBY64cZq7qG82MUnebRZDgz3r3QPbq86bfFNr765GFhARoqcc24GbqB46UlAf+28LV0Jg+Kf
EwS8IE3EaRNFmNV6ghXD7MWUz/HkvaEBCkC2K2bVKrqeDybunS+xq76mJ+p9ZyiJi/+PaOc2uWcS
mV+R4Ndg6xu1p6Vylz5G3Ht7VsgHWPDdyxbrHKo3t4AGjwF/Am21oDON2uBIvQ7QFY3HJeRBk2OJ
oBHhZX8S9PUROjCuk2MSXnjzmm2gUzHvoCVq7GfcxCcdNURksJk1MQ2/s2qCrUN2vNS2y1C4eH5j
pTq2+FmqHIqW9Z4ltwDbn4Ga6kPLkrSKCiy6vRVny4frzppL+KcPypjR8QUFSK9LlF+hjeIgrt+r
KIR0JerqjuJO8FpeNUH+5vV3w13olVWrZ5aJ5nP5tydj+3VYfy50XDwVLGr5TT1SOkz6FwBzv7W8
IQiftK1PPzOeWafriGGW/xLZBT1qUhAbklNjnvmq/iB1ETMrReJABH0741jWhQ9hddF/wkeWZaQG
drALf9qXwA8B4MqTwEEjNAz71AMYmYg52m6kqrCXYKuMph/QfOf0qaPODJU3B5H6/u7zosXg34on
Wy0mXkL21I/1QWg4L9Gnf83iFrQj9WYk4YYeUj7YA/rjZYmdIeullHJ1BqYjLGJzaJ6iOD1BzIal
yRine107mQ7LrasYwurAmPkmfA493DmZZB3TXY2DOf9f6MyWvhiA7vrtdgRxpr31YtoyzD1xRHZk
MGv/+4g2jvDCkWwPB3rjyLCVymcBq9dVDj46xlM5amLXyCsXL30OupfLKsxVeRi46Z/0GRB7fOjj
/fGZnXubKStppVg1mBlDDMRB68TNwqBCNgGjfWhC4e+2EW6D191fGRp8YH1aacm4tOKqRfyXJ3F8
z7WdRpeEOB8Rcp6BZh8j0BXyczMtrItZK8zQWtEj8ZywsTOzRsB976I4OxR2QZwfWTPRP90Rftji
6DuXzzR1HV1jVbpfxCHrQMa0ue3G1eBT0fN26Jt2QQ+5VZSlii3JLUwCBb4Xc+DYZ7WSG0IjC6V+
OWDueXrFroTuTwxlNw/Jtsf6hkhHui7oHQ3a/idO+ScCD7Yhykt4nJkpcJa0raxoOTbemfI3tFkz
129UhS8tWADNRf45ePSLNZDw0C1ePsSSS74TT0N9WKLPwe7UyKEqRZZsrVTj12ppgqdzG7zIbw6b
v4UPn6yn45quHPHF0JgKxJ1UbbsMjUzNyOb1zqS2sb1QSCcaoD6HnTt8pvcrwZjie6fTKUzFZLFV
powZnRy6PbRaj/iQSDI12E0fS9TBdTlSqMfirpYThL6s31Jtx3Bvtr/KE/F5pYLmJZb2bXli0egT
1F5WPmxSLDiwIOqu3LpGlqbszlGYa3MeBdCJZK0soNFUAI/AK0tfY+2C03sXGSO6pWRAx6xkBnqT
9bFwCL9fb/HPERVl/pBWFZFWkH9gWzT728jRpJLkYfXAStIWk8TbdawRRYP4pd0XhFKf4i1J5l5Y
2Rxc11CDBa7Xn+s/G7iow1CsIR+cZxHjMztYiLedYhJtK0/ZJdS14oN2koDfTzBgE8VMrwtP5qWf
/8fZh4tdWeg0H2fwCJuQxUzegiystks2HzNnEw1aldHhwrWt3o7zff1KC6AmBT8MUYkPRaM/au4R
/xh/1bZLuNZyEFW/BDOGKKfj6wLw7/gJ9bp3NytZ2PEEpQftjR5g50C5O4npD3gWZwE3TixGZYSe
QYkWa4KV0nb4C7Sk0GAeHEEwjvLxQEhM6KbwWLwUogYH0qIAvrEELOw0S/HWRQFagUaWXshyQrhg
XzYl7uTfH1PpxJKKjAB3p3/4JtP2GCW/mKybaKtFYJdSXd3o+CCXCeIyyD30VTWaKQNCrKM0imV6
xvytyoCkiMEJcDrOt1i6B24NfNPOzHsbJQyd3XrpZBPZ2uieAJEC2lnB8Yo2KU1v1uNsYw1/fXnj
F/+x1EH4H/wTlq3gkjrYG3MKESSv+o4D4We33cp5XWBYxaLp8IFDEUrbaJknc/oUHBJ7sNH5iIVa
sHI2kphH2UvbLmtIGxnRXq/ccZGicieHUEH3yq1/GJq68lfIKoXz1VohOqsbWsO/3e+A7Yw9IV6p
jvuQlSOxYFRxhZk7WkWCg89Bd4azscNrWOMNZa3X6UVvq8oLs7+BiACZeyoM+/0PfsDx8D1cWmpi
xFB49v+VxnoQKY63gEbkaqI1h0gSjcPLgeu/kyc4TLjtTVyDv8OHZpiaTGUljD7emL+NPLRtu6E3
obUgkSrLCHyMDvlb3F+ClPlauDrIByYVrgbHNvEQ8nc98XEXr/fCM1ZZSfWbewW3v/OUr19T2HiQ
+Vr8zV6vZMyqs2bQFnGwW5+K/x5NQN6fNiGsmN+dQC12Yr8RKMSTq7hZcdY04pdFluI3QufJ01Ax
pZFbVVig46WUNwgayfG40Ow98LiuV7NPUSSqOJZH/5QlFujYvqAsw7FRxGXTV1cGJwQ8OQbyYRXD
KpN5ycawwAvICtAa5gSbxj18mk5Cj2c9pdONERosEZn4sB7ah9RmJHjAyMt2Q7FGufFYSNId7PDS
hRr65XJEyg4+fysLVqAS+MAL7cwvFvwjASckn3QOoqPvrfSBoow/C0V+FgOim+7KNAa9EpKRpYkj
yPYjnAh6t8pac1nWUO7Bk1iK4avDnPCJ8lb3nq/cNvhRE5wJoKmB0HRUNgMf7MRCFDhcjJB1ZOeW
Y7+ysaxXEFu2KZiGw4FPWHWcGnho6tzrIa8NEYAhterlYTZc+WZ1qSQNmvNrJPw+go342SuFefO0
wiYOBA7To3xyS/0koTJetgNUWB1dLmwGD9Lwp899HGcg+Jo262AcyGZqcOwA7xabKjNJVF5ezRrt
INLaK1TD1znIqAcuAU5KFe9dl31tQTfX4XHoYVkGkHSCLc/HuGUWcLr7/e956jHs9w0m0noMudTQ
g1kVCZYYDk0XndurqhJ5uud9F4D9RxyNHZRzuoZZJDS8N7T/6DEIsfvvG32vlNGvFu+pp4UX1m2c
7WoJlT1RICGlZcmWlbQOLT651QZTVTUVh6Xn4H3QH1F+l2nFMVp8OuLTLVK5FOm1MIwuIehrKulh
kIxFnlgnIgRdyBSUX/pduqOdoo/ktT8OMuwx/Li/3lSAxlt0vNbTPhaytEhg7MpolqsT4E3ABORw
J8IUfVEdsakHPet+z9MCbxwrIzH+dv75RR+3AJsJd82aG4ubvBVbW3iinozcm+kYKQuIv/yJ3cr2
nxJ+atPocwIxhy8jGs+JoSrj3jjf4p6fhY0J9sg/imk/WB0m862mEtSp9U2bT35gKT1TTlqggQTh
jNrTSh7G74d2oIoTxIE+HCIeePXFZOpxX0jmykC9ZOZk4vrf32/4fz88Y/5dHLMUdmXSKkWxGKdO
Brv+qHpBOLyjbZ2ojhTlFU0EO6V0er1045R9zynq1jNbEvW/8UwVtCVFRkJ9rSdH+B/FWulB0BFb
o4CavQUJT4Rd/Owk7MIVndrMrZ+8Cz6A8Y0wPSdW5jFn4nRhlqOdW627SRgwuo3SLLIjmnxQi9Bi
L//JnqtcVDFMSwhmXxjwjn3g+XSoLKGjXJl/FUR/bHe1Gcp4oHX5merUSr6fbFr9pYoOwuG7wUIV
Tamp2mC05/eRSVM6e5+mC+MQSBEGUMgihPQKg9uEQoWshHceGEHq6kr6hgstsHjmViXZ5tN+rMW+
NtWcalCKlExP15koUB+EbTrI2hBJhS5DZ3HgcRXfB8L9S0ByYU5LWHkaX4w4krh//19GeUfWkITp
6wopjZplqYKZVQG/eV+XhtkKJOSFmODoa8rEBGJ097cg++hCUP7BD0Di/m+si7zx9jn+JIrf6Gem
9Byv3In6iYyDsLhM8M7pnTLa01n3WnmYk3sYnzYPZ2ZJ540Wc2lFtm4BLtKOCF+0IH1fV/g/dkP+
iK4bh0+oDJ7zM0vaov6903U+I5V5iDvJPNL6+3yOkaScXbQqZGnpAlLWpBUn+XOysq5G9uX1qfs0
vvpYbtDy3yEIf48Ou6ZFX8WKNnUVHUEFhz0nZRTzw4866yBGB2fTJpOYr9r3GJkRJQh/IDpwtKrZ
IdSDSe9pgt3XfZ4pO4m1pIIAfzfixmemyTu+7GGt8iKV0wC+DToHgM5O1K5zTYduNoxclpmMJqyg
EcdG0Sfsg7TUjEXxafDSF4uoFNAjaOyQKbxfSvWFfg7mxe3/EWsa7OPoAjbCOpqYpkRppIaW4DQW
uGPIkeGr7Qy9ivy5t0nD8Cv96L5SAD8oOylicNeiRB98rnMbEvGFHwvVpJjcSzMV/EyN+Xbe4VIr
wby+pxUE1K4AVQWJgnI/98ffkif8ERxn8cCbcxJP2laD2Tn9VHnkvTXvWC1upkSBFxajWnXSTdB4
/iKXalugdDRvlZnf/TeaI5po47PiO+hN4yKyWwZ77kP/FGRiHn5k5SX4yVEXxu3P4VY+Y3PVxlzf
ED9s6eNm7hraYVF6CXLJypYb2TbGD2vao5soEseSqrLLDY9eGiJgzhfmfJ3qglTf3Qwxi9rnjMRH
MZ45MTKnQOGuvGiGYGg8Tdq93NDfdTbT7pJFxg/kO5Mj+npVZNck06HjdjIzsOxG6AVhDgNmwh5L
k8FTiAvPSafqCRgomEDfr6M1Te8dYJiwHfbFN7Hy8uEg/+W8lAsZY42LNKKYeFuBiovwKidWM47m
vWZ8weasXmrnsxocvvYEgRj6GLDTmGlO9qhOKnVJxFYL09gKA0sDIJI+I2Nov4D9FD31WFo7iGJM
iVNIf0SuZ5HP35b0ajnMMOu4P1BHFWlDuCou/VzTaLxBnxoO3cxvm9uEl4bDUNNyuhUDFTz4TF3w
gAAhwQmEA57HDnNr0uuss9U8C8Kh7RZ8jselX2hPCGxrptvxmb1tIw3gaV2lCt0LadTYAfOapzWg
H7UWlbVmXkiME43Irpz6nEgr2iuXHpvOu9IQcbQkzwFTcnsLtNjlXwFfrxqOU0QExTi6DMSW5XUb
szWcA1Kf3pDZRXXYjlNH2MoOyCZ4NcSTB77/Dl5t+HO4d+q04/wf11RX6KjKe7ks4EvfdbB8P8vX
11WSl4uSOTj8PtQ074siS/oD5+mgVWgVl8C10wxWOlwG4aqmUpAL7SzAtGgMi0rJhfYMu0+D+xme
86FHKQo21MkjDG+St5Hby27H2g6ZsRdSsO2z9SGYGrzNgy5OGMFx8n2ctJpVfELLmCsbzQyTZpS/
4W9ovmsJetejtHtutQoKNDk2PJxOnxt7hE/jDLzJNMwCLya41+GviT9xiif4k3BNe9Lbror/KFVM
a5myNo+c7Wb5gBaeMcGG6bEhnoZDdypeoDVBDOl53Rlc9rHTll8Y8pgBcuRr2YhfUIskfmIbM+MX
pyRsdor1KJzBG37HOFKmzc+GxxgM4NGj6SEjjy6zhw+mi663IBvVco2djet/ahhXAaJFjymOI+gD
OMB1RnLIpwGPTobTdt6nak+I8Ckj0thNcWTTpQbS2pKlhU8JLiEC0mODU3158Pv4HdhrImnLYcU/
4cdLonq3IaMlfkgNkh++BzgT2xLmFsUKj11ksinUQ7YwaNRzKAZ5S78XqE1BqCGSuzh/w8vlWsUZ
KzjXdTgDtLnY7cCIl5P6BIcghLapz5c6275cvoXWRcUgMBsSqJdRlt0YXA2LZp7LKR4SdeSL6i5m
eU2/y4cFPmzVRkO4sM9bC5pw7dlmYIWZ41ly4KdrcCW74gcOcNwhLi0U5i33IjquS+5vpoml3hRF
kWbpQZQ8QqKZ16Drg9aizzVCnFuLm5XHXApT85FIvwZ6d7OiKwkHcIDwbDDGqR8cefpRiIc3//u1
HbIl67k3zhZuKRv0t2Db9vmrkyzU6zNB4Col08IS6jSV0UfWcBFG7s/q50d1LXT03b34Bzxy067e
pGeQ4GuKd+/Z+09UxxVJO1FAalR/8AD7RMMihR4F+dKDkR0U6Hy9xYPCV6X5O5zxndLzalh1yASO
ngtMcy98maMM3FeYDbvMu8R4WSr5eDVYVkPEgBkaWQAlE1F2CGmWXecw2fAFPQBkT64bqhyYTmKw
YXjqNl+4nzDSJ1M268zPEs7nTRYaAirTiywLq/p6W0cmSJiq7rxmbkNHssAEztC1yMphy8hHPaQV
E1Gkcqu9h7UlwA+Qf19KVaUzdIZaolVotzEm4RGKGkYCco7Ym3RQFnMb6Cy867MoWN/NnwV+/AbD
d43Z0/ZNWVZfP7K7pmpqw5nvPN1pPgPsc/qVOk6YDNDj04YS+YbtvjoMw3R//AFAIxF2kAqZNvaP
LVE5MMVNFYOewRpuXrzZgnftEoy8aupFfwAAb4y+5jFjE5EP2R5ZIRjt9lCIZqingikRD9d7BRNA
0YdwvFlXufgVZSMBa/PO6MBMsf9+PNCJFDjxXANBs1JZdw+i14RHsdyy1+psTjf1X8WJyd1kNonk
WNU1s2dCEWbraadMaiUZeuujXDlDgUx4i2Xx19UDUzgEaSt0d4OyVLoD0GYf+xo9ZOGZRQpfUfus
rWTVwb8AwokH5EYaTRmK/D7NS5I+khPG7BNMDSEL5NFx2ZcwAP5ObRVNz3C7iB1oun7u5srHfIYc
Frzzb3LYEipHfcLgTK+m1ZBuD9/IpNibc/92o3o/yy/c4syN1ZJv7lGiyolBIbZGqESb3p6+AK5n
Oa3Yg4fW9THD9qPa8eE1Jx+omTC9M3TrIUGt4D+3Oy6suyC+uCpuQ9fUZ+++Uj0XKi5JPThbwmYa
AG4feBwAreJVNcmHm03DmMEqQg1wRKKJOdDi5T7t7yElolI0hNUR8P4nwSdybX32Av1vKD/6NBIY
0tuWY0Zwyv3opKGrGlcwVC04Y59DdGHddTaIGECSddvUwjAomqA765SNVEhECZyR/GOw0i8P5vt8
TlGjN7kc72GAxEN2jljWRAk3FhGgMH2pegIqJKmDFC4KbMphsHIFMzKqXcoEBrzSxqeUIz6Cg60m
26BqlLmCyAswvj5P7B9JLtI38lI3+uH9kBNHs6YDMtU7jkr3w6DWFUvkIIXG/k+VcCukVgKKPfsM
8j1MfQnWmSFJdZ/uF8rK2mVY2pPVIv6bjc8MIJJ6Avy/xr8f++TLNEa/MchBi7oKpcgCoVmAu4mJ
q5sDDnZfp98TOvuauCEGIJ+2t1r3wcPGewYpsuDk6DzCQ2QrRUBA4YcyviQpaU64zhzRb230ObXf
O1EbboobiWB3GASAtuRCBLogDYTSAnSzUJNBNQv8hOT/KMew3vpAeZFZrIc/XWWnu/KduicAF4o+
/PiZ5BRuXxLyqb3HW8/ACTgLNpwl0naZuqE6cpJ3rdx7EkXyALG0aSnDL6wbVWn4HwCogH1V03p7
UzehK7vcRVkrJcM6/i40yJlx9eBOoXMA5wkk3tbnQiZL+LUhTgCu4RznaxAGBFZWms5oOYfY+etA
sfOe436mXeDMlExcT9vi/rsPGGcZg8W8mr4d2C+S0TvBGt1bJDYrV1+2g4xayCTIIg3/YgNfv7K4
i72phuI2MfWXmDWC8wOcbh3qJmQzwj9ttks5oIoDB/SoK7TK7ep90anJ7t6GV1UToLK+S7eNNCcx
W0QX0Gbm70vjB5yEugo+WGTDZEFiy447j6bYnL+5jhMg6dinHxuEi8xXByhtvdliW9fPK+cNIeFU
BdGPXuBKo0xJzyJLuEDfMG8TpbKIXMTJwndm02tN1C09wM5kUJXEePihlkx/ZjFhHLYdV85jknRA
HgXjrS68yMt23kCjbC83glughjXPR327zALlc/lhKy+/9qUJo8C4qSINibYYv0EPreSLLLWTHA6T
cP1WmT5kHbSOS5FxCcJV19tBIbKsgQGqB0den+w8Cf6Bg13OUyE8EP7dG7ziulMRiuaVkMnlNwfr
e0v7NeLdNO9X7QbzD/fT4fRhWEG+biwuaK6RVeuqrZKUT267ZHkJbK2pjfEO9W/2VZDMn8tWllwc
ynDkfp18jVzVMOlUde0iSZkuRlamHYTHQR9Vgd1Cb7vK5TnD3kVGGFdw+RdDx+LgNIV4peSZ3NN0
rhgc9mqScG4b/TTwsIIsCpmRmkL1vLglj+iAcyICHHl49uvsf5cH8egtm1ykMhB9gmVBRjQIf7DG
mpoaM2YZD1UgDMaA/ySZ6dPWmLkcWeHDWmXZuHT2VDlZRei/yb/GlmEZZkELca7M29tyV1/WaZek
rJFuPC2p9dPpUkcF9Ii5YonH0O0w0/PgzNpCG9IzFnStzCtVa/uv+GmFMeUQYOsgcoRlGV4tF6Ga
Y05fH67wD1acjVPdssBTY7wHi2Mqt4ojsAJo1aeSJRUksEpbUAQGKlTv8CEnbOViJo7qKUKKp/uo
/rMr9U6CpMPzbmprmHz8N/Uf2wFh1QpNuQsnYNRfDAr+04goxNx5p9CUAySIdTUa/bC6ypmRpwai
oBrk5Qrs9/DdI0Whgosth0KiT0XmL789xB2D+UKnGS5Lna7Gpn2HRJs66KvwSfBcWKMPgEDSZRyp
CyAOWbgMpUxrne99EFEZGUBWXsso4hdGY+NcX1kiU4+1pYpk98Ys0MZxnmXx0w0DjrJ0Ihvb8qUC
dFJ5ncoejA/4ScWA7VNLTMyrE0995fdwKEKzkzLRsTmygWosCgMrD/MsxGoYiwk5dgLH7ixlwQRR
aeRIK5v4X/ajzEG0pH1jKtMxwTBrIqQx/7O8il00akWtsVkZhkxBZ4PZ8qk+Ium9Cn5cXpXl4wbj
Hc5G701SSbjMhGEZBdk4yFlbMXhySN72VYdZWZ68ISYzrIWaUjcCgDwUPLqn81ftrFSW05mm5W8E
MUkrFZY+fewa0jPog1aMxNT62LHrLOfT3kMHbxbbnFy/yZeNIdJsCBHecBkw5Acilv5YfHX3pA08
UjwZcBVMkWQaBSrSv4ASmsUDnXyUsoxwWwtC1sUT953oZW65gZWsyb2E/eZJ2xzRI6fT5aCeXJmK
f7SJ+oL1zMi3Q78lxUdvD+MDdAtC+4aTk9coZ6lwouDSSSpXm7BxN/FJqRwKXFRlEWSjd0heIh5B
NlJ1Mq8NcMlgz6m8c7OhNlIKMO51hFOEHVVy2JXmxZYnmoATucaR9thg0XX/iGs1kVw45d3QZ1Yz
h6orTzNhHq6chf8cHSt//AITcrNg3W2G1B4CbM87Ozgva/zTmZjJJSbECKQ8Pm2cAAiQZPsoooO1
jCFfPQMSnZWvKfFzTpkSYlCURRAVDyfqiN/ybEELRwiiZvEabUpxoPeDMzCL8K+XDQteWT4fPYHz
XRX/3vZOsYm3wR2OE/FLYprspayuoboX2hRiG1WHtnUhaI6VZxepoB9oTUSDo+4vX0KotDBNA/ef
bX5taWJ5l+59JgDLaczIFjTvIoyqsHzaQb94wlzy1P9g5NsqZlTXp64A2wIwhrue/XncSn/nd3Pk
amoPUD2AjRnRTUjArO3UKgu9i21sg85eb4vrLOI1n7r3AOEqtwwf1rI0xn7lgrhs+LVhkgW8IPuE
/3DW3TuwWPBHaLhqYVmWBhEwVTZbD7A1O5AJupmA5jGOVUd5bw/cE0CLzlpXbRenBctL6xnx+uGp
tu9HUCma+Hf4AkXvMqWkSk6X5IVUdMymcaAnKhtcJOnqE08P0BxELUYeGb0qXw1cXBjtH298fsyl
69a/V+nYt4/Mlf5URc8HEmTV+hs8EaaJaVCqTlF8bzvw6aR1epA9JGc1XTqts4qKxBYhENzoKEy9
fFewHLZ7uSeVMmgL/RG0ym4fb4/v+F71E2iC3iP5G9RqDr3zfX4iX9t/OKeGmYyAR7GMgZWvYH6R
s/nWKiolQBYyhxziKfvPAgI1lCBS3ac2upPEU+4KWLxeYX2tRojLS41wyDKic3cntCncMGW8xKTT
fOhQGExmsX1s24ts8uQRNV0EsZRMtANZitCeCSHskHrbvsaPQ7uPaDSY0zV15BM9gba6SfhHgwd0
6Ac92isVntToqerizv2yTJLHLmQ/4PKe6W0PeP27rzEupJuiCFZT8WTAyZOIqRWSBREPOMCV0A1X
IlKWeVJGHq6BTDnU8ldSM2lqPP5hHDsNjwblO3S99FJbHD9BESzZx8D1OOc0MnwggxGYCsUZvm9G
mZhjOi2EYvV4nqIek7PHVUwLkvxvnA+k9y1NtgsFWdLqqu4dSHHDVoCBiVDtl36wx6WEVKV4Zxxj
rJkdlmePwlhZhxpJS104H6mvft94HxpWDUhVmh4+mZ4rV9nVJP2NjqL1onma0Yv1KerwTUIIG+nh
kvx6mgNZgaMnQaHXzbaBaIIqAnSlV38bgeP5KhJ7FktjlIykFj55M6Eh5012Mpu2KKVFxTxo3Y+Q
qtBQlswtmc16WbGQn8iLl9xN5nEZvIst5fwKf2N0hVaepkbhiiCOU+wgqY9fmA9Fqj/eocijfNPC
XoaEEQNE8aj/qlIgwmeN8fnBPWsRY2S+JjwR54n4F5DW/qKZZIj6yOXn/YueYggKpnDYJGIAr6GF
cmXgxvo+S4vY10XuAjCPD3qzm4Lv04p1ZcvR901uZ+Fa1002Z8Jbj9Cftr6XosR1tTPOVAiMKrHj
k+XDHac93ddLqDvSf1wzZ3wqNqBxryBWemUm0w5G9VMsA/471Yp54PUObjFEw7+giWlZByTkLPxx
cvYrOHRBF9Svojy+LMQG3dKIR7r/q9sk8jf3btTCQCthw4jOyRp/FEuFt9eQZik5iJzwXHmxo6TD
wD11B/f9uGEdjfvQK3AW1GZwy1nB8G5ZJLbh1OT7oDTbY9tak/PtZ41RjaXh1ZpL0vMLx5iA0LoG
k4kYNJTDip3FGNqTkJzkz+OuMqs4GIIpo8Y76YLQVZjEClZ0zdbiuXXw/uL2Ns7/1kxrlcxf//yE
tkB9ISAWzPNHD3TbXaHk4tBMm56PM2SjA3Ux5XmZvBN9GWMeiit6ssQ21kjJrk/l5ApGSeV/+6a8
kgUVyEdFAiJiYbKJdiIhTq5b7vVyGTmOQOQ+wVIR60HeThA1uONHLM0x1eRGyU4XtACK8QQGviHD
Zy4NXBD4zhzxMUzNkO8JtjwzdxwZ2C3aXWIFm0zHmLgO0JmMFvl3i17X8xJs3h7s5740uGbwKM+W
itQ/3q1PBlS86l5A2dan2lLJxkpt4ckH5U1p75v5qaPzGdg3TqM+bLEY4a1iBWui9jppIDOIkFyw
l1UPVWkVe7WWXKE6diV3jVFOBjrDmH7z7BGJn456XH4dZORCwaaFwh2JAHQ7jMpZbIzmBxjx1WXt
CwQTcV2iJBL34tlCGUgjmSxcSNN5bHjo4BVN9K6SaQenLu8T8b+cm8dCXiUPFxK1W+4+s3rii+mB
YSy4bfUP4jwUa0OiVUhb7+CNsc6gkwefGUgmu8ouTn7zCeqLTuf6/wNcweh5KfOk8nMaCnHxNrob
UrSiE+sWZPB0X9WBniaFXOAWxKM3VMH6+kBvs6nHpzw+i7R2Nx2x2rIlntnDcPf6soeC7pwQ93KX
Lwt4z76LAQWnVAP4EY3CdB+ZB9Y0yzc2/Cj4gpUx9rU9YGFjGg9P6oeehgTIQ3LTpjW6KC2qnKuC
24+aimKi3VyZ7qEjxM/uXMeO4jwAF9kbTbFbjxSzmUnT4jmBeZb9+zvl4MWXW2yb0XAAp7zphfAq
RTtNkIriTX67yso8f8LqKSxZFXEBuY3iL8C2/PhWAoTvrrx4VihzgeoWcx50F3sSb5cNmBTf0c3H
xprvMDJhGxW97sWn/c+B+ZfLeLB+absPxaQbJUy8X7RoDVGuS/NmUG+ZlKShSoO5hnGc1qX9CE3j
j1UI8S+nbfjPIAdyKNlKY2vi5+s7iooM9FhluDDY/U0cxVaDGqKlm9+iag4Rh97fAUnUSom/BXdG
PxKPYYeSCkE6S5ey0yJkfGirtBjtwqpQjB6JCCAyGUpifL8aqiu/M3p3bSlDtWYCjQFylhvs6nh0
rbKR+OTcpFMxumfb8t8y0M0o3zH1s+QgfVw7WnqhSq6X+ZZ0fHbz34/jaItLENWDGbp7wzBT00Y/
/b5FY1IJwNnTLcxHxLyuQK4LOtvAOtTLOD44A/W5CMqOdFvgqkZgLzZusv/WG7xM1s2Bqa3avDnw
bYFgwWwfvjsh/sk6cV8EPjf4Ptw+bsw+PfaRVQG7IFHFbWJG7VODHfJRNf/7y1OAxnGU/IbzlCMk
ZTytmjDpT1RXAXZAqhOyRjJLwXQQtFJa9cCJnln9eiom4SA7tRniLfnByoP4StNPgoMOxEroVtaJ
/crEfp3641ZQdr9rGOn7+ntpKoSdBGswWjEdd/A9oC4icDca9YhHt+y7xnidlVFdWHXw+S7iGzdb
RQdFrnSvx9rJBUnfHG12ciPgHmdK3fAeGMTWm7oo+MQPb08uVSX1PyWtLgeGPoOEvSiXtrlWx5g/
k43zuJIJ2JEpHjhzhCGB/OtOq6L6ndi8VbkSz/RypiUX/2PMfXhHj0/fmIpo51t6t/K2I2H30ZKv
NHvfIy2KyW9DgZeLDfjY2N5XwpAFvToq5KLez66ihVOiCM1A4bp1Z9ffDTBSNyirCixCXwiivQwB
kebruLjITQIzDleIYfb0FkCK8pVEWfDuoVtBW3V6a6ZHO1dI1R7d5KoMXcaZwXvc85aIV/+wlv7r
D2cfLXz5pwqG2KV+tYQ8dYde4/BO6SZ2CP3VwMSyxd98Ww+1rd+zRRqEFiT1YkqjXBvDkRZ/6d6d
yarcgzdZtYj+aulFoobmh3leFgBGPzVvle1I1NJ9oyUOWpULZv8Hq9EuQki/9uPWVNw3Dzv0hBFX
I64jeUQ8uzxUWR2VPDObsrh9ToEj/L0uFyqqV86zihHTRABWawsiPdWii0cXn2FQdd7Q92X/Zp20
GTZIWvfgFOZ98sGJFHjGq9erwvI8ejim+FRNYwynqRpSZEu4KOYhNrlJ3uO3Ntnf2xqZc4luVezD
dipYLP+GDW5VH16pj8ZNLo79Bih+1BNFPCuW2tv7eRXmQrIKdCNo8cZU+ExubkAQVZm24sAaZ5zW
V6j1BuAz5LLFtgz9EcUMQh8q5cJoViVGGTPu2tIlsyuF2sH3Esssg7R5iRjKtnLpO7jXvd3/SHsI
sOUVH7PEN436TV0cGBUmlYWbKf0HwrRtqNmr2f8MbwAKdEKEoCZPtG+kIYxoplPnWpWMY2t+1MSQ
ko7YLVJEyJJsVUy4KC8QNfBrLVGmXUsCsoS4P19rY2MSIC4ktLMJEsVegzb3jNe0Re1DEAja8Fl1
gZOaBwGwPVIJakrpXV3EQRAXKDmtLL8C8L7s2BmSuRiEJXYJOOTEB9p6LKLUVIxO+Fg8wC5TvAGL
CuDBRtVjPUCMXJhXCLnNZ8TWO1GiiR+iZk4zzo8CLq+8EwLNFagxdpxeeehMDLoJMCdDdSw0B6+3
iKbjqofWtPkIafTKOnwYY12DZBLdBWABH9Tll1YHKX65YlBUycnkt+cIBbKRuAYLT5fcFLBu6L3T
4TrMu6GTrR5fAUKWznHy4C4611uVilChA2swS4ABvCvbcadizjwNlMjDEwI84Hlk7RGEJYt7RCUC
Ei3KuEWsEKXokP4RExn33y1Dmm2h8PDZVhWcy7iF/yOwhMwADC8zi3hnZjD2hfIU4lUWBAWX+pqf
d72Pp3WcEz4H8ZPiGvVCWo7uYUYiYyNG7fFDeoe489soGhTzorOR0CQIsoUyjAnX4VZlep821JsA
OkBhgO25/NkbDK9G0+Ai8nScB52fQlpiTj5qskz4PplGkL8E+s2aL9QEPUxMjkpfLkfvfIOQQQ59
a2YlzjeStuXidhtKByw30H61RY/DA17cIdiTzAg+iRoR/t7pKhnvjbq3N9t+8emGjPwvbDMVGXI+
tQno8pQXw4bIUpEQaKXfQiGflHVhc9Dsyy/vWw4lk38BHTy4aHMTmIYEPvHlNPLLrfDTAYmhg0lG
+shphOE9Q1qErjyLNydp9a79OzUsYb4pcBQcK4m73Z7oe9nB/w/AIqd/p2RvDRNThOxCulPt1pPz
HkSnDL/mnNagQ1eablAIo/FC8NwJNuL3VskWd6Be6hX9lELRidFMJeg8cVBRgw/QNJg/A42IcVn5
e1Cg3DBp0/sQQzwmV+i1K6GwihV/6OXTw5EASrY6NelACK+2PJznv84OiGDemUlU3pUuS8DM79Yr
w1zIx/MFBRvy9JLyV0D/1JCfEha3KKfdKHLdbaTFn1gi5TcHIa5Mnr4SC0hqOKorQSUUH4sOtvmd
JJ4EDzeWCkSEFtmp979V1pe3FkqeUCYFAu+HUyyWgQnjpFMxcsx5lAJtnp4qFKtD5pLz+qPPC1j+
3Z+DfMkxMA+/D7pdzpm+qkr14rXisM/D+kp23OutG7e77M7QYIaZNskD3sTWG+V/EHjRF4TWTgcc
ifogIuX6KzrizQmQzWv1mr6BGI2aBYcDwlkxZb6d7yk/BKhIOZGdLYyRCCLGE2iSH9+Z03Vr7std
hKbir0s/cGktvR3YWIGa/KIPXOZ7yZbOSfpACmNfTKoLYC9lqHaxycUZol4E4u6AV8cJ9ff8B6CE
fWusUipllKnLP6JjYblABNFVn+YBNYHH1mf9udowmQWpwFdZC+m2l+GCGhHk4mc1PP6FSEoeVe5g
gus6ajUT7hMoOMy0VkEL2pA1JWJMk82dAIp9iXfqQ6IhQgk06E1bLcOoJaC2Oa0s5AbrZEoPmBpA
gls7zWsOfjTXdifUnC9oPwHZ52HFYO+E6wF6T5n06t+kzw16qp363EOoOFaZouZ+q6ttJyfSk0en
wMoQfVDX1srDa1vdHo9QJ6sdngep0rGuDi9O4725/zzstG3Ln7OkWqTnVEhZcP7v4ekNQn3bXbJs
MrjFAwB2w07H2i6Nd/R89bBh1hHvwrBj+QO0Dyw7BVDFWp1nuwgofsJl+JMchSQwf+4ZoqPZ2KpL
XlFFahUQ+KgDD9e/aOSef0Ze/SAvIQZ7Nb5qwLQ96Hms4lc2+cTqKj9UWei2Sw1qHGuY/BuVxIN1
NkerGkqJc6ya8JT//DIIfCPesRdMSKJdV02UetQH4PT+leRP8OP9UdzHMYXAs7o3IvxmkYN5EZP7
0i55c4Vb1wjG+YUN9ULSlDiLpyjrDXQA/4OY7QvA2ATrbM72Fj7eclotOHg0ICemXuFnCQ59lF7l
JVlb3xYPsSGfgjFauutIYAwX43ZZ3GNLM4QRyopCiizhhGoz9EnKlJ85DFsZtYHBlc2mW8dRYcjI
pdUtEu6QL8cFJJ6RpEvPrUlfkrlsvigpHHIpAVJKSdqXWKyK6oeRhFcEMh4fx1R6c0ndzio/02jy
2/lruHRbHoU/XaywxJ2QP1vQTUjV0HFHwBm1w8DSPvZN+yW0cztfBehPai/3MB7jOrKLgSCvHAyV
vsYKxHQCchFWq22VK+RDqw1ZJvubCBmCFY3lU8WtSgnjkk5mtBa4hwXErTYxtru7gGuqQFbixNQR
hKkJjkSAkWlYq/tpETasav2v7g1crh/jQXh0+b+ncXT8RZjvMpSRHDDzyHIUlJHmgqzlko4bvuUk
60SR9iDtMH0d39TszTNi5obATm+NsCZTu31R2CLL9jmGSYJKzrAZmifLDyRGceWogFR3Azna0jmD
EoyKKpGHmoyuIowPcu+EJzYrVvjRYqGX322PsGgjvG5O6y3wK9QChAyvulSMGxOxVpaO5G3Bzo6W
afLnG8FlC9voxj7f66g5O7AUqJr8o8z0GchY45IvCVbv0bG86z1Z2fynO0kE76kanT+e7Vg71qgT
y6kcKkbIV9/kGO05b7tZ7Hd/nwhARGvefJ5fHqE9WdvENTz6JzAdVM18+d83eXFxnOFRBFtqkfg2
AOiEehMSSI+gsXElJi/4eO3ceup1gPoQBQzwSugQ29mBI1DRgwgss79zG7emY24zOsw6vt2LUqld
sbZIP4dRT8Gow1nqnAatbMH2ECcbKV8fJ3Oew8OF3y/L91xtGrs8G4B+mAHzbaFtEP3WF9Bhlx2U
RCHfHgFpBVHZh6fFfcHMLDO7cC03w9Xczz6NBmJueIB3qxfOs/BNXUzG8bBPtYsDzfp7y3BP4PE7
0CQIaelXFsHVF68upW4/EvugUjcvxvxlSjibtX/7QQh22lxAnK8gTY8ZQx3oRl+jCaek/j8ynVv0
+c4yaJjPXCcszPCrIRZGwrqNMBd9U314UvhCB+917lZO8GOrCUgCbcFK/zpd4o8StGcc+c6pAaxW
8dmUPfjVpEGXGM1F7e4ndd44C33mjqgG1/YyENBsu/w9ZCOhTSSBJm4f91QnaTwLN3fBBGu53WSr
O+RaQQm0nvfDU87j/N6FyqZXYWkGxw7bhm6HNYVBFk7ezanQ7CtBx58xP+uL9VGdGMgR2zVtorSc
vsEF3TtTNwqGnVrb5mGzjw9yZGIQ5xx2JF0WKrGfy5gcajHBZqIQ3s5Qx0uXlSz0Egs8+wstm+B4
gyD0zN1v5UzVDieucxYWFIk3AMRdp9F4iUJLLVFqo21BmGG1Oz/k0dHX3UGfwGnYYAnVZdtZYHqn
apDPZ5+LvPKMV6fcRLvjzkkUkAdhetCnmYOKCeDHHh9XZG/185Rzjc7v+HIV+Lcir1Q+OCs2Isez
Lf7wy3NGAFAl2AmM3wc8IZTXkLVtoyiJ3pxR79a9rlkPwk1PXtPlVmM7RmOqElArbUl9BqVUAKd0
II1zKQabnuQJEfbNSNy9jJlw6Ui7tAtKs7Qr5hh1moXIosQ9hhsn5QWqoY4vivOERigM73CBe2NU
5/k5+TdXdmcATEReeS6/QG3yX1rVxzRweEYKSJwN5+EaDw2JY8LzwBiojF/H/tSuqbJPBY2n6zWr
CINVqLR39wyC+SsLpaztknW0gVcxtpciBRDBWOtDnd7oR4xFZ9pTNbcq48vs+7Tw1fcckRcm61dl
JF91LjuAbdvvh7Ss0mpF6aHmEAUYrYCaEDOUPdKw8YhldUgAEoLDyVFJi3PAGrNJS9UTFql+yMX1
sz2FHPLsdQvRlh/UJLD9h3ehsRU+wNHcSwsesxkxDNmgw4ATk82PKfHpurunpXDCSWOpU/2Q9MTX
mLtkvwBq2aAWhx6V06OGVxrfRl400B/38eetpDHkjrukQ7LRwSWGPuR69lOGrnQslIfr10oszwMg
dPxei+AWoUL8F3D0PVyaEf2VC3OihNDNGE0WgOpesWVZhbkU10NfS/Yjf/BVY75Udu/ywvGPiX59
KJikM/IiPX1UjSUVj/yQkXFmlZBcEkK2/XrvwNMLGg57zrZAUOhuJ0ePlnB7AHpw2aXvVTUx1Gzj
AgMrVBT9hVqPwG4anSjHfQH16sZPqkufRRtazeg25ZIis0kXSBypKhrMzYehOaSqTSGqVfffvHEC
8jKXlMl5d7PNZVvajhKKjzjRis9DOppmcsoH0hc52C447aRtDSBb4fXQ4Od0uxpWGbtOnxQCJD28
HjnAzHhDovaZGWBK1pbLT9FYOWgTWvCAqdBzq3IbLEKg9FodPhSaVurcurXn85kxT+SxFLfVxQlP
aiPwAjfRrgbI+X/kwLuERT0jWuQ78e6RRWat5ZpV98T30FlD+JpgBptB2NZbJXz5T5Jl1dLOpwsW
wk2ldwHP34QkkITuFLKJrD+PMYuUKKhYjOMDXZ9R0pa7EkBX+Q7WxWSw3IsbPwBEQLeXBCYyHpKe
d+o1ghZG8n9rQgUpMeDxj6r8vyJnbb4/1+Q70jfTRUwl+7QwUzkQ5JG+954AS9W7xNFVNmNl8aGy
Rj+8iudqPX2X1AN+ZniLnvHnS6/9FLLqODLMKQDMiSA1PORu3IS9uf3y12OU6Hp6XmbzcKjcvO+h
j+R5QqxokQWUpbbnxsruKOzUpz2eVhuvNj5KbGc+60VepgonAalRGaIoDtwF8Ysfk3HVIRsM/Sa0
zXMbDFoiqX+Qx3ibNtCn2xRJ/KNqdHk1UlkyKYrFwCrBOeojuCwpKt099OqHkiV2Il8ZREscBbUG
d1roU8xpiCGl7aXqy4YB/QhmJsK5pZjknjQi63qMmLHz9JZXnWtDH6Ai1ViF5E0Uc2ZzF7N73ZVF
r8KzwFkxgbHNPRJrwoWnkSom0UFITlKwMfq18MHhw46KYrhYkcJvOK0CeQgHfa+6xZrQOvu13Vl1
rE2r5ko6XqpcRu1qvorBVgsagLuhp5MPEbXi8UZ5ehLWWUPo5KBaJoEIaj0PkhVdNlmX9WujA8rm
kI2hilZvO1R/9zM3LG/c2+epFkuvrf7WRa52IhO/PrBG/rkOr8lZ0jJpHmCS7US0N4ZC2QbsOazz
vlwFWNCT+3Wji5tFcrrPNcVXyvTuBbclCkoix8lRWi/Hf9r1rbM7CgQ7SDp2xvOuwrVHAFx/eSsd
spH8FLdj/PM58ITyfqDz/mSvse7T55CB0+0oNjE4iQ/53YYQwsSZZFwjpbTXiYY0gjbKbaW3pRT0
rzJxi+kltAcivwbfkKj17L5ODUblFuVQZt14dkIuA2qT6UiDeUb0RI7s0sqR77ofjqdj8J1ZmG2i
RI65ZRLwGw+tJjln0ZqHrNnyDhAzMaAcxJWnehAiZfclP1uWgnr322g5NV4Nqt21j62fwavIZlNU
hOIs/H6Jmh+ndNBtkBBhp1M1ZND9WiD6FK4J3l9ad8M2RnQpF0IvO8JRrQGSfiLSfAD+cWVUHmfy
sYbZo4ZRlMS+8jxv7oIMHny/DY0JOUsdaTGUaWpOdQ6C1qpMuMaGR+5jIQflSPnieYT1XxLghaU2
5yZeTkhwFm8IX71F9iips/lzhkF0u5mVYjwpjqB25Fk0enHW33j5laX1qa/TnpOavmQ9YEVr2W2h
A5I1sFk9nn0k/voAZ0wqqfSyz4hKs0uxbqUc/s0c+3Y7Tn9NMCikWM5bbD7wdrHaTIXuhR6jR8XE
xIgpiSoOci4epMxNaUyFnDrX3UQ11eIEMp6eab+UJIU0xWg1hi1WLNmy20tBE/9Lc38hSNnX6FYZ
jeu4fDcVperb+C7ajlpmHg1Necyvoilmu02sdFtnac39BKmpSg24t8ZdPrN7cyZzFDC+iWfCot5g
bm/EqtG0WGJrGYG8y1J9s/eEd+nRepNHe4V9WxWqckFv83Bc+ltUheEqHzW4JRL8RpzbDgX1zIEQ
7zz+kxgKsMpWk6qr/i8xdWyJOz1o3ScZo35sU0E5j0DmAd/aOmJC47RUPJAckcO6X+n9fm5tYRyM
8TcBTc/P8vMtGL6SvTMZQSb0bE4fBbzZlJdWfPcHFRpw30G1vsyhdGS2SD634RuPlkHNCr2Gu4K4
6yqiLGmyqq9tl3l5xwr642B/PToxF00iSValHp4pFZoG6E3eVL1nGlY+JQh3e7Ual55cLD5VEdVB
BoBu2QQdKYnBzRhOIYqSHXCiWrdGxItATukCvYigpKc22tYw/eZ+EoUmgYmxpbYnyx5FsjuF77Ic
jSherJq0oHA3L6rnQreSCjiM54G0bXZwoxCgr6mpZw2PkA4I8xPpZwCSJ50uaNq0HB3uXhL+7m+k
1nozSdgtknObUp40avxSu83xS9JxF5CRho+smfOdzM8bRiG5SZWqPxGJsYgzR5GC0vxbzfhE5wAp
w/HbIlGWCjrZ4IQK6C0bv33876G+kaKy+LiXi+qWFgUSEts6MvIoaD+3ib/FiPk9Z0CIG+nqIU9M
ejObsuLmzH1FdOiFo67TjCMVOaJIgLUzbmta+mtAm2D+wUhwWxuijRdaVMiJ5EZ9D2cmzPqKpF+p
YuIKG/NcItfSCFyJ3LHmO4qh+gOU9hkqcgwXtfOOHcvuYJMjGtv8MYri608puB6A20SGOvjIc2Dy
ugSdhqAeIFqZ6a3xeklkbxI3HV09rEtjlAvWqxX0/FvBvUXGCqJDa0VCs6NnOtkWREQ2vw5vmvH8
h9kDoUVbigK+BuRuC7UsPetLsovd8jizbI0A14Xty/jiVxpZgGla9QW2xBBJ+RJT49ef+VaaZASF
KEbYYCtREi3TKLRxHYgGnDQM9jgagwSNqUVC7JPOMK0SCJrEjpYgXGmxEjB4Cl15p0dglpsJY4zl
TW7kwZ47lkjnJ36LPbcVBjw6PBUN8n2ZynSH4GS6bBbMSOrkuSBrC46KI2z+sh3wfilnCHRqC65m
KYKnaX9N2rCJGBsP2KiPOv/Aofrc3lZoP0uvSsGrJZs+t7DG7orvcjslX4+j7ppIgMiPrKTFr0Es
H3uOOKxzzZXGmwpsJDMv8s5uYA8gJH52tqZ9x/ZPz26GKPRUFAZwq9ILs/D7xT95KnLppMgFYC+T
aK7lRsIop7dOLlM1kDTUudrI2RDezDhS3+riWLsnR/gvj8cdAaiiUEot0tdNfOHa3mKey19UJoS4
J+Hwm8jOAVTlzv54BVigg2wb+xZHQpPBfLYWOT7Hqrb0Prwc07CPpGZnO8znJGUNi0QY6SzEmr58
bPpgXv+iogtAwB0itdhdTgroIrYQKWdNSXjC6yaPBUvDpOwOZlp8IdsuQI0WHlEK+3jJ5QnfYxkB
sqxB9RVsRFuTHkbBM28NE3hLq8g3kJySHUOMwrtrGmSNeevjb0p4X33jfJ19/72JmEtWhmW55Tfo
NPG5s4uTVO8li8uQp88N34P4tHPa8ypeQgFZKn9mlRog5poDOrTNxY0dm2MMO9urEhfIcZb5QhDY
IY2QFs+MtswNgUhiCWoZUIn/+GEOl/Z3Qlz/f1xHqJpV+LLeb7JbkT2FYpGj8J4Cs+VykUCpvADU
odnV9F6wXTS8ukNYldatbu9nZ4hZivp52RRqFWg84e5zm6jchs+sq4HvE2H2e0lJo4ZRGRsW/VwR
a6nCjUlLzfaWOt9dhiopvCsGDpuaA5lVrIeHuBgIdAYf8lYeejW7+noqG218SnQJW+2LY7cydvY+
F05RsAZBknhcK+9UHbbXFyCSfNVg56ef5tKM4MT0B7MqceOoxhZUgpi4Pc4/mUJcbX3KAPeP/+cY
HhoB5G5ewmK4KcJ1ICJD6KLdovduDmou4S04+itXLaJRpv0T9pmtGIKMOd7Tj+7ksJl8sIJlk8r4
q7NnWdWwRBynaas/2WcMGu39n0uPFZN/FFRne1T8uswV/wMlv4ymS3PmH1GDsDWgVjTs9p0FcSQf
A1o6/z+MDilCJMdlxT+SucHkIykOHJo72Qyc+izj2M+pXGRPDGOI+sYSwDDgc7gZFkmZ8/GmtH2H
w5VCzlli/B5irx7EFBP9+PW9bVdRVNM3EhNBukMY9CaokSd2itOkJLQg9mzCO00iUMTB+OHJNS2l
lpevsz6p1U9dXFxXUKXa249R0/jpbO456qsmqswjLgw9dCSWi7l10KVOKgdjNYZeEPCMk5mNVKlA
PvVzBFRDkYE8N5j25uvAAxhuKugVJg/jyG4PrInld9n6VPwxp4xMUtEnuzXrYC5CrEd5VkxCR2id
9f140pGBmH2OKhNoNKqf2YgLVo3P2D0043TcR/c6f1wxZaCmhq1RaBiVmheciMdHngtXEGS/nbwb
sh08mauOotdK83mTjqO9Ye2b68f7YjCXBkUB8LpB7jGzGP4zJ3yCx8EPnF4uEuIu+OXE5VtRreR/
OVfW9FqGsaJ+O0FR+4dsjROhGVrVqdbTXVyLY6QoIlHoAeMQoie/zcnGzIO4cxbGbS7Q9sVgzfF8
drXLNqKOLXS3dBqA1HkoDG9na2GN3GDt7JOFC9PejgZwZgXrYyKs7JXZ/LeC4G4M2pV6Pu+TZwHj
RcbqRiW7t45Um3vcKnRSTaVGEaeZ1H071dk3qRiykHxh0k6qMowBeVd7pAG3CW8ukdN+KUiLQTdC
EKfGbacylKqf60GO6wzpP/oO/fciLE7L9xGlI6kvUhQRwczibBwM8qAQnoNzvefxctJ4EGz246te
J3Ez66zzdE+Trz9nW4HwDkjn7mNU9n/qzvz08C9RlXkLp4SqYVsw8IjayN6/k0VGZvvoKTOR70Z9
P8NwHYXGqOSMRPpq2okCxFFSlIpE24Cz/a9J7JPp1OCiOucsS0gWG2Gd+b6O40CLMorv3RyuPRvx
FJEDny64AxHd+WmS9Cz36lpuIzssIDSIGKXsCDcOWo0g9dnSaOQbDoSlF9U9RdZ2lxy9zfoQpF0j
ZSPmA0m6jKiWPUXK26SwMIyn53jW61HI74evfAn2cDvEb5Lt16W3qoRByE4tAXHrt7edOCCbb4BJ
XmgtiTcODslhskC1HXQer2mv4ZpJ2H7Fr4mauu6h0+VOzDb+hbt5wnNXAHiZ6GlC85rz1ZDmi9K4
B8KnSFf6dCIMzmulaqTqYL10E6W7YALjN7U2aPTLkvpHcAibiQgivVD3E+NkAT9DIPfcRc/czdOI
r9MNxYZpCdEiDnxxft0RxNAOv9+lSMUjPRoQ3ZVW8+3v4W2b2UgYHg7PLYqAT6sOIi/3/wBiH/Gw
ckuFdnnBhAVwL65bVzwimdTSUUDS5ACh29L1siuCK0VjuOA7JqKfYGjmmqNnRnS3Xn/3YvOHixpp
AJDR6rd1OomvBAopeSuQJLqYYuyWy2qJtf/lvsYAgBOAByUst7biJSF4SfzFAn50Vunb01lyM/XY
iHQYV0REkCWF5MJCMtajjTqyIoAa3UF468ht/w0zJYlMoLGvTBsSyUFnleI3C7tidmT1AkFE7/xj
DJb8kofeZMXe+/CKynNVPvyyCoDFJ8bF1fqRUb+rwReOhxUHUb6frkNIwKsvS51ICtzs6hxRZBaU
6Ltx8p9WURql6KvxOrnBNB+ZNJZLGeiSIa1zOZdi4L3OSU0jG4er/f/hYbrVeLgm+IWejHebYXto
AZLqmnEnZkCjZuuHx3zZ2UyZMCAbKs/S1Omg/DWTmsJcbeEj6FxZkypQnVjC0DBZW7qsvsnwhHWX
ebEUMcRkb1IeE8C31namqHxx2MqS7MJWB8B6QKtB7Li7OZXIgKAMsXc8dl6STcH94pCTdx73aNOw
Q5LU/tKSARdr2v3Kog52KcrYFlJb4CmRcOo41/NNf9iKM3baKzcpplldGRXQxhyTmqrrcchHeubS
MVykmhctDQIkcxW07/y7ETxTsSHxvGlyVlmO/YRLk4oqIE3GgadoGyBYXt/FhAX3OX6u+JeG3bZ8
qdkOu+AeCC9CCZ1te8H3hZEmIsv70WC/vxmD/Uwc3DZjh94ZedplJlB1qFsfJeqfij8iV8byO/pn
PUi4aMWDUrZSY9NL2TT4W1Knlz/gnaNkSSzJUTep6cTGYMtVkqfJNGz/lLGH+Jlr17Xr1m8y1osn
DurdQdSWhcVKANq5ZrbpOEJAaK3uSgxg2sG0VG5NmLPTLjVvtA2En8mG0s8h7Jgwc5Q6gU8BYmIl
ezQOqn990NB061FEj7Obc92wmxOmRJrdkjk2yIK3cNvtvObCgTnQdo3CmBBB0eSq5otCCEDHZF7l
CjY9qRdDrpXNwo3aOlzKNyQaHL62ZpSSIGftpBjRDBt+S+ueywXO5n1NDOZ3qXkAYvss45FZMbCv
/LgiZYdBZXao5Kg4kyvDmdbtIc3jilAJQmHSrYqFl8Pw7RhY2B9LEWEd1t6KY6y/mXHRYpEPZe2C
HKX4wB+bydV4RsI2YbBxe+Y92gVvLtmllRY3F7qsubhAMQitV2esc0TQMXLa0StdDW6npPvi6lq0
WtRb28mWFQ/3tbe7CLaHfZNmkueOEUb1zg3SgRtDaVB5AZHr/9PTNWg83aofET0wEP90/Wcz4gtp
WNG5MR1axWsGw/55NvQRByMqxzsSH6VqW1UvTMGJ+j7SqjnTZplvtOOdtjEgwB3I85P7VYw7Yy6N
9osoqUxxR5x5QQLS1yJiVwGi6lzGQw3oL1+ZxWaWAYK7WUe085ynhWiahffRveijJn5U41tnn9Yh
kD4xTdfIuKWMKOu0VTz3UmHJuWIfjtl3YUi3cpYQtOrtzt9hrWiu8u78irtu6xMHmOAYeLRV2M05
MyvKf6G8ihuy62NUAOVxfXiCyVWKAtVsk15DeXFDr52bD2/XmdQqGqymktxtGZaQRz+mAd5xpfvz
IiNffa9+fjo2CxeN3Z0PMOJtsOnFm+SG4BAX4ygImPWSbwHj8CQZdt0tDFW+SFdJyDmYQCKycQvG
d/gXxVYgz0dM585cCpaJyaT6jyfGeeYl6IC9t34owKY/Se2bV+vKqrpdbzMN6WjIFcYY2eT580DY
0XnW/nqxpOA9Wr/l1U+jetP2cpf3nSWvU1ukXKgHCTJgpoDYM86woh6ngsGISY8IUrGwste2owJ+
jJBYVTJnBdkt4eULOty6wFw+9OEy5+soWgcTJymfVPk0ChUayxdHWmBoohw7DjA4m4ut2nrK01t+
qKr4Tmhmvn87BW632AXIp4PfRzzVudgGlztrPzW/YnnSD/XjjUkDQ67Dn/vPqAMpAanYVDohihHw
TVvbqOWE85LyvhFlgHpInmiBNXLFZGUi8ApD0E+sHLqhH4DlBFnFY/vOcs1RXs2PNYA4M2GsAIFh
txYKn5DQjWlIbdmznqkG3dC4l2ld33bFuEFOQAWrGc/e8/zlyHXxuxPmbuUwUrPLZNkNib9HRmBl
VVMoEbCE/g0/41dr5hdnYx3pe3nXbpI6aeG3mxFZ1R9kJiP1E5mNhpQnWSByoYj9HhtOJ6Uzn4tJ
zRtqo92Tw2EEymOO7j+BuXWa4xkYZLGeptzqML/4EJWvCm3oj8C0dw+M8hkgz7DMZre8kcaBYz4I
0gVrKwInfXcg1fDmZDwbcJimTFl+oApT5mUM3oBGFRLSl2fWYh42K+MDFyi9E4K2QovDiqu2h9j7
Q5kJZweOcUFkxSXnSbv8bH1/9Q3Rz3Ij5rPlTCIfUq6wCgMbXlZSEoaIoF0osUXpik7qGLrUxie2
v/8exv2zqq8oXuwTLIwpFgLutexbijgWGjCK7vRhqszmcYtNHkRtBOMfkriZd2DlYkzw6bbLNHfZ
OQL7CUcMz/o+vcUTJaNcwXuCKvZnlkiixm2zq1do4+Bi4bZRNx3VC+pgGvRmf/ADIr5Nmt1cc8Iz
G0gLN8QdJIHNwcN+RtAlPMZYATh2MWacc9mY7CvpMPRKNuL0LhMxGlTZqOj8ALPt0KeqOJS1uwoK
R1oXHXjHb9YR5e5zS7U/Z4Ujp8Lzqhc8NQBLHk0TZoPzynxzVdAEMmsLpFoyLZu+R/us+0bv9YGJ
1/xc7mUOksOkSFJKKHUvEHb+7LQG4vbQWwb2xBdpl3VNXq2HU8YhXthG/UzS7RUi5luSRnaFqr8Q
bDw52SXfD9RiBNSOrenhoIynPXLrgQaoaVN/h1SmvXE5yxQLXHfb4IBJiyl08tANmIDtsVt6W8lr
Yt9u8bNhxy0MSSODgUZk027M1xaVo9+RNRm5tBeChVkgaJDUP7uha+HdWb8I36yl4VfJVvJ+gTUd
W23ndtFSj/0vkKOOBq7D//6sSQpDhZYV+gjt4uF2Mea/TBWonvNDQisgUZfBwmCIjDPSWmf2F4am
0UI+8igR8s/w5QVNG7ilC7lXCgOY/Cl3bCdf1+x4aYmxWdmWhgCE5HzYeOlISoRQQPxQA4hAjZiD
iIqURY7QKWHxjR9u8RmLghNftU6Yd/C9Hv7NaIk9WL1Iqer/crJ5BqGYVJsq4KE/Wf9EKr5ETJQk
15WXStvOs43rB1dzWwDvbafd9UK1d5eFcf/q0te/P6fXBhdvA2NWISqtXdpIbwejSPqh2+hrUG2x
MGgHaR0z0dDHee+OEXezj6yC5zspGaeQEEmcH9C1nJyc0xo6w9FCE32t0vj+2l5I/QO2UXno5MPH
g/t1oJWm/JUCV6tS4OMX7QMcI9VuBup+Ghftb7xQaTj8r2KsbhqjMQf6dtm9dyrTVNoLo/UeIycH
afBLs17FGoo5qio/jTw1kay7Y9onaoQ9km9ij82CrEMpV8/zZgUFwiO7LEHAr8P0uXT0e+a8+VGd
ljBVpW2JZMIPNKWb/ddUys4xyUYmTn0caeFo7uUlQRq2PfsvJXByIxBOo1rG3aDNlcCPqGT/05KX
iIMxzzAVR3jVPVk8/pl2cAqk2An+a2h3wJH100a8Jjj0pYmGoH7a/xYHFaGpKIKWE9hOgmV3O9G5
tgp5oPUBhDplUgV3SwO0LSbDXe5vdXYpAw8616AiHN4Xh/LmUXFzXWodaeKgzOna03HoZMuRLbCl
Ng/d4upRQVbavbufI9KpuUhBS540PmnIOhaB9gqPoq3Vf7AQJ6UQHfLuEMJxb0KXJly5pTpxluhg
Buusp7EtOosB8Zn3YFLMlDf2B7bZdP7J2qPtpCLPSoiCmL9siTrTXo8XA59xCOWa796qA/biARYC
GD8dAxNBz8pQtlY+zXMsB9+1e0ge9UFgVvRq5BAgGOkF3iFe/FaUs5qYt9tRkvsVgs4YKViMZH4v
vaaPJO3ccBBEIx2sb4i8QN4I/J8xCeRDvEApi4429lqThtEItqMj7Q4KznWYDe7CHamoBenL17Ie
tY2bUzZ2o+eT+tJtytFVkN7W2WVP19oELd9qfEV84wouAVlnTJ2n1VtjntFNYLNwJbJoarTikvbO
f5UPB0yajo/9pZs6yFrAygrFwjaCf+BqSjNC+JQLp5eyl9g8BfaEBWT9PZaKElJdSTB7kX9CcOTM
6kFPcZXeDRhOyreKAJgoR8oE8Pm/7wr1Jc+LeFRBq++YrRrdIUety9tWi0Dztd2Z6PKTXCMl1Qc1
a8jKmDmc+8FBGcdcPec6rH+l3zIUs37D2mFLMxsXTfli4BT+ba//i15+LgUA3L/4BRwpMRgFyXsa
dgE8m/tf3nKRO7R7vwCnYgfFp3PI6imuqG38GSflPFDjPZxQYZHun61nhFyaBl6Jgl9Zde0ZnHzc
5rbk8MAa4+lA3DD2zlh55hd0aWSRsFNrjOZmCZS0UfkiJ1wcrlpplnexOL7bIVsqo6DlywVnr2cx
+pPv/1nJuogZphv+PCVmxs4fCbXFBjjNEWd1uXK4ik4Unj4vqBxvL/NXhzhsDvQD9KneVy5ER3p8
36WiIJEp84OL9Uv1e1kY03qBk3b6Ft8v+aU58EJk1L97q1NrwSiRHTv45MWQOFPIS9/i2i4xsZDd
03kHJ3jUV/JFGXtJRdBGGH7mvsywTywDgAH4ySQG5jBBGSX6ELhFVFAKdu+9tLQEuwlmDJhCbZXp
YkmqELX+hUMykFVjTs5AaXcInCC0G/UlvLrHNJWZCeQi9WLDgxkvzYoVBoz+xi4PRBkDilKDe1FL
G6F6xeuptxvMrWONf13mdmA5hGeA3bhYQr5zFKQW6w/iSVBsc0V1ZnilGeOyRKxuYI4qGtksURgY
eOg8LqpoqvZKSmA6yGiGYToLsRhv8OAuFyqI2mq7sHx5xsCYsRULpbTH3ws8blfVFm5YS1imrGlg
BtWgw5nUYmf0rYwP22yQaTpZzs7T0yobeJv9M+nIg1ugeWswIlTS0NaFywoAsCRDA/8xOOKiKknE
+/0moNsZ+3a+oy8F0hteNMKW50d8uDrjFcxk0HgG7nzSis9gLD3XHjFCjZxg5hh3mlT4bgs27tEG
IoOjyT/QOSI1Y3YqUiR1mrAqRFNaXwevy5cv6NIqmhOYHPlqom1TpAuSTjuzOjfUHLa+dog4/ARr
+5rvRQbFdPTLjiGoPKX17bfG5W+MO8L/SgHG8K6oJZJLKAKg9QwADLUvhNQ44OY4KV75vPHQ8ueJ
yso3XDy1xNPBkctcfR3DA37okDtdBhOEzwK7YJTUCuyNPRlr1qYbDxT+89cxjmtZp+p16H64HoPh
6Of9ADpJ3ARzogCTw0i8M1kCABaQOriqG9LscfDgvJZMw5KN8pI3A0zMId+dJDikTMN7V0PSoT/E
PsBZx6zPrDKUH5I+UZ31BCxLZgQRXe62bknk3OIMG1AQUYpdfqhoN8o2vOxpS86tGHzuqrUcP6mq
cLqkzfVSQcuwL6no10p4tcERSaEj0vwpiZYRDeORd5ecreIKhODxVEw7MkPtzn12yyw7eU32qaQq
mzQwgFqGIOxABIUB3HnFpqehNeR5jyxdKIZw9K54B0cN1U6FJyvoaE1Fu0smtf5VlTYT5gpz1qkv
vabjXoSGio7Dwry64YLUcpF0W3Cwj9ps8UTIsdGwomWakLmShb3ZdAmX8vvDlsX2ETQ2uEOizrj8
G7OhImYA2X9ARtdkSa729krx22efnQDP2YG0qBZ/3cAQ6gytiMKbtYv9DkviPbFk2JLiUa4n11ox
PzNPgFlfFbVEoH386+C1sS4y0YmerZGVo3rkPxINYGfhKNZTDX28ZK64d+B48CM1I8ZOgaPagClL
7BgAe1HcdLAlb0dtFFcV/E3xivR2hRR0ouKgjlAZsYKSQBZLtl3+IIkZ6jC531Q2DEHWFgyGfOur
hmIOSEY0PiO8qDPsifxhXkhJQKKDc0AVLcjhsG9SAxf7P3r3IvWVgpIBjpxnboEOq6y5F4SJms1E
DH9Mp+MDJnSo0POvhYJN4kENtetbXJ6QUcQqyDIAhb7kmth+5Y0lK/757w5pwFbcsT8seXiTiziB
WTVlRW4e7NbU/qXmWBADW8d6baAjh4eIqumfcDKsi71iJ5HN/5ccxDpOQaf9NbZFEsN03DOEc1yX
Zj2f8dh3BRYSx1DwWZYOO37/tX01ubNX432XDfzDnuX0aJ4jK0IrA7tX8R+PzLed7lr6oej/ccNn
E91l9LkAAEsPnqIEL2FJlKOF0MrxfIlZ7Bw6yjktlgx9OP/DVg6x89mksu91HXhrjPJZEaAjIFBP
mOgEMCbHNnwhfUPRdgdyE40UiwTbcwBINUrgfMGpq2KWiRCwRVg7Jt0u4YNUCv+JILdMaoOxVJO/
NWYOu43pPtwg0ifJz1gEPEcSYWHSTed37vO6u1QLLT9WB4DPxRWkb9QmsWonowmZrJqEVZrziW+8
l0JD4eTDte9+hBC2B92IDHcyAltzbdp7AQuhzbdkl7TLCRd6lW5vRYtwM1Wm0wo04x+lxSE768JJ
ayBuipYBUyZgAO/CxxOIDkbTg0iGQEdZMEvN8oTMWpV1uUVGGR9xj5bXSjz0fk9wt4E1adEUvw49
zOWdM/DkDQ6C0qG+modpAzFT6ECCLRwJZSKRpesg/uHC7lL/oqn217AX62KxHXKb7s39x+1cuoTS
ztAG/0y6b1aWYTEE5/yyQb9mXKjXjvi6q7GOeK5+/TCNGbLXzfNjUv9jLJpw8y8IMj7MuZMGmd7U
7L/GVyj4ZzRns8XlvE9Cvjycf0UWvBq4/Cqc2zHtefFuDsw4W8/aT0HAGtgsqsyQjXRrETKLMWLP
DBMFsNt5iHcx1Wejpd8gVZfRZihF+xljgeVtRPmWlu4c+TU561wax9j8no3GJRnRiVrH7EjYgDCu
Ad9C/3KXc3QShijG/ivQ7Q64yHbKu8Fy175TXDZVhopBMMa+xubSC4xao2qvCbYeQBVKNQnuyNXf
hLeuL/b5vY2hWlL8cKHCvvd6pyLR5XM73N1c8P0fhF3DCcuohFl82cr2fbeqP69XIFEmKd0B3lTE
z3BicLvcQEpHktFMCD8KzYPJT0vlMOz+1mg/yYmMfHh1LolGLjZ2sXOLyplI8bFZ2nApNxZUoGIP
5tNmkuLBzfgqqRykjILqVMj2TPy5D8WGwSwdHGxKbLxGcZbh/cn91dJ9yVyHyG6ZLl4flzJBzVNH
fJQu4MNPxd1g7sfZEJR/3W/d5OrcC/Jut93gmTbxJ5HC5QlSpAn+1YT09uLZRbHUzjcUf+Tje74E
5KY+cdbzUx3Li0c6EtHTBFktUdaZG9fp3IyC/J2BjfqsY/sl+ezY5ZfsLbfPqcNrgz6dQZR9vHsH
5L/1xF9ezXlwQqht+na/c5YK3Xkrw+WlB/a5uCov1XX3gKAfKM+aCDuirE7921Dp3WMbDIqOoAPU
wAx6SkyOLEFVgq4T7mrNqsCaM5lVwNDlDcboWX406IqlEYbtIFcim0LL4zyVVRyWuzrxgfMSZdnR
HT9A8F5M0nZWU5wT1EbiW/uppn1d9Bmk88UE+lbxDU6POAdnw7RVviYuc1fWSDrzleu3lCWXJzOr
NeRUxj8IeOusG0ngeYaAhBbuJFcabdreAtg8hYElofN4cu3LR6J9YyApBZaAeb4Ji1y2nQqM3xQC
RHKRN+1sFmVhuavpWvDSNZKYd6ksme5rfmCY9hxpYfXrw0b5ZflXZnoRO3+RiRXNFbjihLqmXf8n
GD03+QS+HEzzC7TJ9hBBDJGiuut8KK5+OqdRnPfxxUJGhjmzXNbN/hCcx3Csve4BX2ujt32U9uOF
29DBnC23cyqlIoG6vs3CF1Bz500UVHsj61NwZkPaLKfg2DXu9HNnlJ0BL4Cgh7aHvQWh2Jd1aCdG
wQ6VZp8L4D/gsOj7YJHq8GyKCVF08OLTAdl8UBnxum5P//Poe68rkbkLi9Ae2a3/kFXXJ3OB8wWu
Ijw0W9v30bfLYODIhrHXiH72YwZEPVgCLTZAR51KBarNiqpBjVj0P8qovQezaOHJcBg9qyehZG/j
GHNjBwV6fwxA2nEMSeO3M8Di9XXhcqJI9ZoqDwiXYMUYygmAc7NwTr9jsOguifUDmS3LQGEFL36E
fYMURwQgC4GEqJc3cmsk2Y7+ocHmJJtFzDB/iJqsQ3cXbgDTOJAhoZcs2MMCC/kwUTVDi6OBInnO
wsrj1prNqLJoJJurgEXTVrI2dFnpUyQHHuz8fk15Qj2N7e818BIlos08dGsAICso0RWk2630Uuw0
/X/qPAflnVPaBJZEYZHdyc9HNuoW+FosYoTNZe16oDu0PEG+cTyh0Cc97mBM9xpfhPfvcsrIv5XY
XedSPX+BUJSGkXSQJsRMy8juVMPYQEVkjgwysr+3AR5nPUhQBBzYm7WqO+jxJD/2Lm5blZl8Fyli
JW2ep5v8n+SsmLb4oxF1HBEcyWjg340B5YkQylUfn0FxGc9eJYlt+UcMHpj0ZFvd6FH6Ig7mnBAB
l+/WyubpbFDyeHfRSCawsDTS2yvmJ8AV4efsekLhvrlia/VIXBW4TY8AlMDFV8oudgfOKoTTJe4U
33aBzCPa9egQ0EUoIjc3gR+VtG7sE8705LMLSD0bb6JVEvoBSV1X1j9h2NvIg0xW6cPn/h4xQZAz
JSzZPlGwXg2h/jGFqwbt+c256g/REkPdwocdtPLWB74j6aVwauUoyyXxBQzkzz3Oj6TdjDLdWI9R
gkYLGZEEAp2AviPKODT1LlXL8+RYSEitH0iFaHGKFjE1Z6Ras5cAaPSefHz2Ap7KSR9cWLxVT5QY
DFhSt+g4T3aCJITY4TPgHasLvgCFf5vjCIhSxK58QuKf7AnXYF0KdpONGe/6oOZeo+Sf4OEyRIew
ZNEAZtaaykRiYIXh2N59hdEkqFepCPzbH0JJiQSq+Fg7vrBLNA2cLFM3+pbRmxc+g/ux5pogRrov
1r4OBDZPBGNEGeSV4ExZeMbn2PM6jN4E1N9edZgPYXz8C28Ho/2v2DnkzRseCHV+tiHUN9b5M+U0
aTdw0hSuinwEa9gbt3bBg2IrHvf1giWIgEqfCkRXiJ5XY3QvR02OPBx0g6b8m/KuORMorxiKfKT/
PAqwrP/O1N4qXxCn2wbtLsK9IgsSyY05XO2GYplQay2HJ0CKrvVWZ6tscnCifRNPHFTevZ4a7JZg
UqyMGqJO7I4vmvrtyX9W3nH/xCRYRGorcKk4Bu9wugK7zjC3foAwMFeWZhZQJxaTW7u7jScWMs+x
SbqNQX1+nuXcL1l1hbcE/Ag3sZre7wDawPo6QWkOqcSb4jKENp5a0YFr4OT6a/Mw3tnDjHyOI9U8
P28rNtGRRxeR+EPwxAl4KremqpReKXcomVZ9Jr5iARV5BNZK2T+Vhmm9DoFBVuhMl8/6D7c3xt+T
A7meKIcgJBvLy/ejajFTMZ11a3acHPIXAVaEn8uakRYB8sUN2glXHsSARgy3usHRfxz2Jzxq+10D
YzqvcKymLksGbhf/MgiiHrEqmKFe1OOenOYbe6zbzuCj6J4yJpkWp6QmIVoAQButxHKnJJK9RGis
mgf/wc32vXdzSqZc2RJ9nVCymgZFoAV0uv6+PFgtYd/VP0KR0AsjX7cNwxK3XmqtYUMvV02z7maC
AMXFQ72aBV7cdK2dhgfXifiQDuxnlpErgSyjiDAzpVM+zmdHngG3GB6HV6o5s/BfrvYQWR2JK+tq
scgshtyoH86/fVwz6l339sxVoBhkhbDVbWrKB93pEQf4SlYjLptqFs45Us4doh0ZkjB3GXNXxKjP
dFP4h9IKZlKd2j4nKFTAylidHfsw7RtXZKHAV4xW/KvlDEoesgLmrNK2DESxJEbMWzOdRq8Dy8DY
m8VRPES1uY5TkpgRoYI90+Xb8gxf2+B5lmsd2jwAKODKd2UyqcCd9IvBgPT1P9gEbmlXdNEdpBhr
XffEiLG7C91lWIf3X19sPPAGF6SWjjsZGgc8TiE9e6f5G0B0zNkScdiMW3C9r/exKTtUUO/tvSeb
RXdD8zGjXBqWpLd/ADD+/t2M+w97dS3EsWoP0rXdYVkEFZFgmSdnk1hhrHoxhNAeWvSXaC0JURnX
uS+VJVuyP9VLHkzD6NqifhLV5pCAATPr0PzMdMr3sBZB1IsEa7x4E7PlnOOMDqOk+RIM4gzd5YHS
Q9tOUjGYkZPbEzk3svMm/HyLyeTgS2y93WFbWHP093/E7KyUbhexH0J3sUC0Ky7JPrpTWa9l1rJO
KSfMBATHtt3OeaXkaN6zHCQ18LWq7p7tzjwJm2TIW5KtkcbqMoEQleuLLjMI9P0GhTUTwRtB8nRl
Pkiuat/ZqF/ur2y9GQ/REg/6/gyYk7OEgY5cpLQCzkOLNl9kNfPdGg+V23Uvj9Gs/WieaF6G2GtW
AFVTFDmXggLznYqo9JXp26kBfEhnh4ekmmscdH4lbrYy1/yU8Nd2Zd0tERcc/Y93YEIU5MUkFLqJ
gIScWZqnC3yjmcemkRrxn8tJH5HWPoKklDIU/bMv0+jikB8x71jhaD4BLsN7R5RLaSj/6oiy+Jds
vRHemHQ2Mz0L9beYo+3jzh4Ds5gWVchruQO8VUvWcv0HNG+qKa2r419VEoSkIVhxMHACM73SGtRm
D/FCqzZK15zvpcQVax0st5eJmbzQEmgk4zQrinlrAONq2qn5Jv2tv+yIrEm/egy30b0aHElufnS4
QgxWDBq0Dcw4sS1NJDzOnIai4azo+9Ptn1925lsv7SLX0YdDHdh4bRnOdbIPwjdqWSe4F5vpMtUu
NPwupFN9R8PaqRd6P27dxNQJSkzDKn4BhuOwphezoNS3odUc9D1mj3oExb61LzzNtXtsNjDxAFoJ
O3W/xOY/Co/QzVOAoL67/32FOaz2ESuD3eToGs/DJrULvYFoAkpkvULs6NPSAXCHGOOHlZaGrur7
KjpKmmHM6VszEqGyLFUOJ3kBSvZavQYQtCJzjPs5X1D1RvX1xore6PH83WWCvtO8JqJOX7WOlxU8
pstVYv53NF7jhyvkkE4khl9gcidvuBpzmDFBDljQYsjmO+DFB3YavnJPiJq2ufnn8HguIwjqN5oX
DTbYJk2wj8u6TTPEXrfSlUs7oxVoCCQF79lgOWuPeiFORGnOUx5+mjZyHJJPof3sGvxJW60NZidU
40I3oGjWQjN808H+BDVbWEc991+sLs/h9e6FH6BDAzxEned+LJbHI9eezdGxIkhMvMjVpNIeltuT
rQcf/cKPQcZ/nJVQpZPMJjArHsbt4xTIh+yCyappltgodDIqe8rLxjp2hzX3xHYec5WMlGbpCmqi
1Hv/LjH0//k6OsomGIjmP2zJU91umwFrT1dav1SQzWJLXFF6iIClZ8eQJXsZbRlJdqv60MCDI2HZ
1W+H+vRc+u9jEOHxRzza+cDs3TmJckXXBahqZ1HXItFRNkh3hdAQQiXFgRXHVeP84cAPo7C+Hfrh
DZ2vkW6978EE4aOKZkFngxMI7cMy36JqyGo9hy5gYl+lb1/RD5Z4vVqXfcMaQkiAqUApE0sQkN/0
Fok8HwlqGXaIzli1kMFwEubLtZ/dZJG8AD+5FGj2UgDgIRmd21g+aLvCW/rnIv5j32wROM4MYZFY
eod/uA2RZ9dSk8hVCEB8gcW9FcXIXkinsGlhiM04HnXdWQ9ZjndQFLC0rlgeCmthslKw4Q1naRfN
0xXix5NJGs4aH0Fnj+5OSsNl0TIcmY0UTIh2M9xP9WUvTPG5TYxT7IoSIB0qSn9oyubZBQbjKwEK
o7w5N20KUxSiSpR2xlTSk4gKnB5J1CqpGGPJ+E9+i04lyY+iNFO99FmmAEwXEGUhOH/xZiadBcan
x10qLt7ciXH4Cn+O3ecNd3H598CnTPtDf7DuJac5NSs/nu8f+pv4J67pTJjNjNfP0HmZLZWc0UfF
Xo/9vIFA2k7yT1mn6mLL1/qYjM08aB91cb0ls8uJidIlNoRZJEi95Va0/TqLOSFWG2SjHN7Vai6z
v8MCfY+3AwRWMIKhEPaNf8Ot1RLZCz75ZXKwKB0oYQ8fSUu18L7TMMLKW4ypEYBHY5NwieiJvpqb
Wil74rJauM61AU8WgRD/DK5ieO9EvUcztPfhvKsMejb5K3O3Gp4nhowtvNFHplBO0I2nVzY0fZQ6
2g3ZE00O+XYflEvRfQazTpdHok7oWdbHeq6on/SexSOOj/IEiH4ptkpkAB/r8Zj+mQEc7dKEHUPH
aEBwvApJ4Y/l5JBOvAnDIoGTNGRv1e4q97VHwiGi2mx0uXoIERQAQLAaC49JwlYv2i7qE0I6puim
Sh6IhqXYn6CXWpFy3TZdIJ1UqMcaa3qZTZspo8zsvyQwKhHUx4AzUuQNax/Z2T+SE0Cwr/ZKvWnR
a7L7ipII0x/2JW2AcDB5xORx9V1kHJWYqoq3kLSIUystCXuJA4D4hyyu8pr0xClmF9h6Kms6INjQ
/r9nTgP5xGJCgiRsTjvNiDPb06Bd4cSv5cP3hWJqDsbVYy1jQGlTo3r2L8IICFSYCp89ap2wIibw
4A/8EU/SK7D4RtLizTdW59EtnjGOOQwBk3VaAuDcybIX7ZqWVyxcNPX+PHiSvik16kyYA78JB4P+
cGiwarL0VGlzyMuD86KCZ5vAbunVfSdzPsXNGPkpbTBiSgvCMI8WWe7+oeR4Ixk6wamLZLr2fz32
9Grq2MWhA1eNyYGpbshH0zRVdLkFmylsO1SgyDT+ALJqGQtTrs0YHAjRu7DjCDo57jlMy3c9/J0t
dBJtvTUaEDD+5PlJ81SN4bj9wGeOH8aWWJoo8n4EBB4Visy38zXX1eZECTWjy03ZS+29v/cDihAH
nNFlGN/zJ57Fe7Lc+HuvH7MRRW9NcTcNZaFCIplbF15CxAv0h1SC3YPDlOtgqFjy79P4DtjOpUai
nM0gO7eOuSuZewz2BvIAIBYoTzxy+hTweweF7B9b9Jsorl9rcvdV3MbItYZKlM40U+wSo3TsWXUr
cu1Edbcv9FJv9ICrvkPewZ2m/edDG1+CST3M0Mf5GKJzf8v9q2DbbkTB9T0/LnXiHUQY+5FY5lUN
5Fwm/3uP+T+3samZaXxKwDyGgt4jeRD4rEpmeRWfT06H8dk+ZcXQKbyCpG03Wu3bK3RtMNIKA2NQ
w9KAeStlc1/rMG2KAp0eSYoGSRAyvAIjX0nZ5hgtwLWmvrSo+Xi5Nz/gWTzmhX3fbMxmOZL44l8E
enV5g0Ww/I2OGgposaq66cRiVa8teijFiCd9sPyu5oQVVBCpRYrsh1lNP+ltsOPSqACThW/Sz1c1
bCxWP2taIPX4Ej9l/WCY6fbsr+pFCj8n4cVSs5nRQYq1kiUlyMfgwkef+/Ny6fMIktuW9PDrAYIl
XvucI7uCwa/+mmex8pyvXe9N53Nlfmg8GPdze1SARFnTLn+CW6NM9z02GmbrJrLYDDvnml6Afe82
XBTV7WNpXn7DAaWYsgt+/0oAp3h9bcYBZ0zvDZExW96CE/WeVy9wqamEMF0V1acQ727BLgRQsFoi
3SkZLCyciGFQxiRzYT/zKyHVCU+W1MyB1sdI0gPad45fNG9xmFQLB0FADXXvrKtbWbHoN0/M71lt
XDwqcC2oieWDYS6Rh9xTUQNhEOiTG91Dp21yaBB2BQfj/sCR12+PfZOsQL5dzj5Fgo7/fql1l7Aq
+DBxa7EhJPauqpEXd7W16v4xTJ/2Yk4QDl/MMfhYwRtdCBDpl3eDZUJbo/a7C8Z+kOrITFtDIubq
W1w/gGkKN3rKZqgK0c6tfM62A/oqZyHpK/G+vqpBXJg4eGNTOgd7sGp5YNhXeeICmbtcT4IkinOT
F1zPfABhxeH4O/pimmqo+Q3mM/TxR0ykyVKjYm9RnrKUgqVy6yHczP9t1WYt74N2KqpTaM7KzxFa
nuMqwpRt+hSkP2dyyLCVZcrvbZad1BTtEzOsZhf7AkByfXmhjUIPb/9r2RMBQhXJmVrn0yY4NS92
tmcgmsx0gtd5L6XR8DquBIa6O6y7yikT7gXPFeEQXhiKX5vtOGJxag/GhLmCL7ZG1AWIngMTdA41
XpP8+/Xf1Xz1Sv3QZeGzwc8QABgmaQHhHkcg7mAxFhUoPZRvCDh7xwOYCVpo4DBI3Sc3VbS5YggT
mWzASXLAe/9Rv2/fYBJxtxeK87uf9w7JR8yRaeg4k3QKL+/Jo1/Y5KVD2xGJnOYNyWDAIYwVop5y
8lhV+rYlTZV+90b1hrIsJ7oO1H793VLNpTvSWBXffi9BhibEKMdQ9Kv07CxcX06/k1q523csT1P/
qlbGkT5ssu480IGoAyd+vIe0Cuvz1lik39K3QfS8mzhMsVLEvnlv66zh1CItmS0eKOUkHFYSg3a6
lYHkpOOqHIu6cnzRvkcDK3zd58SuHqKHmGar8LsTc0trwi9lo4uLwXYVItOKfsHRTFPuLdhoFzXA
oiBPm576pUwQVhXLICh+elsEFtX3UyWG1xwhWRoW0xWcv8ebL+WHgh5Wd8sY1dIQT3QAa9OsDO1O
3wiYOL/NK1k3JL29Aa1PbD93fonkSJPzxJd2KnEMbD5J5m5RuXAUNw3AWF5Ko8VX6QSkz2B5IhHc
mjnhhDjrcyq3yHKv3yGlT7/sM4Kj4C3QL02Ju+vL/X/aQSWFamWKEdrpv1fRdKJiHRQH2dbdZL6T
uR6Uy1IysmxRYQY8XuIFyiF6d0gfGW8PWdXipsI+xT8EigEmwAEnZSFlu3xzIMaSwT++Xzgh1jfm
qW4SbgWy9XfMwij1PVUEECXoo9hRRvSZ6jOcUwDy8nU062S1t2PsLDT+mgOydLDgbS3Icre8S7L9
PbmuhLl5UuywcsT1AOe69VsaNawC47MVt5n14kUq+ocPx1gGJgWz0G3XMoGC+yIbgrNgzP2uO3lz
yVRJvSizhExKuetncMqQtl0AWnVys4lfaWFpqmhk+DJUOt+BxlsWTlNb+OhdodrNIrk3Gh08gdgR
r1/Mpfu/TCNL8vFEL2Y+vrlmrhCZeKdNIDyLmMnSMN+o5SL3cI3n21Bi3GFhYBylfYEAI4gWQ2vy
FpZgJqZzrUbsMTUMKB1v7gIy0hTwl9JhsQTe9/LKJM4gVhcys1yoLc0v0J3qvwd2r3FM2sQbk1i4
SVATaHXnX3I8MN5k+hvpucpBAbtgbMu2yy08Wb4uc5gN63u1/XYuwZ56d/+uVylvXexw6iZrsOjh
f3b85kltX3rZXjArxXBEAvqTVcju884X0QJmDIWklJEYE2FnsvXQQq4QRfJyqmbUaQ58e3UVXG5+
zqPiX26sYhPmxkRsLw/wxI3/GO6QJXW1rPSg5+1pwMyCXy12RbSO5fjTBHsTeTxgB3NbEV0WpoKx
IrA9cTjBLNh1Qk4ims2aGeLnLyhyW3ql7poFvyzV+T225Si9JXdJW/OBI5cpjEphDf9OiFHontt0
umiSKVLpDVGJm8gMwymf24fqBlDEZB1995zElEXo2v3hNJqVm3QMHMEMcMob/zaQvMEBiqotLGQL
gZxuoNSP9qKB4ORNT/wB/J9HjGjtagZtepEgKFXfrfz47Xr9Ih1bXkHy89+6wx5cC1RceqmIyhdh
xYtKU4rSJMInDjP30bE8Xx835cgQydRxqi9Q2T9mL9NbFI9X94eYBhu8Zot5p7gcDWpg+SPmZXXx
aTKmKpm/3RQX5hZYiFsJXl7dxDKiQzJXRBaa99oTXxBOAAWhpwwitdd8+XU2+lTzemaP3oRGcmKe
Q6i0c+LVu5jCNdlj8RHJ3dwvRo5w1zxu0Zs1yRCCha4fVmLsVUt5f3NrPqekI2K3+9Sv6LEmk8nh
gJCmqplSp808e4axiCUreA7ezihWETJzdiN3RY7j5Tdo2fG7VtHEtxf6INh1P/zb23eKawstdcJB
YgtOLDsw2L6n3PqUV/2f9u/IzXbDqG8kh/F+aR6Dl/Np5kPRbDgrCKa7rLZJ7RSQdplP+AqOq7fH
MBk/4gjalIkK0lBIss+Tpbc0GXUtdLcmUiXkYL/EgMETbcKKB8tzjS2ktpl5jRI7QBZxQlfhQOhx
puDQ1MFQ39UphymkmF7BsbAFI0b/XvGRcRfIglGyiha8G6Np0rnR5RVUXPdP1V791w3uAARrIwrD
N15a6KVLlt7ebSwC2RRJIboD5z9EeTAdk4j4t+nhL72r383KE+9cnt+xBMvJolr860rZgfFPw8DJ
feKG/lxSlTFs0I1CylKzzTT7EmquUNjTjjXzMDpUzBVhiR4cNQjmyYILjEKbLp0bEa6J7DanAqO5
9Zh0C3ZNf0pI/DRk2K0DPmXOwlVwoYPhtzWCwuo9Mlk5O8DmO2Y6NRLDkibxOUtwBeW7+iKCvoC2
ezWJasU5lyce26eSUfvR1whhmAxVfs4PGruk4kmNi9mPWKkvN/nZOxFE+NtRqIxjf++EzA4Ki6F3
lhPclnbwP1jS3CAD+DVHLz0AZpTeYgHjzt8vaXgatAlKCW021dydQhr8sYZwEwS8tIE7wI4DDmDO
6Q8r1iY3464/bsCmbUzES4xTf1ze5ODUYt7u/EqKO9N64nRVcNYijp9u+5NBXbpHu4x4fulNZ0wD
kKpaD53+EZN3L9D4CsFWPpV5Bqyg1/8qyIP5RxEiorK3y0+idTQtJeeCZt0ohueBAPjUQzw8Iexr
pl9S/g9/2VbyXETSQjMzWk+GJL2P4vtsq5Wkc+JoZRayC2Zoyh1brFHWe/AGiHmulgXwxDuF3PIN
BOVF0avcO3z49DX2VTpIGiNluGuv5nc5/dwmvPQUdt7R6LTWqJisx2KIALkEbIc2g2JLpB+VxH54
ZeUvncmIXtm6qLd8/TePjDkuKoidH1yUSJCO/5OF3LPLM88Aq0OBkua4WZei7Imk7+5r6hmZr+cI
bu3NAc7z2UWUIyh7Vo3hirx77CwiCJaS7UpWvkZO+8jEo8pQRu/9jadV/CBXxIWzPdh3wuNUvxA1
i86TYZEdWEIZVaidUwaozzrSEAnhjRgQYtt8KYN7PskAba5DVL++DBwZl19cwaBFieojDtgYib4s
gJsiji+bk+bfx1LOMhUgFswC/2GJwUQYvUMr1GWbKl6uAX56iBvIN6m557K7iIqtpVk+KjH9FFXM
ytYzXFbFCDgsLhS+A62Q5j6K6xBuRPK6diH4miB2GoeoCbGSm16GQ/IxxN7qeyEqZXylqED84L6T
KTf3+MM3kM9JayBRL7wKbsvmjpIuLMaHa6HpsWZak4IskJD9O0sU3W1cXQyKzEZZw3glC/7xxQOf
X2CtcyoWmiFF/L66hbv5miDJEtmkocLVVAz7O5fe6Z0CjG3GZ9Dajsl8qMtKgdRMX8rVbFMt3NIr
8IPShRiydzV+0EEPdnPbeZgUqiKo1xr0YFhL7jpXyNuYa/218aKpsoL5G76KoJsg1cZtkEQ/+2kd
7y4bvXlUMiq/YFZvRI+YKBVh7A8F6wBXdumRs74QwHIRZ6sbjTTWGKeW6AKA2oaD0cM+yTpY4kpn
CEEtdQDuUEQ3iYnO05r5KijQ5hu1UcLP1SF2vwX+PC1kr6CNxLGbTEjCmC76Bv0AmYJubJodqSv/
70pmDT04TxYH/xfC6S3bV6y/Ya24u6ofcCawB3ObXAHtoPaM+UBG/oCs2RyP8VeMtXBIxY5PEV2d
PHzwyAMQW5CiTcN9d7PAksV3fw6+9T1QfHNUhW787thv+iUDUsTiFDXhiTLvy/frDeMwz0oYbQuw
5XdiE0wJaOf4rpY+5W79LcVIHQUxFFHDAc8XeAO62mJAJxkQWnvvwxQ9rDTO3jnQFWP2rcwO9w+u
D/O6OksGBsTNldL+WorUNUx/J1A6o6dljusbojA708xuZLjSreTl7Ei31K3P35UtyceHNzXE4lK3
FLqVHwJ9dYbOd2hPHx4S3KdHMICTcTqyV5osFmLKdIQ6BvQunUgoz3jqNou5r6bBnNxAO2ABB4qB
6Y71aHryqaao7BCDd2Q7h7/auSm5mZKbjWs7A7piJ1V4JAP6NDRGzJXlhYEUQHsXOuzdZiCCHp2w
2KYfaRDHvoI/kVJlUQngRcDyJeFN+NUz3oxjqN1Chtwzw+tw8RFW42LdQfeXOnnzSikj9EmptqML
WXynTf+Eyesr+LPWA1ruIdkrJkfvujzpvRmPizhOU5lx/ixQocqnCeyQ7aV9HHKAmBdUcvrgHzdj
QiN4hDqg+ZQGBpFcT9eWlpA4ULFM2390bgfeFpK1j1oT69f4S6Quyu/XKlD47cus6f3++edmARXq
SGL/uVLXIkCwi9iWVmANNdv4UyexK8Ukid7bkEO2B8sxKlUeI8fgqESL9h2m0hrJhIdUyd16gxf9
cKORk/5ir0UvYYMZeUGUiHwoR13Vf8n0vMaC0Y0xXqUJaP3vY5Bi5zQCov7qIoU59JJJk8E0JLRx
7AgBH2OHbgHDuPYTnvnm6nQXSt8bclvAoRI1XqAhBJJ1CIDSYziFBKcdjFSLmXkHIwHIEtcQVzS5
5JNQ28eFtmV9zSAuGmOvwfJ5fIUDBXSLw1KPc4kKbsD1caIMjouMf9q5guomz3pube7dbO/Tp4DX
WsMdYCj0SIn//mdtz+xdqVqTCfXBdx+L3K3PC9uqpumuMEMqveENHE0DcsYtO+PwPs1mPpzRBbA7
Jo/sVfdV6fn7BSeSkK8WQ/8DeDT4CgivySDnfU+dn2utM8tEbUvpIq9t8HbHAmIrCrtnN6vVxAQ+
orXrWaeFdJQn1Mq1ktzD1WTmR7Z3oX4k5dnyXHESHm7TV3hghXvendief7Eie/507Czy5h1qF7DL
mqv1Aw5q/KRVZTiK3aa1/eWPH8kWt4sQW5JE8DR4sxl060fGfqpBsPRZNmQ3mFCbeRkar0aDUr/I
EACTqtrvEywZNTMZaAHmemoSVBgSAP07chLrbiUEJDZ6c5xbSdiUXxmJwOP+Ew7agQKDTfN0ddsz
DwDIAKbUe3ZN5hQQvgbrj0mEk5W34ZFUj8qhaurjsvOJ/DLUdlte69cAKaiN0At6L8VUxhl4I1Dx
XMVLRJotFav+URiZDnZGPwS+N/DXEP6j30nfE0yEvhj9eIe7FEOkKHP6cH/EuCO+FkXhGtLugMC9
1VNnh8H+PhoHBo0ZmOPirsgnGOnwFFIH5DrLmgONl0SQ6HUO7xrNXBj3T+DHGdUcJFYdEVuGEfol
S8pi3EmfOXyNuuPnuv4DjH5wQd3uVnjetFjkj0zFEadkjfTQvOtdzoHT1ijEc0r2ft/G0ldQIDMT
Dy8N81yuyQJXIGZHjp1XmPM4ymW2y9noYRYVEUwHe5ZEJEbtFYusEzLYcDcVmM+LesCj/JoP0fjc
4oxQcFicnHTQ0L4bVktJsaiTh+bQI7NzgalU9l/7Qvz2KdvSYEpLFotkW8ejyprci7rzrg3HNdai
2ihuf07Rn0G4HD8LHcgjoUt850JEPmMuz8JvdxvHB8wbBu1uxkXO0/R1UDSTex8M4hWVflzYad7X
8JJLi9qW4lHTJfhJvFXvbhSBqthKD7Ggypoe8u6JqXKWcWHRuLRBqlEOMVBpzFUxUL9WbY/HgTO9
PCvmA4xxAGlTbZkldPA4pWZQKcG+vR5btXqYu4K8HQpXuvXGrKA4Rq2W1w63COi4oxIVsaPv6zTo
sOF/cSl1LWsYCF+bikjYVxMuqU8AsZU5mSnMytwk0TqcEqdjy9SDc/uIPE8JJm4CB4XN/7e7tXWJ
vCZxO2XUemGg1QYLETqkLs+6RX0xEghnqJq2WWaso4JejwAWw3na50Cd5QLwQchOUE8N5hhTzwb0
8HFA4X7X8+VoI7+nI8qP+lHxsdbPeYG8bSqezLeKYhXSkbU25meOCKvtclywuUqURTOx6ihjYYDA
TV8zbmgbmHR3vfURUVcH5ASBINAuEhON3t84YK2srGoYE39ViiDylNxD8bjtwxjYdM0wQLrC9r4c
3+zWdCnsvD+pXEZA7Y80hMGUmLC9PaTUBiqx/rWBrN8F41k2CU2zZ+qWrGxwKciOGIZ/68DgOYJx
Tn9VNDX4/IOFeeqV4B0Rmxabwovv3VpS2BnfmdwlW89gl30FLfrue8Q8kq6NakIl3QEZOBuQYJZm
i/Yhl6+3d3xjSBGluJ0hZAvNJe42AKYqvr2dYK6Ugp7a4wa6qJywGtQNs/oK/LnymEUXV5KRvwrT
SH92W7mtAbAwuzqJI8uF1eyWobLCOKkkwjz0gpyyN4pBlUPID2aQHxHx+uMnI9c/NDsuQ79WAyCg
DpXUKOLqPm+skW8jJYuX7MqaPEMiovsiStRO4u/pka+rxoWRMsu9tvFLWD86b1/cGV12apKsqWzm
dN5bfJBn3HfDDoxmpNV3hijqrXoTCzfMqEhDxqWgWZf/K10UYFvD65rzfu3QklpFhK0V1IuLVuj9
8cM6Boz7wm64lU6hUDvUJWCo0GVG08S5VAT7+Axmiu5QItO+tzGCw5kQNsfwtGc3ToOlZf2OFJch
rjp3SIWf8cqXnkhTc4Sq8AjNcojIfwQKVdDckpzSMSZTJs8pWHcuJNeK51ws6OnhDAm8jgyoc4zR
MOtgD2ZcWeIYKHIN9JkNk9vcG1pRMkwBrFi99kLE6LV/UeznJHJhQmbMcTQeve/chGl4AWdeSi5q
9XmzcViWECOwTntsBxGDOdaweZwOTDMpeLMRIbhkZp/swCFmO/ww6lAX3dOtn7mYUTpHpfVP+frh
rKZ9M5rejCmoRHIjuYIDN7BVo+9EqN6MjEQ0FgwG5um77KVm7EtfDahS3cnGh2nhThP/qTuOBiNL
KzZMobXRoccQNZrdvCFIj+y8XiG0iwP0K/B2YQabluy1Vopwbvy56BImr2POzNBzOhM1aUn/UbCh
BzwXY4CKPaMelAJRZYSM+DDvlhHlzeefdXfT7DQJOUNYJKNe+JmudxYIEou1G0ZXFw9KI6QXoQI3
yywf6LW4V8+E5M1U0o13HF0TorKYerF4FPKIl304NXtWpqjbYQiCRyv2ugJcOz5Z0i/pSXxZpFaY
/S0XSM7ZPPVaBGu6t0Wd2bg+/js5ONDerzOtpEKV/Aw0HA5EuHljENEfDwYvBiTuSbE/XqKQnuWl
oPkedz92eTZr0EiBOVCzk2ZnU3Cof0hKdUIEfotDmzoj4VSM6APUhYceijN5D2ztFKV3JSroTvNr
6P9vVo0dkwL+ysUjQlMI2eX5eiox/MUvrhnjfxnBV3qtw98mPwJQjq8GX+GzcigHjHrRKJXRvLaB
9NRUKg5EPtlliLzfI64g/KBdaY723/BFSP6KhrIxb/pGtkj/fdrveqnBLo/F4c5y3PcnXmzEnZz1
lOuQJQ8t9zrDFiocfu20dM9uHK5d74Q3v4QsNzfps6VeUWS1mdfJEYLctqrpNKYqBe4GlZ0OltKW
3T3ysgEQgPb7/7hUpD7cf2YZX9vKBW/xhum9UEjOWk4/oniC5fHOWfv6w2zJC8NJugSdWsXDXdP1
QgutqOs1TU+Ha8FlcLKxGJ6plu4TT7rKA43JBxyvFpObhkYqOtnQczpmvqyQYWv+JXlVsrvTZjP8
3+sWfFAXY2W7fxjJQ/rMQJ2DmvgIbBX6LCHCrUHSnTWM9Gg/qhv6e2+ERqwGOBfZ2MZ4ev+bhUW7
F0WXoXcvhRfa+cgTyALAxTAYRVbkeRQn4Oolj4LOEsVSoDBoia5yd3SeAm93La1mock/izGZFZXQ
2NruLUPNqsAlwhKJqVhbmoVrCxWTvGkOoL1N1C1OVumfqAeGI2RO6f0fPgnJ4KtcAEDK7QF7k75z
1jEVYouDJ29pNcKi/AcNrcCvTOvKAomPGTmRlgbdYsrM3+vDIkyCT28R0Bsub1uCK9XfCR+18XXh
E1BCaBZGFxfpvTs7cei5NGo5HAZOjreQZ7L3NUY1SoYYIvYKngIvDiB8G6dbbcafqEG23kafRVIN
gh9PAtql2GQQjFoCWioOhBorwo+m4cGaqdtoQiVJGmMnPkF5Bgpxb/ZBMoCvI4Tl4zw9PyEEn2cb
/VyjB52NNpn5iqVLSYLFLHNluq1igHeCRbK7xHfqVD5R33jJbWnH7tFlNX3Xz+d1tgc0RA57xH8f
sV94vTwx51AUS+2cBMVzyXqOCR4aAswDAmMpkFEFCl7zSDZe6bBZ1PNMxrtXGl3DQEW3KhSOOtDA
1KozeMHCARx9nCinGY86R6Pj5CIRUcI+xqfpod8SrUfyvwn0BR+N14/48oGifNmyNQ5IT7Oz8Dmj
E7wEkyl+gI2orPoiw5bE1HBjac2kK7mTGxvTjHPrgmjgMBZ+K3Er2YkxpDYNM3VqI+xZxkCJkoDU
MDgMrv6GiCuCljcfyqlRYLhcDmxH3P1sSObBg3qMVLsitlwd5Vr4D4fccj1ElsHcH0dcylnjNYcA
bZ1E1IXAzUUaOWr/3Uddr1T0MSClF4FMHUsrWAL9nvioZVtVLLPqyAUjHFz9IpYjNHdiG1uhJe+/
WmJh+Bkc5wELBNdfg9B6AtQ9D6ylpTHdliRkLNXHKlKqBpzf3xntEfA02sPhbvqaOrNbsTSdTB2h
YZQ2G87wflL64MyAn0xSb9LZrtbe5Duk08KaeLAeXDZ4x3uBsRveUPtbt0psbUmja3Zugxb12d5D
urs9G+xa8ND4DkJN9GFUNzqNSLb4NctlMre+NqVh/Xa+CIrp+YeFv9zprYnV2xRJKulmU7R/cJld
JqiTGBgWeZnVkxWI7CI8G6krPiLJe2u8N67an9MwC59t3IDIs6GAGZVJCwlDL6202qfgc6EaCDT8
XJGbvz6j9Aqu2QurKj6Qd9hL6m0zK0bwfGZ6sVX861tAo2G/aGhbT2TMoct9sdOZirK6o2Lvm3By
vdP2SOor9Zky+GomazL9E9pFay5+9GSRdeODC11yarueRQtdUZha9WsNzv+EFOV7tjKktJC3X6u8
FFQmFNX/mure1PKLDR+tvjNIQtHdX0Y8dlX4Of/DmSp5k2xNdItKQA7q9k6YyW896dTsx9bKvkoE
Dz02zTc8QXLzBxbzx0GBjojuO0NVgkKYv/59NU//nk1JMGfHj6ZI/6dFLhkaAbdMAaicbrhguUGx
virsApjKbK/xK5w5/Et48+PAGgf0wmkmEB6kL1v7xD0BU0rrX3PFM1mHPgPoMygV5Q1QkmnnnRuo
elv9C3vnI1NELPn5XOBQMxlCn3hVUPfRvDexwiZ2Tx8F1KfOMmFTv2rHocgREpmmVywwcdL8nqMT
d3/KMbaOqlvMZC4RvBs8H6DJtq/UDGIu9mKdBXmhwZykxnAus0qoqZAR9c8Q2mPmXAKJKTx0/2hf
aWgkQ6plVlXJNlnhb3o7TUF5B6dj2DlDMEUkILH3QwKmrzykn7Tzt9Xvo7TTF0LPVtgJMqMdmVak
WtTD7nKOK4sO8yFLgCt8mKXobyk1PfHilRsav+BUPrccgW2P7xqdsNnFAAPprLQxXqgNKc9fdXEd
l0tLQB5AkQGVQXfxII//KN7gZRzjXVZXE61hx8ESsO/mJ4vJpLzFzqOUP4Zk499bGvI1h8MtGFUT
OVceTahuD7tLT1h2huJXd9UpOTOSqOU3eUJnYsvosT/fnIZznV7OvWyE+GfalQIAZe4OSURZuoQG
TZJWie00ppqNokx3pS70pYzcP+awAg8FXWKTXlT0j4UOV9O+AObE/NXtuSPKBwy9Nouuoy7IyX44
Nv7XsEiBGESSmJP8trHoLIhjRgXNmJWWbHYCgmOH2hZuktQr8fN9SfvDh/Yha6qeLmjq1KP+EZp1
8g5NlyKiCMxmiJ1w2aYSLJ/J73tCb8qm3NyGBcc1ubHGX6u0bL4+ictllCzIHAEyDf26gMbC4xbQ
xp/ZER5VeTttL3hBKOgWPu1aBXts/WhOQuHiO4aBE/Xnu96pKwLuQ2aeWT40CkzFJiMG2VBkU+l0
GKWUuLfu3bNd3B1OTcj7z9Ou5UWD3SzXjV+EYcuZAvc+HgOraDu8CvdEQ2+bBRYAa63hjKBPS1Tm
gUAcmUDhHQ7nMqLlQau1EgyxyvUDv/BCObPplymajlL9TxueCsthVBP8fY4DZC71Xpluo/Rjaw2W
yyB1j8Yx6BUmh3D7A1lPT1Ndrauy6jgbBLJxkCBbgmJMOXg9BOTcA9KoubzXd9Bxj9vJWFK+TG90
Hl+ef4yYRftOIQLcME1fS7kagEfMXks8NTTdstC51VyR362+GnEhhMWECx+IvWvTiDmZXJyv6uWU
EnTK+IFU7kwdGdteBAB6RKpMGG8kzG0387KP5NU2RAISS/tgLvOKOOYyDpw244cPz1e6rMBmVQjD
swUZd9YSMTGknvyGz2+LaXBFkZepzyarw+Cahm+5y/BVzvfaOpZPUY0nR+z7oBGgPcyQdM4gOQQj
brsIrVNvL1PLE53STjpbFzm0t4ugflblRM9ujmjn2fG12v6K7rAVNTd+9SRpRWr/nIO7e1nDPfDa
1Ip8sBiDyp6Z8wnrgff3XilXTbd30ER/HYYWl+sIlkn+UttH80ITeA9zxztthbjWp0URq4II6JnZ
FHpV/8Hp4EhOxCZPz67h9JqO+Fd198QV/1YfQaMxgaEOSXeupT+gDllpMVFPLwy7D52gxvPceAmF
DyVoW0vtA3v6avwmA/v/D2zJdBA8aNalO0x6Vt0VBvCzhV1PFgZd1h8xprPRm5XoVEE9gFJkOpI+
BYZ12xNRscf6M0+aAmEo/+eS/stltPXUDPLuVVl07U0fc7hbvlXUbzfqPMUayZaGbXHOtwRuGg9W
x9iy6sHMZAmmD39IS8496TsNmiKIanbG4n7LDr/1FDPfcD8QwBBoxs4/2HBf6uS8c5qmiyah3SIo
df58h0AaxQyccVIKDUCNKuRmbL130t9NFI+WQH9T8aS4RzRteBh4awuAx8o3EJ5nin/gv5hIctms
+qtoaN5r7KzaNGB/ufzB6tdooDLlm0htz53FJTh5yYeCdR/0eKt2pZ/HZM4JuCIyjo4neo3zzV4b
zF7JO2OManfi+45pEpoSvEWeQmtfFZ8rbqm26I5pIXdLHTmlIwKAKZbJ8sTp2ldzg94gBNyaaSD8
sB9ppqCLIfrOCS+eleU9w9EI4rZE0D13WKvKWWl/ardZ8gvzgMJ6OsPTXhz/89TJFvqjWXbnUtLK
k1z7jekMiEuRdvyLyq0GT9db332ZlvaITp5S2x2fesntUaP4HjT7olsg8Wmd9NxfT6IqFW+bvOgQ
B77BuuxUZ6mcnZmXuOtO0DUeD+0Pl88J3smLGz2kUHkTzyn077HTABdpOl5lVkrt2FYOgQ0IwUrY
ntZ3bu93iU6gmHga+wyoi0MG3U19TwBKVH8oxbSz1l3zSzIEOMppmHSXbjuP0R6OGAhYsMpUazpy
ZmRgWdTicocnWo9ibWTAHxpviCv5GOGGCUQ8RdH/ju/EiqQP2PMr9TiASJrIVNbaVj1pofU0d/7S
mfMyn1O3VznsbKiLuMGnHcqpmUtAwK3lXxDGVbGiRI/MWlyfikt9wquKIg33fEJSvKk76/PHg4/p
SekHUia0Hco+HjhNsLi0QhQoelHd897HqZ0VYQgV0o9pNs+Ld+aQ+Atd3FJyVI8X19vVxJoYKB1J
vBMXBkgRdzlCJjlqBudWQ/+DDxADnt+LMVZPac4CSy7DByHZDG5xvACVSi7AUO7GtrrSm6gjbzxu
QUTTL0eehSspfOkYzX4KFh5RDHYN8dk3VMG4ZlsHF+OTPkoXnJkJSydiOyKaizAv4ygv1VfvzjoL
PKN1kuTKbniOrSwixlSTnR7WxMei7jUK0pmj2sO0j9DYIsx+hh7C3AsdSc2lcwUJGMbEqYEUeRQu
fDMuAgpzR+d/6chqE9Hwrq9vpfBz0b9OrlNef/sCgyPts04Ke9/5REkkRic5/pu1jxztP1ht+Q7h
t5boaFdccDnmuT5iKWk0BGh/6s+xZzA9t0RN3A/+s8ZvkAAGH//N3gcrNqndf6+E1SH7hphHY3VF
oDmDJAk7p02bG/wv0djPu40OlnYtYgUH5AtrIDTrXYvwgdc1pT3PMOc9IU93593S8JJMwddmZjsI
xJGrhpcao2EhH5fBrPDd9Gk5bwQTdKGmatm918il5YwIhBcXa/bK5QvQEdQN13008XI+bBcQSpXe
y2GOjD4wZoHF//IzBWV9VOFnCWvjjjaJGeZUXhgvbyZhdXgdxPFn+ztuC52keYDdFR3CaXwvTUOH
NpgH3iZ0cIHPVxGxNH8qSRnlyGIf/hCl4LpUZeZAEERvF0TitTxAJVz4nFy23l1OOB6pQfrPlFw7
Q3WUWeFwTDrbzeL/iAIHAYqaPT+1PqS9jCg9myoYiQiis46VWKztooWhjPHQqHePWBBIGdSl3x4C
N00OpIBj44JeB+8pMqfWj9L4LXgJVUT7x2PoFVgE53JKgc9RLh4Ei/g0pKsvaxo7Jo3sg0MiqRY9
uRTJ58MIaODgUwPJJiuMHu/N558Xsyqzhl0a7oKGusJkiYUDrxzQd+uU4FgsHB7ORxxlMrTU5SJz
42DR9U6FFgKjXacY377v8Mv7yewitdEbRL41Gf39tn1JTNCQuzkO66AQJ4XpTDLUrnIngroIAcIc
YsrA964F9zDkgriKfb6Wq3zo46Hlk9Tz7zEYcwEBTgaLeB9UC4/5KZtQaQhmWPoTWdYUCWSszjLh
C5VvXNq9aSsELP68SRDFIsJsRIYVTbfdRoQj4qGTxWzcDyKS12wi5Ze2SLuUl6b3qc+ImrdbHjH5
V3k1eMjkpTwQPKfUUg26bfQn+7CsibDKhuT6o3zRq1sgtPuVOFZdNWHpq3n9Gr82P+GkGHJ0G8KE
Bdssg/v+QrSh8TMSsAN7BRv+zEAFtxy/JL/rVZM+cCqYjZztMWgKnn7lmZFolUezjUvvaOeS/ifa
7M3ZHFQwBnV3/u0HEWJJTdLLLE6IaGp91AAAEjvhmphVq5YNx+6TToC/hYrErOf2EnAUSnSJuUWw
msPZ5UYgqygu44Px5Jvo5/DkbYgsN6kABjvKCtVyelXp8XaGkafPBdaRUuO0hnZ+zdnqtG2/ijj5
wiQEB7U0qfid0eBgGkH9nN8Q0t1tWtpbQGqzPIZlJlviSOCrBHPbPNBQ8RolpJe0PALcAAk0AbfG
lDwJ0M8MKCx5nYmXQqbO2ghf8yF0dI8eFpXxE5L7SSPjTqdKo3NsIzZrrmq7QQhhpKf69OknjfPJ
jiQ33irR/nfAcHykbyKDUdiiQRMoYdycbSh0Nt9ypxMNceIPRDDl5F6wmaukdd8UEsECKJCWBEOR
iXDzNLl/2mCJN9T9rbuCOYxcwggoys1en73qktvad8mYuKqjEmbcfFIbiCa1Gs9w4CKCmtndUsks
ZgWvkbJcqVIZXRpy7B8eHL77NmsC/EIo12kKI13u9mU6EGLytO0V7KMcf/VHBhoXet//U9mafeQh
cKhgG7TrUkFAjQ/nN+l89mMGr8LlpQoyOysnjIJQHJog0O+j9nvvYUXK4LcqCH8Ndw8rydoJsKFl
c1AjQ0qDWF0RWAHuiBbvWUE/207C+PeXILBYYCu42IhWIxVbzlazcex+1JYovzMVZIn5z4bRAjHV
IdSGqArn+RrGqNFqbscEUKjj+IBL98CcMlxxgJTcn/gydelGYkq9Ec79AIjSS/wHAahRmxr/kzwC
ksn8YQ9Y12yrY7+KUXdry70un3EKtYdu8oRUf6jx7S2X7avJVEyHHz7S+YnDRWX4jRBn0/JB3gVd
z2hl8Kby0zJ1P9unhi1in2P2JQnLhE52xZblPj1Mk9QCQcuc6xt+XqruAXYX/wSbR6/Fh/NfbG23
CyqHUpvXFlk/+K/8Lx1wTxaHyw7y7rS9R7b4bdWPNixtIYNtIe3wXm19fZbkFsIzZNXCRibnuBUI
4IjpjXGa+l9xuqONYmmoK/DULnXnOnV/0j5U1Hvv2dca84Pt4K3pUclKwZrVAKjxHeStLvUouYaW
FhY4yJr5AW7FaAO3944nFPL9fjVi/+Hcz8wRGDUbkRkUiACJKSK2J0ob97iUcWBV5n+F6yG5hgAx
wmLT37c/kb5xrhARdncABJFGAiviumXVKH6WUlKOOJ86+CU0Ktf+ivmyCTDbL6r0VOUc/5D6SpV8
E7rRUkpYeldu8Mjl+2BAINr/fRqK2XAiCkxgrJvq/t9cnPv4Ld4+VSpDEGraQb88Y77K6hwzcv3E
goH3svdouAkHTYODeRjnfQlzXQGTo/MhTyyZJFXgl7oie4rctcIo62kILgFtVB1u8gDAT+k66HSj
iQplnY26jVvkyPe+LCJcr1kEqczJKf/iF12R53NjCgvV06D92w5f8kwAWEu3KjM9+KQ3q2bWhqdJ
67pJx6+SyeZqrozXvzdQsfTXf2NtYrpFZ81vkf4i/8aJLwjd9vImhAsJVdw6kQieGCVaaZeXsPqj
TKuqHbXqtE4BsbUuIkX40Eh5J9IwUpetCN7c2G7GPWIp3v8ncxI4wL2fw107eezznJUfU0Gt9j2v
i3TDpsmSMQMyTh7qUL0WBOz4dcaxO1ucbXHEZBiCUWCMKbto67V9X5g2msAOLG/xGrtSYxYl5oAs
x7Xc+0a3087o+D1jAzvm9D9EdxPqCqpWoxgcEqDACgqVphw8gbEhHFd8dRcJXj4WctGbH4QM9Jk2
/tQl66j1x05eQDb2e/6Lv9Hnpev77EP8ZCS682T95KV7h0mcwIuq9oVgudzDsfX/JQygphzzZHM9
RDeKtSCFnG3SYv56QbmoidJ+2d7PMMRpRBBXtIlM7C8n5PT/qXe6DaNsF4wGvtps4SetCymDGps4
3V9XvuAr8gTGQ1b0/pLDZWBtZZVN/KzpYyPA0FXRxKVI9l694YqjllN/EVUNiUYr/GVWF+M9avuE
qZsNh5h1Wmy/VdZnZqyxVmYRe0++dNkHn2haR7sNBTD5sRmwHS+rxfXcsyPovtfTL6InyknPF0vV
7N4BCoq0JKBasBIs4j1+tFuIvd0kCfqA4Wkfqzhr2h1aHxhzXAcXgXNnv+2nxQyKi1zdjzvQ37Jj
Ub+thtk6zUOmuFgxa2VMskQGeTi0whPMv+WixE1SJcVqs7IEbzh+ZobVr14NRqJYNeZOAQHyP8vI
iZ15wpFdJie3iTKkt8ByXrhzHaZkEAuv+wF39JcFGOwZFi0wKV69ZMEnGAk+d/cXRvuLY+JKErWf
vmy+o9s1PUQLaK2aVfwZruUUHKVKuCmR9BxbjqQmiMjWnVSl1oDEHCQSzux8/tRD55TBMFpTcSuW
iJ/qwHBq58ZkGwN2QIVBtluCXM76axmZeBtLM8kqU4MsTErY1dHQoirX1tG6aXvt2NyVR8WtkFw4
uhkJlYg/+QWuYUCqG87H0S1+8KCWyrljJJHAIg4LbMBqthF/w4VL2YEEkLe6EPdCeJICb9gWZ2Ka
2P9wayBuohYA/4bZakDZfMBH/+ZKs2+14R6cO1/dIFLEyDvMMZ6M99HOhOft/LgZzvGbmdkNo+wJ
ueydr5Bjmd/kHykvUksYecLAvs1TMbLIdeStceIJMwxDqmYSuHzi9aUouJEPblH25t8hHio5YWgP
wCToLg1rvE2n07yUZJggv2bw08zJtsIsz5Yi9eq7crLenwWSMOJgiNZ7ZTIVAxa6RXuhRxdZ05m3
W3RFWfkNewrn4gOa7QjYvIQg1xx4ucBrzsVLNzaptrKQKOmNRPl1tvQIRemgN7zh9pvT0pLcxjz7
d1bn/kWeEQ73bRtqo+nnyHk7PtJiRHmMqLaj+3Mvk3jlWmfVs1pQb55XVCfVs7k8l62l5cqcuogB
6DkFj1XvLFDzhzLBsQJRA7Rd1NRPk4OwWwjhVDVrPynU+qXFd57AzO92GqlBfhUOcbOEqU44i5XO
nsv7+rFXo3VG5PncpaZfxKTX7qzDFmw7zeygU/w8j13mdxtYSBqmaFq4iIaquE6frDb1aHlwjP+d
sPr3YVYM6Zrv1WmGR4Jz1OxphiMM4GpBm4B/2Szx6MK4Mb6p8sKnVzvVaEWwNLJmu5E9e1V+Pd7H
pXKD9T+C6L/pvcANwttQq8hwTPp5PtXwsYZgMkpfRgGxlpSi/f2zOiKtPlD2tQm6pByM+0g4rdiJ
PYpA07wQT3K+UZiBHd4kX9tT0Y0vfKSicDcRzIJPp1IvrTuS4Q48QIlNEob27I35YdEvIZ0g1tWY
LgljGxcNQjXxzDPqzrPZl4jOuUy/wvM5G2FfJt+ngN9PPbwkYT8UDoAN2JGxFxEXu54my9t7sbGE
wApJGGqIcOD5/gaH39aCYMH7DXcvcfppA+PgqZjhYOsgkjif+PvBO3IXbD/g+sLmwZU+UN1TUHJg
NrQcLog16tK4vUalgXpipfAkx7U+ZIj82OlKTB+ntBXG3k9TKpYDQA3S9ucVJ0G3HWkh8vcyzvJ1
I2mmEXf49UO0M1LZJ59heLkVI0Z5p2KgA6AO7wbWvTgN4EsiKtI/AV8SKHKPkmKm/tre6KqRU+W+
TJvuLWEKJg1LGhPIUfXp+8Ni/S02V1Jmp3t5Vgmj/FmIf3WGKtcNm33sk8WoTw4dZwFsc63DnnqZ
p17YYQDFXin7OegabjEIrr5VbVP2theN12BuKKz17wi2/9G7viYVslvYvrYAuuqGpqhT3traWTaX
OrXGrezh+DdN/1dB1sZ4bn3yv/y4x/aBtprrmlUUvUFEV1iXAdtCAX8dXALY1LFB9qs2uovi0XAi
j2nnQPmBSI/cP+SqQviVSwa6g6MJ7BmsPpwuCTW3YiiVWfljeT0Fa00YQLH8sTptElbRt9lffVjV
q7FEbA6+TBE1gmRQQ9yX8kgcNDjv5K7af2ToRsRURj9VOj83zaoESZ0imAxEvNVQKezRwW1XKw4w
PlfXPw3ELz6Rj2/kqJaXFQOj70cr4HykfnjC/eoqjqjXFzGhJA/syS0Rakt69uBPfXBJAdfahS2/
WZvLeLk5fw8+A8e+7+W1SVYjJarf6cuzrm1U7diq4wFmeiHtmQeCy80ZRKrUygwORF0hXn0GWDei
Fh7zDS7vjpB/ks/kKCifiZA7jeSZ8MDaQ0jhT0Doxc1S6NXMAv71ERAbPJcVgNRrnsa6EZpb1v81
Ld0QG5G//iULLgErVU6s7e+P/PRNIvwNzpxDETEyl/MFztKR47WyKhAtbSy6Gli4+eNTQHQi897P
DSG3IMzF1GOw5QKqn/I6IwILgS3uGrUx7AQyPwe5/njByFDKK93bQXy0Vr6hA8hYphIadkFQ0kjl
ob/waZgGpsplRuP3++NIum5zWKg3llGKyOcQ2qrRcBdoMuiXaD3ALP+JSipp+o+gfAx6hnt3UKtz
YgPENFEEmVjcVfSIJu/Ek2GgL37bTF5wz1m0EESfLyNGdC3ojQUNHkHl8yrIa67w8gO6FTjawIoW
t3JXyIvQdFNppY8mfmHcvP1Dcz4+RRlS+8N61CFt83HWeDnmFCKyIkL8Dk8ciDHxMg4JTCgzkHsn
09cVeQ4o0KTxv3qWzASX8H/9TDuN5Peg6jgVfQFguHU8FTSvhUnCS5sMrShrc843I0s3x9p2d9V6
Um0XclvZBLXiwAFesi6vi7OGvgEtRfq5U5jzJjOVH9YatfqlOsDXPdzf0nN956UdSZ39bj68C3Jj
yGvmLjmie2q91l9gfXf3Uq0KQW04wQQ8an/rVUz9FAjIRg+F0M1xDVVkULQOKKs/V0GaJduIsOhD
UEi6o0s9FpBi9qsdUeXg7Mew4OSuN2rWWTq1PbMrbIUiVz7SGuuYSAxHCUR7SG2My+HJiwi2tgy+
RHKmczq2nWnHtpVTcFGfsDJFZlznZxV0yz8JdeOfO7Qw1RTW/KdjR6Io7v0AuWOiPjioj7fchlhn
F4sCxxmnzHJlfkYC+oVZAouBtES18+/AmvfilDURdYpoz01eyqldsEm+0GOl2QjuKoJyqHAIPlfh
Exu6wcJ45g/5K+xLdF/Nyi+cgdPFN5ITZuGbVn7azk2bP2EsP0bMm3F4G2N5mRa3GvdLCzBY0i4W
2jZYwMngdIuEb9LKWGUNBAG15fpaCCSHt6OM5uP/Yxg4vVVq6UI1eELhhIzRFPkvGOpWSRVcL9vZ
pU67PG1Z5BKBeiSSXtJnbnUPzzyjtosVFhXKmEASzPKnj0/aiwLMp/DshNHQGu5NLB5bMd9DGiFA
JDEKYBeVAOdNxY0jEVEW/LMOZ6SBU6aHgRXLKkI+VuuxiEQILsOhXBKxTXnNsUkXe7xoNSN/S9JU
7QhckDrUaWQy31p8EXIsZhKBEQLX7MPCHY7/GbhF1ZxV8VpR7fJ72JkGJDCOwRNbqbfsuoEaOtdt
JEuyNgq4FbMMfLTOYY7U2I8YUiboCKQHNmGxsZFVXq76692/OBGi4urX8ZzcUbZY/7jnS+3fgFoA
abzgp01NoBd9PsrIxUoh/tJ2Alg9Fd9OnhGBn7MHZFcej5oJxTriPSnBLtv5i0skrvWSoezcpKPV
i2GgtU0UOpkoycd83lWFGbpKmaVuFqtqpnYmD2k47WJhhf3L46ZPgd0nAMiB0m0o0QlgZg7hR6lc
b8mQj8uYqCB9Far55H8oA45KnilqYMogogD4Ipa1eJDcynlYuTMrlW2FKISqVsKOxtlNi8VE4K9B
yYV88AKoKhoWq2U0XwWWdpGJCBM2Bk1DHmALYvONWAIUW978/x4P7OxrKp5KK9l04ezzVBuRdVgv
zDmIdQ8YjxzJMbRafsBauin8kKTOWkCJJxdl3FQy32EVRT+RicDw9aqYpodkto11U2HbYT2eNavk
Cj5iwIOU48nsnfunlG9J01hER1equQWeBbatJUnibvSWuvnvcAnKS84hw2nGEuM/QU9dk4kYIBtx
ul12xxNtb6bwH8r5dbLuGOPVxaGQgCFV2Ng2nmlKdSriFpZWvlTTDPPIZRAWszROv5dDVC6cHeRb
+fghuoofUnVSUkner85MM12y9zA+Zpo7Xqfq+xT+gRJCxWTH61DJzWxTZ5yQ2xqkuHCpr7NAM479
XH81LJtvUWPNx1kDlMFRslW7O5/Ucyvc73JH0GM/dmZFB+KHvqdKF7BLUxqw2yD+nXEaxqz536r8
O0CF0PbmEdAVoG7ccBWdWYofqmojFwh7x4Jm7G1EElWEejklJaPS0kCRz1EiUCyP/D/g7jMNrAPH
XWM6AEGlbuk8aIr7rj5yRf7EXVxvDDkUrD9DmtVEoLR5ycVSJ1/dfKODEPj9YrgrI89redzXJqi6
bg0GlCiS/ajNEw73uGDhv7Yz/+PaM6PnGxBieAbwhMDdPRngh3mgdMKVge6cEl4bbE8Pznokb95J
8K9QRV+lmEgvRRe0H1tM9nqEfNcnwcPFRL0U7OWiLloEYGFUpkzzWziDOdbz5NRn8QFAgrEVUGlO
8Z08BYh8gVbH5JQI27SgbPn6+b7tYcVufxcNDdUF4vOmg0AgE+tw2pJqm52VCs2AixM0Mms0OfR1
PH0n037RixUiLH2Tl+aOWXy8frA8JF2+5kALQ0X57HFH4W+0iVtC0KjK49lOZo7rsPzkkw5Veob6
BbDtVhm/ysBWDIqDStm89anV71LltDrKM9SuMYLN3PgSNUR+Na36WldhpZ8FM0cU+Shx7ldw6/AE
X58pTmTyNFpByAnHObClmYeCqbPdabYytnKbyYVK29PWWDU4ZeVduze7kNbql/gVzfUt0XmUWtBW
y1C6vqAZMtR7qbbPkLlIYJ+dt5Tbpxm13/dYkFI0ZH4d/H0mn7EhAdtIoPzwsrQEfqK2dMpwgZgR
cIkz8P/lXWoQfcYZPcZ9Dc5Tpl3S6ivuBJsodzSJ2BuPoARi+ImGHR1NSs+40AFzgdJ0LPy7zWxd
UlZHkS2cBixMfHEefLpMJLbMtl7JaK+INFVorVcjOJumZP7k1Aj+8y1iXNKeM8bK2M+yjbrKI4ON
kjJwROXqxbASxZEdP0nyee5vymAxrFybtBQAqmnbCKIuQQ6DfGsvTDDZTWnZD0BOTxWw4W9dvwTS
ypftKO05lr7UsRqhlcFSO0UtIERZZ/bSetI4qS/W0yBBfaUm6uWd2IFkT0XD/MvriLMKLj7faixb
tzdAF2xEBqiYW9vbinjscYLIaIzgTBCOEYe4kET5Z0CcPoLN1frMaGPCZowCpNBy7SqSFLMOBDtX
dpwxcE2sLIsfxKyb5yq23ELvoAjWJ4zJcLhTd1+bgaCQh4SPXeEcIuKTbxb+eASVrII56BjWA9/x
8Cd7Q/b8BrSrmvA5y7TOkRb5mZIpQ0hLus0GSdWQcPMTHCAr5TnQbQx3onnONymKJdxvOqjVdgQ2
AOg7UnmpMJJCH9iXsFrq3vx5nOrqZgyzs0kp+iDSYP0gBRLg93w6lYqGGyzGjHMMH5sSu4zIMNbR
fx5sm+peTwnEidWiEijCyAA3fG6etSvEERUhJ9H2/R6HituEPLOdLAIWULcOPfT8B6OJ+9lmmawh
VmNh3Jz2sdiPwhGzLi+cI4qQs7GILpXDzBcC4BO3ynFvjxI3PKQTrO1z+ZyOCpakWacNAr9Bzz06
Ml/kd25WflUIjJ4/YPMGjNt9RqDRhw2WCgFx9CYvZWghqutN/44kZeFlns1of+NcYL+UERgQLoeL
BPY3Ia1Kq1qo2qnBo5fsr2dXF1BI6+X8EC0DVgeChGwmRM40Aw1P1EoBQ1HZSPk3ZgedC4xE92Ek
SJX+JKXbWw9FuV4HD1ztPBpnwGF2hmT/g1/K6+gUQWYhMIV63JctEXiQ0ZKsSRVC6p/0dp9+zquP
7fXx2zNdKalRv9XrBUwjOJIYbOLPk1yWdi/WsdKiRRkzBkEbgYfmB5A+5iSFEBeempYV7JWFnEmR
Ebn7H1EgIcng/jFPQbPCwVDN9atBi6aKhfXs+ArUnajeYck+tL73vW4U7BidIgE79ODrOIrrEww+
9edv7wyND9vwi2hZjQt3AlwSEGGhXxtykoWe5KOP4+iHcf9bQ3gtEEt5yJA8rKxFcxhFDiDe18f2
pMRa9+XJL4SVKm6PX0ygtj6Sif+zdG2VAH3xjEh9aAUzQuLw/G++mI1V7Sz5TrTGLtpjXIbQ14SY
LNALx899OBPa/gpXja92ACo79mzmNtZQasMUBNvFAYmRYgyR+M0UwACwRQNno3D2RhPTq62OFyWQ
LoftI2OIK3hPwYD6eVyO9O76+EXvWzzf1958pLV0p/mepnxftI7+TO5xGZelhSpUMewr5SN3FrXY
mOtKHfwnysIOdv+1y9BnbzQIcBDaFr7fq/d/zTL26ck4rz2t6X09ngC4sE+Jb6crEWwDMuo2OcY8
C4O/bYCViWWhS+LL1SDrJc4Aswbs7hIetjO9HaWjnCJ0TnFUBl92x6rhZVc7gqA71n2Ie3aLFyn3
FqvEoe4mUjGIVDD7Tvl+gYcfdWYM9LFzaHpw19E7SqQrpfIY305vRPwewocnel0JtSaBSvPjjp/E
khb1Cn3aXmkppkrrBhPjjjxhqBuySh7kQPrcNuxQEP0Remy5YgrvrLf6pVrTmjHMr3uNyOzthYTt
363larQwkr0M9HTNSggP4yfI+58LwMk+6E9eZilde7p9t+T9C6q3NK3gRVHH5z8mDOLPHdGyipUq
6crA8t6pgnGwiG3DK7TxcNFjZ3rW0cIwfpW6MDyFmYTZq3ul06jnZmyUN0YC7cmrc9tvgprWeXS3
lAO+XqSFQvQA3h/G+A/T8Y4djrs9XWVsTQq6OfqepTHIv8OCXWYdRNFLZ7UlRSWIXd68tHiskxMt
MsTzYCb3LkfbOj1sIGhggCKzU6oBa+Wy5H/sVXNpk3iSmOmHAcvsmZgYVZ89QU7OqiGy6+r1OtMS
o3XNd/HV105ovzkK5e2+NHMydUvx08arjQA3J792W1yUvC/DWbYHCsaM39gCulX8zKjMuwC6WLrZ
KdpXOlZfWeLpDoR3efgVP46oA+P/m3tdu3ksuYsZzmg/mqPI7LdPIn7W4OZgxW/znKakc6I/O/PO
j1B0eveUsXr/DjYHq9pZ0duvFAqRWicNC/2tIDsQE8cIGGCRZfWxQ7VvR+JU7p81HAJm7s1PRffX
KPkydguyDl/5w4fHnhzC07oyAGdSLNalYzuEb/CmXh7kzf0B7ba/MYXwIvb97x6zD2JKJSCmHRBn
X9U48VN5h9Z3dj+W3lvpu350LgGCKXJAC79rv0z3DY/ayDtL7asUng5qJlioJ7IY8h9Jjo/DW2sJ
c0pRbBAYSz2gI6aBLyTe3XfyoQ3Bx9kxxd1M8dH5fydk2ZfLAtG9COQhIEwX5vn6bAnMaHHDiqQ1
Wp2OIqNW/J2+KyooD0a2VFnd0LLuagv3UptLkMIMFRG45uPnaVRPliz6P667fJeke+AN3JrZHuhp
Ol1XX26xGO0efKxQff3iSvSOh19DJ54Hc3A7gUOOOqkH6J6ePpayaDuKbm5WL8BNyUMgWvwmijgi
b6vb1lUggKrqiZc5GkqgWmknKxDuqq3TsVBdX0SDwt6qntm2/kGueb7WTnJZxo4KuVYYG9+xaEz0
JZ2/zMUcBlGukKsJkS8XI+8T2Wv3d6GwPidyyZnyN9dkEOo64S9x33UrhG7cObHJnmn20MJ/Fvii
MLctC1Pb2XM6FYfC8Ym1knLauBcGHKp+1IIg+xtB2PgNXosfs5GQWmEYJfwvHeWH8tl/pSyndk0k
PpZhbCLzFvzPRv1MHJhKOEfq3ufS0bHorINEqfS6Okm5MCR8/KgMiDsuyaRCSvPHIatJXiys2o06
MfcUAUrNXDlUOGEgaU0PrWhMuqPHSh243l4e4a4WIHkVBjWajh9VYwmVVJkxEEtiH0A9jE5oJ9/g
vTgJMTU9CS1mhXxgitfpRVqPoCicESq6WuYk8sB2mvpy7ckWEl2Q2MHT/69XgUBw6A2dww/ouYUP
/izkKt8HSoCGx2P/ru7XPEEBx6rAGpIe6JBj1k3D+pjSyJ+Sv+weWqAtXmMKfJwoogQ/WvQ++NdZ
oUkeCS7D/CXPxWj2coXbBT+52R6qzMXI6d/BGynQr6c6kvThzWSeICzuYq5RyYzXHa0Ol0O4HK/6
cIQCzr5kHXqtDdEK0oHmNXjVyIlcs8Ub4Vs/0wBm+ItHP+zwYEH906Q2Hcjhejo7LNqgWPTp1gVc
cg9YGhGVOky4OROZNLyHNfhnKchSHGRiczeYrRPrtHv5ECKdnr6qkQGlGoDHreTK6byThHhcg0Cj
/3m9rmqwg1Rk/v/dpTTFpJJnZ+s2I3J2ZR+QJXD4cArldBnHNuoA3CNi5at8PY7oH81cu7dDqkME
YpDyGW5AhnD2XrK5IHhb/DUE0Xw6K94aiARE64yZ27cLQrKEpGY0nwm4LmKgitQK1zfCmyPm5vq1
2v0KZHosVphLjll4UaZZNZO4UeuinML6WZ+iYTe7ycLrtOziPRCZBKscPgeVXXF2J1WAXFmWbg5N
nWEJMeOTPilQZh+yP3Dwtc2MSmGeu4um/aQFS6NHZAj4Y1/MrszPhDLAqvYHuEE7JzxBru0cpC9A
fmpcwWK8+zrIwqagNVLQy2MiqCUYs6KQKS3YfvcnWQQhO8bfR+kSltsb+YslT5/B2kUwjYWQAeT5
4JDk2HlSDSBhSE/vONnvgXL47aKHYRdbtEt3D03gzlZFvsLPVtPsI0KCNkZyXfpw4qBR2C6NehyA
4a/no3Z355MVGaGXnKMP4uA5fugzGb7OJhE8qO+y9HkwyqjgzXfAfgAIJ8PQQ1yGmLmms+HChAIg
R0Gneac8kUiBTY5pIoGIi2iMXPUtEZFzPQfvFs/s8D3UMrZ3Npev38Rx4SZZ74LTewj8zAXV1YFR
ElWYe8hUcX19XH8K5vgEHuQtqgNjeEfQf+nLdNexNydt9afIKGRTlOADTSmTU5LXQmi2cqSD2AC3
YvLgfiFOj9oCaxmlUn6isQEXIrZaDydUIOPHv70pcsJvkcAE5ZNM2z8ugLV1yMDiutyxlyDacbcn
QQReeBEn4RizguDgQydFx1Tul1kSIy/HQvyvXvoL6qvWtlj8U1yME43wqSZiy4EvzjQo22uGarWl
MWzkpALd/4lWbNniy/9OfiQd0rdKDnVh/XhLJH0Qj/yJBzarBjRngaq79DKTZon8vk770prmB5zl
eHPbnhlwnorqmwNvSUHae+p25fNBMkfRpZsmpvnZaV8p7+dcxGrkLJFTRJjrZshYA4gtSrHcXfHJ
5ql2GyewIy4jmJ/6oP8cxxkD+VaCXNFyCJsEGBpI8nKVSEGgHmnNR/t9/X4oNirdq7NVCus7L0ax
wfuuFoUWl4Aj+sMJzZ90IkVj3LR4bR77j+7xmIry0baj1Bkam7HcDpRdPc04EJf+PN9qDb3KkI1j
77aOSCgkP89B+5kUEVcFcGrV3JsgXLmXmsPVXNT+YKSb+BzrXYmJoPGDkzcjUIzWfAbOxvpg7CiS
7VfCcz4ZfCw0ebFwVy6VepHO/tpxLPbSB7LW8eqybj+wPvevOyijo2o/xsBEzbd3Qgg9VJ7/Qrsn
ZzyufQzykjk3scMo8ICrhcdcF2K50lIW62PrMXmo895NhCYz0Rs8XUrR/LtCtjtZqJVOBd0swgtF
Ldryh90PiA7QCG2P22XWoqReTQ3THmKg+NgtRCRVCEzh7HcHRTpfsU+87J78bL2FcIAVVtZzGsjg
AZ5CD8pL+4/33F2m3/xkGUAGko/BppFVKlvMJS5Jm5QF2uLvPU9uWcnsw5kb3vT4Bb7cOsgy9kNE
3xUXqAO3mKr/sPruFC1PkRJgrftyH2/Ucajj8f1q/2pKRcMmdA2Q3TKkX6B3pD97eHsXAwV7eRd8
iUNyw+/bxMYXCCrgaonJm7zBQH1GNTnqZBH5iklq3SQNhW7GKHuI0AkZXt7KxbeGXiKg964QXVeh
uDiewglPzyKibRvDUToHo1OE9HBYsFN78SHfqxzwqyvlnWGD15Xvf0ASolaGxnbFDb2RAeqOla2V
ZabAfNAnBjEFXYndQ11XzjeFhphagKL4+CnWtlpb/7HWmgcc7pGkAuVA8SnqcqdyTtHo+paUrEo0
y94Y4HmAs6Gk06H4Dnc4ZqF6X3eybXvDGMQg67seJ74QxMKJg3wnoC3g9LsRDFR4QC3dMbhMeCp8
1BOPBych+IJXfTFZVvh7ujL93EwdLTVSZQHLnZn8Rfa+ksfcngbozMBfwqtTEdc4/s4Vb7+Ilz/Y
tvtun/lOfV6IapvTlvuS/35VxgOqi//Io4/oAh2f/J3AXNpmvctKdWdTV5jMiA0XbSdMUaMMMvM6
Af1cBmchHBoEIdmY0uwfhietlvlA5CCI8cVydMKiQQ5FjVmIaQ4sXO0BGczMv+W6/0uXK1L9sdyb
XAldywNZ59ynvEb88VleBCtpqLh0vnRmZJkVWf98VRo60qkL8eA6Eand98J4vdBWGmclIh1GicV6
KgmRJmP9a7oq/0rlY7V8yGQcY6fghkxYN8rfKuw/VXd38OZSLiIHZ+rTb7+gwvI/hNYKzq8lOkLo
TyDuTmaeTerKJw+ttVN4A1kasXOEoK7o/EXaFScdwtvhMtTYs/++tWeJKedLBEl1n9BgPNGFnrlk
umpr92wjC+TTqN9apFfgrzV9s1toiPEZofUIhfall725ez+pe3MjPRaEbAMVM4EgyPZ5R4xkEONR
K73CFY6gmO4glFYLGRhirtf1eI10T19/SdgCVLl77PF8ZX00d4F5iW6E+G0uitH60mOlt2Z2Us91
cVGj5tcHbV7UMf3tzgPoenVPEYx6HlnDHUldYKIVtP9BkYoq2e0cn8SqkLobzb/AqOaf1C3/Rc68
kohVbBDKq7W9OoEPQl6cBkLTsXurMz6gou9KhZ3DafOS8KlPE5D+RIpO5jWIyANiwrvF5iH7Fx1g
hxnOPaiR4d6uQJxX6ewZVfzmdFhbYCxUQ5WkXLoiuv6yWV+11xM2xuxnfK4Fdc21cDqlFwTg6bCg
P2JZ+e3JWfvnPnmjbwY8g/MZu+AsUtYFVUsNtmOFW7/qCLyd2TyxH+EYAyBneiWarueLurEb/9RM
zxylk8fgqcj6/Xekw8p3bR1j5Cs+U2WuEc+NSHSivB2O9kX+nF2+aaZaar23wTOyMRUoW2bEiZlI
y86omDIxHdNS6tHTFXJ9LAOx5YpCJRs37vM0efOUd7DYO2u3RSO4lH9d03qhKWZq2xFhaaEqsvqZ
h5iwQtLNOIeRjW0Yx9gqwt7OXqOdpqxxATdXHP1Ck4R4Eokxfer/qY8RKrahQK7WdomJifG6TDqF
7uc8d5M1IYorznJ8rHpDJwy3CrNjuHDUIvY8YmpFoJEOoDkRC0OGl0WkkkrcvrrYOMCyVqYr8S0g
n1xU7ZWVZrsg4Hyiem/uU0xywr0nD5i6yilOevndwjiQc0iDhSFK0+Wq14YmssVteoYgOJ6j44iy
cvrmieMGo1VfAAv8dbSlWHk6dEXiWNV11cugfqW7qK9FjhlFUIqKkbAGR+qkkuhocaNvSxjPk4ow
j8zT7qUP6+jL6Rmb9c/85sOB1KxMWwYVksC6jfmQkMB0DWGl4r4GNnAlJ6M3ZygD13c0D0LocROB
gzNG1/lP83Cswo86BepF8FkL8bgR7U9zFsBpDorbe0M5mvKcRu4sbU3SbBgUjV0Ybce+kCgEeEhR
UiUpgCnUz3lD1fkzV57rv8lYiyFcHjCfW4cD6G0qo5DCg/pXIy8QZ2df48/Q9NZKImxC0YaM38rk
tgsXKbfwruzFgG6/zxkXsCLijP3YDtkBsdPnF/XjBcpTkP0wGyaXxGgKdwWzne/YYieAYT5Ctzma
jONdwvWdrgLPqzj7PuY4JsNSjErYb1y8gQKWyEb9AMAo5ny3xF60uIandJmVU0aEmgRO6ukobDUt
03FCFZOKiQemYk3olkBME9JqzRohtzla19f5N2rR686bMrFyzOPyzxsXsm/ZL1M57QxLUyOotVc4
b2b3w3v/JIGDVHE3QzIbxnUVDANcvOKBcDtPqXkbNqy6A0oD3c1chNjD1IPQHyyi7CIEqWbXrP8I
AYDuvhOv1cyloFkq0RglDIeCjwE9gb6XkIcL/AxeSEo2IikHQFRnu5F+t5BJwdKvgJKLAG/iP4Ic
zc/kngizVa/fy7i3OYwspOsC2y3Z5gLYIxhLbh29qP357qciW04AQFSby/ZItVu7cQL+d/hQI5DT
ojpaqc7HtYUiwDJqqNw3Y4bJeuxH5lUi+Prtowir/hCC90QzNVHX4huYkrJ3TlWnQrmh7D9VRUtd
GsZ0WnJqkPQdRg5aCJ157ps9uti0vNQIP9rC/FVRnTDeTIVI8bcgf18lU0ID6xYbEHgQxnyxyEvR
6ivUe8TAIaNd881A+SqUoz261OxebxQXM0pzTjmQceuPwc+3ufW42EwN9bT2AVqRjCcUDxb6uveV
z06ANYsocVgWgPG9bE+xDXhVi7ljuuwFjEyo3y5xdjFNCA3+D6/LGmEw+9D3v73HfzhQVJLTXq1p
FXlj5yMfk4m2mreYGlBMeMsc2WRqUrf9YSlIF05nw79RAP1vVh/lDHdxi8F6upmFP38JqbTc58DB
MBycrn+E7cMtGoBKkRXTFEHTxgPJOzJY/sj84MIx14ihE8SgoAKZWTrJwMNxChgUOOIM4aPy5ez+
SaI0fH8P62c9YMipHtctjH28fjWC88AIAnkNS/dDS8+dmnSMIKzYB/+sTeVkyyQKiNDOg8Xu2kPK
7uxFgL2t8a88DDfE6IAIuCw/H66rzazu5ubqJUuAlk1OlJQSODLkaejCsjC4y0qnMQ2VVekuntkf
tEjDmqZFosLfepzsBbFcPzA+5jwRMJp3001C92xuOBh54Zq4fkSJyIa/38/eW8KaDYIXsf/93hS3
4hHbK44/d93u93ErjBZfnDKHJwNpp/3GbH0JUQbtR2KpR/FTo8FeDu7DtQa4WSK6VDhdzMlGl8CI
5FA2CAlV11rNFrUoCqY3eqEhNotdDwpbBuMOsE9QKN+Vf5nFmvoE2PPDAVoB1dX3WaH7Eaz3S/ZZ
877htDGLZiL84VAtnbnBGiOlgPG4jo038VmJYEMe5gGvo4aGwAw7G10d0IXDpyL9v7URa1XTf+FV
AxHoMi8Je1LzuiZ/kYXaFNhKD9mMQD/+72zi4xKJgkbdmxrlTW2bXKxHe9u775jAd4FMJKk5fm75
99RHH6grCMtHyJKr+prq/0OxVmVOGXx8tHfPrZa1g03tBBkYm1x8ePKtnv5N46DUvPd1EskWhS2Y
JJyyc1hrBNn/7UXkNM7xfwYspRKXtriT1F7bjyedwPAPZRdr6urKbrlgNkkU19uuTgQg79/rCITZ
vCN7lvVWMvJwaOtjbmmPxtYjC3prqPK/X8CGbMdpV/ThdD3EpMn2NDDi+oCKvrkFaFVKgfo/khLt
ZyX0rnir1b4d+ksBxQWJmEEDgsYR+8fEHOfvr9xyx3bNJYbKNUirNlflZt5EG9SG1TnH0SZlhSRw
wPWLJLLtRg/pjuBVf9rCc3ApD6oYT6TXyIQ2Lkbt1NB4cVQ5l4S73nJyXPmGwZySURg1Oa87R7B/
+9yhIegHPO8iHMgW1KK1GuBIGeoKqYOHJunKRrS9PDUhC3TW9P3ss8volUdeCmptKfnSpr1UXW5c
QU2q9xE+K+wL+1aTeLJGZKGZjQxypBQfUcS0zBFktAhhEhwRIid98YyXi+qXKj5gYI+q+owuBKnj
ius/k8XpDqwoWJ7QmQ4BVEizR23iQ3VfwGfqdL5EkNLj3kBLqvGBnvuWdzx2FMx/4HjJtS2cfPff
jkpOEkU0Yi4lHIIocEQgqL89OcyWC5yk13Ti365wAZ/rRCRrXtQVkIsgyzfi+AmgJFRVBYjvLsZw
lN+m6D3ZMOcpDS+GsLG8jS6Vje1Set8oJt3AIKKfvgfMU1M3JHTSHmgvIXwXvXHti+BziDo9sdvd
4w0w6J/tDRSAumc4SGwd0KpSCcYwpiF/vqN2egFtBNmflnS0C1csMBH1A0TXVDIM5ln7xbKYfgPg
sI61pcrhjqbUHEz62G5aNrHoiuMyPuk50/adu3tPJOjo+GlWWX6usUwagawEdtF5+b6bYAVuiauG
gqc+YSIRatIIt934ZzByUMdMQBXouDTm9lZTXk43pnYI82Q52IcQOdVtCZI+LWHwby9rZeJGxqPW
Nr2vD+0d9a76xHXxAkUYkDlUIEZSnXlJNKES5tFGSt5XOumJUv+4M8silCbxRshTYyTmLBarPibV
tvzTprioaOHBUVMIOJh/2Heum7KEsduObdx2m6SML8RAA8cnrYOCRzCY/dGAVH1cxQUUvQFeiDcY
YT+aq0O9tMXIR5Ji1/sUHQs7eb81pFRv/gyZo3FqiClCEGKLmEtFLtqUfblQfgG/T76TY13PfEP/
Qr2bO1k/0MYfvV9iipmMwj/f6sYQOt7ygdN9wbvfCm5m/Wva6okV41PIbEtPt+Un6Trttb2ILgyy
LP8Gx2VnCfJ8dcci3Ph/ZaMMi27p1wezO7PKzuN2QscGffe2Ib5aXNUKenpb7aSEvhaVb3dm1gbQ
zqXALTRgoz9+ZXB/sj5xvCxD8Zc5O0jp7q2WbFIpor80bdD40gCx2V+d7gAV6CJmdIN9Z4PyY0yI
4yyK1ScipA1iu3i3PozDiNAuzbYLhfhF5DWILPYShe8kxszWvEMSmB/nmeBLTP+JBhGoG/JaYOUV
yl8f6zNoQYbSExlJ0EQQEqab2vZzaQD5DoLNUz0fVK6TtI5W+Qse54D5VURnZE07iZcqT/z0JjYU
zDn0yyJeJN6ySnEdYAeabe9tOz2mRkfx5DWiR1QcICKEpoX9bVLsk3RYqM8m8OaKh0NgOcqsSC21
Q9DCUGBkOOueh7IT6SNG86dz2pKWzjrdgki4AgtBpeApLlRucnZmWcsz3OM39bu3z9gLIIZumImH
pKi/8OBtDoqXheeZJHdcgLtmiuzY1F/od5BNZZli2iOy8zifc5RZSjaVDtlLzUkjmzzqnP1vL9tO
d0WS5GKqCjPo0BpmafVRa8UKGgRKM2TgBqa/p1+6B9koFi7SKhi5CAU53h/iLJXCT2qub+IC6na6
kNePtrYjx2/CQW0t2KiDkz/49RZn1G+GNo3rAkoDTLxioQrfUw72EwSPMGjJgPBFUj4oDv2uTeUi
LakclFyidBUjBFMEk2G128iEn821GZhFPjhquX+kNV0aQBOLm5pOC55f3r+sZZQEzY7Z6kkd6MgB
KUWtrtve3WCW8QmYy8HdEyQLbucE2C9Xm9C3HrcMPOWKNOtT0m2BAL5sOslcvXFYZbWO2xXOqwMs
5EjWbnAUOPf0F+k+JIKH5aexyzcb2p3sTOFSeWa81gfxsjmTgdQaiWzvXeHlSOz+TzzVxO8e1LIv
W7dJc4RxAoe+t3mXphlM0C2Xem0BcdJmbKaiO324bYiRO5kGSv3ygXDIlGbWT9VnAMZ5TGbRYNzE
/7260mIfZWArsgJG+8eZo8sLVaiN87ltxyEiyxhRt0CSWNxhHl/PyYzHZBfxcCgPA1dQiEeAWmcf
aitICY1LcnpgzCcZpoBmqluF11adDHZg4n9+Y96tKyoXmHFLgsyNukI6ty6bz4jyBFjZfGBzKP8C
Nz3/npJSsi4IwwGP+xpKi4I0ZccS/6/fEOaGCetXJfd5uHiWnB0scsqHQXYX+FphLmW0TbhxnEs5
Zf/vXyUJyKA8+1VpFNAmS9PdBM+ByXaYRG0tewdtVjSAvGTCF6KZhICBKIg/2cIrVdvN9WwxBW3w
nnOTl2VN6nnOXLH3zmShPVGqSZZK8gAo2MOr4TRUCqN3GWLsbA3b9oy+udK7iASNkzCxWu/je9cg
aqBdayN3hUKy3ahNbBkVEQC/A+Kdq2E2/b8NSnZhm8OZ4f9lernSqCwDIFmLzRiWxNwDP4kuZWMc
n62LbrXDLcSdnsrLrrZkWGSXuhJS07O/TSTN6WeHM/9ZoS/rNCtlOjKlpvCNI+ohJrlaxjYaQ+p7
NzwErCJDrt9fzxW6dAh9cbapK0wcQyy1yOcq74BhIp3/1X90tpIVGsM2Aqys4QHH6YGx33jVS3vT
tRHyde8I8X3/WaSSo0xXOnL9ms2v/J13cCRvujsPDDW6ZLRAqRcfLPQF5+y+PoVvDRX1wfoSxDZl
fg1c/tpbiePFMaI+qmOSTCxRxC3lPtkVDYRc/HlvZLVBQkRfVN/xUeu+z38rN1ul5qc3FOmw51mT
lA7mEjSBWqT09Hp17aKDWJ330g4x59owhQEi3Ted5Yk7xyQ/1J5bUgVFZHhPiYWJAl53nVjqI8pc
OGfmhKe9mWImRv6IVuxexUuLJV4DHtL7PcF5mvzAafg8ri3ZKfMLBvjXspv9ZrN+cSzDK09MRo9J
IZB0QBZGaMd2Py/2De+4scG85s17nqAnm0Gr7nkONB5B0Hwsx+p6qbqf/zL6MDxPZ0YiJ8Fdaxlt
Pu1tjBaYr7l3+ygZ/O+DoCo3BdAhUvws84ogVg8aLfMulSL05Ty4q1cx3ANdH0k3UjTIAXc1C1Xv
0XZC9dhysWVExqbWhD6zh2z5Tx29SgeXNeB1l864/9WDCgXfBSP/IBYJCoC9CddOL/E7C5qwItU3
B7UsvgDVZ3WDaIWrFWfzoDrEuSL6nf/bR/C9WFZL1lv2yHwCHmm1Nb2rLKuSyPNMgA7xfYy1hbMX
A00mjfVGRkGS8PFuXrHVXps/0dBL+tycUVuZ4XYtiLpUmAdCKKqd+PVuuppal7k9jTVfFOpni8U4
VA6NVIrsbGl9xJejrsh01OiIqm5bYk8n3kUNd1u+yYjzidNzWBVYSEPPgH+JsQvLXmxHSkACIzPk
5pLZSX4sIBM/H70dCYUNh3bHbo+JQbkxF/OFL73aPHhoGpHirtKEEd/4fkVI3gFoZHF65pFrj+hX
/tzU+yT4TxxZ2R1gpawh5w9+sSfy1iE+TKMRmw4xo8Pg3YBY5Dn/k2JDSQAk6hhu9Gys4Xw7VXbL
KArrqjq2w4dyP2m6HJdcZhPQl9Su9y/WgWHh7i/4bvdyhsyXkVZjwjQJ6OXoyXOf+kxd1cVtZ4TC
THUN5sCc7/NHPbKVCKHnxtNGzLAsrqHvNUl32Ck3VJH5gznY5ixEjE9mjwiLc7Yb7apBZLh5xMEE
Mxkk6NB9IZ7sdFjWrjSxYVnsrwR6k0SkibRwTEsXa296mAmJ6Y8VmBRobCuRgFomU4rXXptnvxLn
aW2jYpD3FItDG/mrbUwYWluISQHej5dF9LcUsTREL+MZlf3DvRnLQMwVr627ZpzsVEA7RjWRnlG1
2xds7mbsSwGjTIl6QCgW20EhR9HQTy3x24DSmUkpWW2ps+OGBpId0S3SuFt0FZzD0vC+V10DF6Bm
xR1YwWG0hYi6geeziar8Js3Znadsy/x6IXCCk6mrptG3ccrnPHQ+DljAYTJ0SmxjW9C2aB8En3HL
wjX76PQ7r+cZ3DF808pYJirMciobr1y/ME0TRHNOA1qTm7HQOAGilrXpvHyuMMdRuKHNzKuopE/S
sLZdNbFvS9YmvTo5Rw50hTly2Ey9DB8Jo1bz2GxMq2RJ2YXutpSv7XT47ELfa5J7eqGTNMPF4CX1
cMcaP3ndidWciTDbyssVsKjXB85r5OrSgs5uftK05DbnToeitujzkDE3l1bshqSd+TdzBy1/B4Lu
kuvipwLbbh0O7crBXBREgqPcoPT4Gh8aaX2IKLH5jkPkUViTN5d5PHnupqax75sWWonWJsfrqnAx
2y6ZI2VxaLz5SELhK1f7u4/eE0/vGoh0g8CSZeV/vta+pMmdDhF5eR3ULniOPlar2JfNEVSME+2u
YMsLPEe/8DPs8Rac1tDnF/ywMvXS6csliKNpIYM/mLxam8SmLwc1WTb6lq5FeETuoTC5o8b73+qo
DXqwaKnVi+Q6781FY1NBEd4U+Ie9IysrD0zVHN19+rKZ2otlZGVM8OwANdmX+8hrvtlA17vg7vau
tI7aMyM/NwHV991afGJV+oQd80Sh5bUJCXGFPuo5KAH7rIqvsOK+MUMRPoQZ65zet8NQfy4G4iob
4STyJ6jDNcXF6oqPn/fNuL4uWvcP2UgYSAwr7cfXhbT3lkNQgg3+UAweBYQL+Xd8Yspg8zGY93aS
bkBtm3L4DSWCQUnX6nBpoG9zO8c95qSBDOtu6Kz4AeTFa8ZlAqAIv7RsB2nvO/Uh5q4S4PZM8IAp
IurKyhwEp/7VwHEkSZ/hMmX9Y3LXNwUc7OyMHDpHttknbopWrUx05SnEEfm9x/9PUlPTdesqKFGA
JIw+OedrEvkpiZg1HXMNQhfW1mTopzifvS21xGpOPy5wk7e5uYs6YppzJWVG36v/LSPPWWu0RbcJ
AdMYuufZ3DAEBGwheHEk/2dBag3bGV+kwoCCh6innGzn+7Pv+wT5hj4dShnAvQeTs1YNs6StTeTh
zKVkeKQrHD+UY5pN1Cp3o7uSIDPSJAs1fcGsrkkbnLp/txdGlvF/1vYhcPidfI1MnGGeGNFpyBlc
GSfq7CkfvsDiGan98nTlDMvQ6kOSpJj2DSLtT08yw5/N1phyzWkHIpRajvnGZ+a0zwrJZdYZczKb
MMVBJKZkpix3O9nWVTrj+VGz+qQZDAN/cXzWt8mCz01BcWtZRAzrG8C0pcqsUUpb+izwFAsw650B
hzBOqBjgjE8ZhSdxNvRtuI285P7k05FcrRjWEaYGg8Aw3D1F2BYOJO8Sjay7jL+Z/l74/MxoZsy8
4zjRea/yr+qCKdqtEV9pgNQwdW5+vBUrkeGQcy0VCc1BSM4KPBEpjoJTUhmayIuqEvvOXpSgWEDt
yZy+DpPDTa58gP+MCopj2YByUaodkDaskcJZo2Knd/Rfg31BzInDltzwdie5+l1C+VmxSohGUiXK
bZ7CL30Q4WoA70lG3rSx236/MWSyn91AD+aggLSsor6SPOGtUosGRBnZYqd5qyRi9jYDB6HQhDqN
yy8QQ8S6dlJ9FLzczPbtu5RbEmPaMLP+hAD1V1f+bVPpftQT0lwJTa/my0ahgKvP9TZN22bb3Pn9
0XgZ7tzmEg1PAumqK637MgGEpdVp/v7Padf8MaAlsB8c9QSPmRGz93QLt/dnOcRtNpotonAjV0ZP
0SSdvhCxxKmwyxFZJipXsR2+orkggK+9g52DY7LHY2PUQH3FS1PHUUjU8rPFxiG0yGtTDo+4oQAm
KUPMbRhP4tm0xDtMkptqURotzOdtbOQvDbpOUcO8FWLA8ot54ZHCEfKbIJexm9YDy7biR6Qco41D
KsBIpkTrABN4S+M2aMWvGiZ6yew5BUfmgqRIadIQGNRbRfQ99+50uLuW2LvzCyNh/Ul7FBsJQT68
/gDHkdBt40/DjwwTAP84FCstZiQQSntXx8vM3F7d2GYXv6ulawe53FgJHoawiUV4u2MHJOZT+0qx
v7fQoV5OFBHLJzsFyWCd0EWQNpASzAkTXaoNYM5+pIqEPL34HUU4Iviz3IXaEM8tqk9d4+g3X5FX
STRFL3kwR88mkkuBiM5yrWJL2HURES8arwBZl1jZPQmoMbsgUuYNMAoqHGXVdEkRoXxu1xCCtdPs
pOf1jcKOjcPAOE89FM6Pr/K2JAGufl7Lclr8Sxd3lZfMJmzqG5DwSd7ANt7245LCERRa2c3kGb+o
Owj2NW95Jex6AFj7+pbQMr4LUzqP7vVOK2Tcggb9p7TIOfZV44SXDe4N1itLohjNG23KuB3QCxaW
lOi0Gagv3zKbAN8kwuYu+H3aAzvgcBYRVEHdIqSh6thlryY9DJhbkQU2dnjfvDS3ZdNYgNEDbV4F
6ukGRX84IlQnL5P8XzmDkRaLH/oHnZn0jYf68MYUQedW76DaWm7HFls4Mxo5rW/GnFGZ50Fm4bPz
0m6MnDlk+A4mgL4jEbQhrCt7Xo/W8DJj3EX302EPIhuQ0HFWk2OoQialnlYYLfQWA6uSyciIpIf+
Uukk6yZkhi7sNpsiBI2Rh67xQtifPIufKgD4N+HagPmnbNRtieLM9ndPKU/mFVfKJGPCwF53yhlk
ViJXo9liHwFp1iJOFy2+dnt/RZp7DMqBTzk7Rtt37PU2DA/K3qbw2n5Gck2xHKYjFuOHvuleK5Uz
3tLZrdItNfW/nXcF0P6cJddJnMbVf/KHh0xxzYpQEoBQvNd9osOSJuGYRv3doanINbUef+p7LAtv
X/x2XjOBTNNmX/xdKb1kEJvQ4GmXxLUZTQmi2i2tCJfKPGq1f0hVzGPg08u4hJCnnnhB8RbHzuVT
9qSH2Jfn8LL2e/zuQ4gDnMVc+dzSx2YUIbUtSq8HaBfIE+BGDXZqKmMmgcR9Bt4mxVWPi7n0T4gN
hMyL2SSK3lZIlI81PNQwdSxREizOJ8NBLgNpQWhdKoXwkXXv2wqCfu6yLjLPXpdGZhqjjnZoKBmD
eZI8m5pYDRJwIri2f9tKEMlxPtfX0MO590fZlm2OtSFAWESrptRUJexETDjrlpVLNW6AahjVjVEB
me+DyhElH2TVQfELRY/ov6xLhdyIUrAEWtyZzYd0liIjQXTMDzrm4EitO2Ag4HTZwWnZuVTeQJhp
bIOgYZ07uzRLVxAOouiW7ClMij7aojitPwESanOyUSalRroQfoEmDWNnlJlAGgx38u8Vkt9c88rH
S2IxI8OTN+ORScvvTOH9IJN09afElVAT0ixkYomnG6y07wyxChnoCqHE2YdQiAkqMg0hgS12w9/q
FC06nF+2Qw8Q5m6hmoYtZNlASlcGLhyIGO0lN0FeIYHRcJgFg9xF+Qqf6oA39gTMWB3HOm4OS4X8
ALt5/MtN1HvJgTO/gPob8Vih4SGllrFnfP6QvaGSKhAPAwXsduJ+SYQx+7HyoLvxtwKVTShvQgxp
ICYSrn/1ML8MabLXQWvaZhh1sp69s7dCTYnO5yduS/pVxvyfAKj+MlpiSYpGy08gtPrQxeHiNNPX
j2udbdOIiRUhu0gHTfHrgFxC/1b3r9JyW2ozy+G9bPHztjbIoy1KWQanRruzLRQRbWs1s2E6Mu4o
Kt+D17Om4F9wwOCCaBSF3RU9rLFqV6sYnNunfRW7UB3WI23rp+QUWT6U9/C7TxGNB12TV77wiPlu
MWsiHNJxESCfTSsdchZEdTkiGnX0DGoHRcb9fsBXheuE/DQYAy7aS3jl9TfVPSYF6MuLLHAs8bbs
Z9F1YrwVQo0Yv4CcMJV6H7ydSkkrUfn1EAqAnivUe9zdtm/GHo8r4O9l4sjwD8Dkyagd28yQChyO
JGFXcBpsqj/6lyquuUw0y7cgha9ByQn4lHVVXDVBIfr0IRaPsUwca2INUyTP1PjQalTe1agKIP8a
8q78YJHjhxAfVftaO2ze8p6fRlCmaYhKpNV+wdsLn/Jo93bb4W9FtU2/FkeKDwSjGwW8wOfE7MWS
8MkezM2xazih00QmU2TemfnZes22JPDVSOuy6zIOTuVNLjE8qURE8kwvxxcF12jlihdxv96YwKXg
uTCXolF95W3OCt6UbDvHT8xS6OO4i9mXBxJYSOju/LqITTK4AWLaoOamdU3KevqqIK/8IDJKnbus
MAX3ktzsfTSFd/mdNmK6HcDm/Iv2Fq6Se+Vqt3r5560y+xdSe6xsIwKeC2+5Tlp3h33eBIJ13lfW
dPngdw1RoUjDQvtww4QtjSY8BLosF5SSO66+tgsSt7e792EuDRu48CaLwgKWYMGk2NzhwsVxSW7/
wC7u9zjuTWGmR2yFSRYT/rc86eqJzPBMfwt1EjqZfZAD2C/1YqD1u2ASOBadHxrLiefblreKU5U+
pKG3ae0YMopCdeZ36iWT4FvY3fc3CGoJaE9rPVNzA4+E8mdqx9KUrliNZDZ/j8O2s5aNgEbIkMgj
alkZSK428oJzfRMjqVxXc7PaANBGmp0hp+7a9f1OyQohbXl9X4r3d4l+X79kfNzsO0eQ9WX1nBXV
QNZwgrnMOee7hGhVOGwUDCq0db91DtXOGeuI+gsOboxtsSN6W9FtL0JPjtjlGqN7tGLUewRS9jXd
JjuP/Z5nt9besWkFunqEnDmVXKOAg4X5PN3ayjyUPvRHQ1GUWOwsizPoQwFe7kZ3w2hiagbr1SVL
5LQrJWwSHgNX0tMpkAypOK4lmPJNEPQ5vuW1HPCe9vxPLg4fOiMCx+5Jrh6svy0uUWSSiybkKHmy
+24waNRU/1dGmCB7C+3SFheO7Q9gw+k6GRWGxS0H37dShl3J9i/PUShQzIxRJz6JCPjc1yyux9Td
LEJ0UiJK8tlJIL1rJyCTYTDXIWsS2evLBHJ0z9LeG5hCuI9TzbDEpreZ9yrStCfhvuDgG2Il2moJ
uOsNwCaxmvWfCBXOtHa9NFPeIQjmUU152vlzmnPrxaPZPGm7AV2D4JBGR9UFetQrSAtQGy6StJrp
hOIsTdE22bzB9WvvwCaH7idp2nMoTTm0MZ7X0Df0TSn8EqdQgIrs/bQUF6JfMbldXauIMkIjM/Aj
yTTNVBwmXRfiGI+ZmWfASjVQ68rqeJDvej4MwHslrdQuTSKBPWBv4pq5wX1fWztzlCOKQtcwAJmi
zfcTlzdRIZpMC9bFufwhtlOlLEuT36hy8f3Lo5w9Rh08tB8msqhdagi0AWBescylL7VyVhaYLfTh
lJhWHB42h/RIhdf+cqQrJ+2jd5SgyOBIyIVztq65LeARlj/eMpzai3LfQ2HO4WuaDVYqaZgLcwjh
oVoc5Bqoi9kIlUtV1QpPydDa+SA8WHOAPQtmbaP2x1pGQ7CpS+F84EJ+Z6Fk8LmktoM8EouqOchc
CGIR33eq+DtcBQSfZP92J3Tj3miYiEb+LdyNQSuabtzwcaZ7obsn0T9JtH2YbQGr+3VY60rK0dyP
446pT3olBCjHz7f411NtjqwlAWUUa3CYvic2FeF0F/vKBAw7zlVkt6ZTsKqJS24qTOTOZ5bKY7wk
vWy2hL/5Nqpg5GFfGDMB7T6fPCk6TcLOxA4wAYW2HHYBs8gfMINLA1E1MTGpA7M1Uu0N6U9jj8VK
VtA+wy3WS4LCEbFvGkLjxy+nbkQfKSLyetj7I+5N+ab8xNyMnTDbt8if9b1r25L4EG7n1z40sd7T
AzpSvznVbmOaGsTzd3UJ0CQ3v0ozvyoitF+aRZO8XWAOnuhoBmV1dQgCCUUt3alUQedRznx6rmUf
PgSEFjrC4TjExs2POEwRqGpQOjdcgqAroTnjmA6dg/niSIiecY3YBz+2nfiuFxdcBfTdX1jTY3Sa
X0I3T8J9VpdgS1dVEpsxEslyYMKNVY9zyqoUv72CINVaYOqKT0nZheM0oX0Y6smYfwha3QZZwlER
mqa1gqxnBgQs3rJApVrF6JNT789v515rAihuswN6x0xOZUBk0cguDP/9qAycTLnfo7E9MFnoJYG8
laPwOIXZ1VUhzd7lqDWXvLLnCFK7baKZ8+L4ATf/Wy/WPjneTyPVixZx+GXxD6d1XrY6oPlsbBow
H9sSlgIXS9if9zczzlfFNri6suCy0rZLdj47M8eGmqhnZe52PDkhk5X5ykKFot1aoPQTAgN+YWOU
3gjoqSVf9RmJkOfr7jOfhdynH4h26mFipKEKg5UjAR4tKRXvjvAFdOzW11k5xztfqO8vjfHr2d4m
L0i1aoEksCygocf9RBbrhqjekltIcoQyjfSSUwiDrl4jqCg3AuE2fF1YgxgNzjvrHpRBAtWkqF5G
QXl3MQ5kvy6LTFFUVugZ+5fefLxwgPTTOZBtockq20D9aP1nE5iHB/ith+w+xMkdAJCVNBqO6JTH
tzWWJU0IFMECtmz5WLNFRXu4pB0JnTG9GeHRmFt2N3SonlyvI+0CjhJUZS/6UezMiLJU0fsJ5jyo
diqxIfgJEssInhQjROzek5YozpKljrXEZrn0av3tDbc2P/3Ko9UtNztceRse9M4tdZCQHLIhdn5E
auLvzMKokzSko1HwfLexls8A1G+Z/hwACKmrcXHUm5UGWEb0htunP+QWJRqvnhRuDezUp2v04Ht5
Gp6m2eZTOQjtdpf8W4Axi3NcFJo52nm8EN0ANE+8sobp1mOuANO2w571JtnOhT80hVRAwJxcYdF1
5TCrVe9LW7lrk7bj3t70lJm32hU+h8/+9RLiNGSkiOsk5qoUY/xoEWHTeYdE5w/HaKZOCBVe3/cl
6ISIn2m31ND9OVY6HrOBAPFP1k/hWG1bT2VVNs8Plp+1kn8iAhwkxwuanpcHh5xdNnw++OLdVn0y
LPFDud+YTTeEaiAkcsT+0o/w6hacjwA2YOpPcEYHF7GzvqMT3kGoXtkYdiWRZ3V8ue+7XGVk+gbp
5EJ4Aml8cllsBavgTbNeoLMMTLVOats8BgC1em3Az82DGlLFUC94nUyWTeWbKcSG59T3U2H1qQAF
DIkbYZvOI7VSBwFd68ZIIe0LS3oulQoOa5JYvo+WSgkLvuu4Xv6fgMKLICVU3OKqZqRPGuxrUiOO
SqOKCeYtjZRsAHqrB/IF+wS2JND4KONLpX3VXLCqRSMXYBjrTXxMVnuN9q+vzUdUtolwEDpg8C+R
KQfft0axY482k1lCsIcwPxEWpSBhhtwk3q58qeZEyKj6v63c6cBQZPgBXuloDjBWAEug8/Bg3lNG
yLftkx9DBdwVOXkFHGD0Uq6vHr2FmFIkEcipFQ/THByK4GTMi4AguA1ICzLymAKzeFOti9AWcJYI
lAHxFiBA71fxekzEB83vc27B4oC+kyu/aZyxzWWmtTTs6viWKnWuBbs43ffJ3xKRr1OcnY1aYG4m
tazG1lKa8IOAYxHO5Fy4GgT1h0xGwVm+b1QaEA/9cYTpifGw88YaP6St/Eri83KTXP9HXP5zoq3C
yHB4TTgN9bIirg+8s2dh7nLOMNtb0mXwR0BJdS/dGrGvzaSDmec64LaH14pLZU8KqYZ7Nwebco6F
ac7IVjtwdUdfPteGUK5iuPIAbY0RPYbxmJ9hfJ6zxJvORz9kqdvSp4qtGakkO+4VsWZmyaCICCdx
2ZtXd+E9cwmnXSgsGLyfF5cCeJ2efRPaGxpZemvsV9i8SLTPdt72z8ZT2A9mYx1B+Sfj1D5v6KBv
26WB4dQlo6S9dPeGtAnVSVBfCwzgqLup79GziHNRAMpNhZm7K2/2YVIyWxK++i0vZ7PFQQxm0OFd
XcBN4pm2Q9hB+0OurFqJ7Fmaq/OzWITr0Lt9Rc9aK2BK5mejXR9SMTJxwfY2ZTZHpdA8ETlEntsw
QbFLTO2k5R2ABYxPPjxNs3ozp+hlSOLxhVkIdozB33MNktBBvBtkhUOTYkgY7cVDh1FX6NdtuhaJ
ID+fnpUWHvurxLC28+czdKT9iiIOJ8f7W7kZNsm2z1tKmZnLUb53Xvtv0rXxxsKrv67FRpZNBT+n
gCHrEglU2FZjSBhhsME1fInXEXmeSjlxienE1ZP5leq5m2WVKgWvK2x4YqSIb8plan8yPF12CUF3
98TfiJ2JBgpUJWv7tIaYcLwE9+dfYOvIulnA4tHuT7kFNefz63zsC1OwRFo9yURa50BzCCZaIzF6
WHKIlUPudzyc9UrexcQKwQD2ZVuEBJb5HN0stiiADMAXMMjONVN6f0XBjRQZ0q5aL3mq6+cBNad0
8ilvE2TXFCr+EnxrFeKDI6nnrGTxZDGA6yhx9V63Tr74IKcvHjRxQi9dQ1qZx5u5fU1K72Zyy3G7
6ZvYxTQ4g2WW/sHp+n4UmLm8GPFZisc4V2UxOsGZPw5qwnEsFPiA44NjRKWl8RINoZjFt+MeEVEf
oNwaHgrn8cB4A1n1FoBpn6muEgjOBkbtvjG7AKK0gd27dQHFs2ZteWtyISG77+y4fLhcFfnQC4Qv
rcAffXEUhkzWWuFuNXK1wvOTrIYKRS9Fa+3DwpsG9mKGag8LklmhHYLpjTA4h5GX4CyG2NcbPu4q
a0I9HkIXITVCbdSDF7RHLl3KMyCZ2kpAW8cKhIv+rMq95R6Les43HAv7yKocrX8LemMgvP3CI+Wm
u90x3Z2Nc2g/PDaykzjGs/71ylKeaMY2Fu4xXuMKGwiqN1TJoU69P356sNGxKZlydimD4hphwhN1
BRoQjtAonHrDaNtkHg05os/Skv/VFV3AygBaei7CWzdgBh0PjUvaSYdTuX/YELfmQ9GvmA6hzcuO
Krj3MucfU4hwsdNcgqtv/VwprvvkU48RwL+Jm41lPZAfoDNnvlf4NwN9+TUjr588nPVcTRRpGP/V
nfeRyO94Wegy+W8lfhn4LBo1kNT6OwZ6qmvpMxinf98CK0y34sPnpWsQlNiuuPqRF/VAuh+RyBBP
YnhSTF89nupI2OSzahJnydMvvJ1F+g/6iukoyn8pmIHDnP2TAVZcUn1R1mY6ZqU1rYYh5Hwph6X2
ZKOlh/Z15pNgBfk+bfh/c6HJc5kd5AtOkAO6iMxBAYMyyfPqy00I2wEmawkgOx0vpmjCx3X7woEW
GkN43qNt02G+Sk5IH//TEPoBTDKHEBRAdkCDi2M8tpmvYGPpsrwwcBNcf5Iz/9to6vyC8xZDd97j
HJxH3jDm/DInqT2tznb8uMhwzO24YiOF7/mKK2HdKjuZiwjkjP2mfAP8x0UeRcSg+DzUgAdfAjFg
5SHc+EPsoN6C+ySRgGG4JsCONhf3XKqVJIqaq5oKC/JACLr23IhWSzj1wOuB2ZJ5cPT4aDFy7IHE
ID/FmICWBpRVWIdPWGMvFdE7TdZ5fqyzkvaOuiNtBuz2AQo+Z1itHN/eI1SXyAWwaSLceEq9N1HM
jrPbYPcvWWOTRIPmxoafQ0svXNb8ceiqZs44ckQy2WEoqGi4InhHsroyuq7ljJAwdiNGj01GgWgs
O/jylAC/a1THTU8djoAl8iwMsnU7F6CvCzKHhqYPLjNMwvODCg1sBtzLvlLLq49ot99eihjbY0my
yMH9ron1mCmEXbBdWZcwz/J1V9izQLgpL9bUBht7yyLu69ITRHv7grtcooFiOFcC1TxGJzNy/SjX
3BAzje0vFVgWJXOnyuwudhGIWnrei73MXZAzGeKueWG6mIhzsYksE6Kny51rgSvyeN3aCjnEhemE
vlLxrGTXIaivChelBqjL+ZOv9ujLCVurMCU1jwJ1gHDayRvlA4VZ8GEE3ZyhDRVMJ2xQs/+ogrWt
Mywl3LZ930flLreuZbQvw8Uoi1oO66GcXaU553DT4jApEJ0J2JFKFBRjd30t0t/TONnd8CIasWkp
6JS6+Ajr9CZJl+RH6u8c8IMud6WAVJV3P7GGFYbJQp+WSILAwshZLGtnD1TybG0n1LCDneow1E1Y
RPHqxxtNk2eYgWDMQv4jrtrBbXPURM9WIlTn7eurHyzcZdY/MtL5bNPBGrztPySouzUbvQgJl+N4
Bcxgh/klTu3DY5ZeL8DcOFF0pME8PfNV0XiAVQi7VD4h0830w6KiDCIRa7kykCeIxnKlbwySQn9W
+nYf8H8LJ3KvVbP2bvS9sCSsM3nEgbl59/oE2EFtE4ZCSXSHPRqh7J9HIfBGdEBoRQUAsGiNQO45
sGlobTYbFGUWyhpFra+oF7U5gQ3mnOO8uN+6i0/MVZ+IkMbofl7PlOSWCMbaPI8hnD7UsiAGiGgV
Gbc/4sSAm4v2JKvondHt0EyW5GLMac8TxtxGdpY8CuhrnzizUFgc8Cz4Thko8WaOS7rjU5jLvfb9
zZVuYJ8ulWedlecHHQmUaMLUfVo7kggLXyQlIEDLK0eGNqgtxXCQXamN1R5OjF7N5gF1+gl2Mld7
5wj5hg4lSxrXWbJQvJr69OsfBiUWrGdlghsCsg5W2QGU8uaKXOizm/UNMBZHmv/65z9UMXUpWhLl
gK5+rOI+O3NoIvQhRKkJsygVd3/cO0kveq9gFS2lL2IIPxua6StERk7cWVucSGq0wL6KDFxA+ba7
87mJi9HL/pMklzKXOsqK4emB0r6oORjRrn2gf7xUMl2FC6AHaGzSQE5NhaWKl2kSokRC55x55LAm
R/+t6czeFnunZU6prVfWqFPrVDILnplZiTkcwcJ13Ttsv/OJdDW8cjhIrBfvSO/dFSrUxBDbJY4I
mktPzbS8hx8LLF127gQvmEPSS2hcwE0iW2lI8oeQaFZ7o7qBlEzWj2EjR+RJfDnEBtjWSIT7SWl0
EW8CK1EZwap2MeFY6zAHcIpxJ5OrqmMU/4DphboPpy+D/MzNVIS5LG1dou9Va/wyHqzpbcTzh9B8
Lk5isQl9kMi39Am3L0a/xxkNd9jdfZdqe0y5rXz23KcT5mNBRBxZ/HMrqA6F8sdPGOHPeK57Z0Cf
vHV6A+RHW91EeTaLipNxbc/I/BRPe+xDs3ykJV8RzSl3WQL2pzEWgog7GrgdSTvHEkA59rVbf2Z0
vX+RJxb4RH+xJ6Fs8bdNWrdq2BA1Q02JEFM0EvT5/j7WcS/G0bsGqY1bMcCTbgehaSuzP+IdWdP5
mlIsGQeXgSuoxrZQRmoVhQVLdi+E6AK8thNtFO0VpotbJR8qve/9OefLDV/q+rHk90J/8+bLfiwe
IDaJxkElJg8TJZTJmlc8Zkeb61C7FQ0ZSbhT0m6I6KMH6ydYjsp3BNRGlZWNM2XX2dob4o4kb9+9
GOtO996ewCHhrTg4Qt/xUr7LZPF1VwYS0O6W09m3NUVsZ1C5nUUF7SVBKeWcNCTAC6QhWBjXqgtd
MJ+QJQh/a8Wp5rT4DAIqbAIQ11KewrNf6yvfXt5WLCWCu7uqjp1+S7vTMY0vzDEF8EQImHISRG1z
8UWgf1xbDUq/jeG0HEHJ8103tAFKtUPu6yxcpG4Ak8i/jeUXioOhjnq2wm4IGlnKmWW6bm6Rmz5p
50+1xm4eGVAFGm50ZQmxbElaqbwhI8yxv3J8DN0FHsenFJ4KF5XNQV60x66a4jnUNy16RPRtqt66
6hZTyOBLiaFSEh1o0/SjdNnpdGNEF/7BYPO3HJA+ozTC5MOaZbVkDPr7+kRXL9bfmn4O6+r8ctj0
nJZTRbwYxw+F6D7MT7CFNSc8fgqIiBP0qxvJEvYhDsuXNdz2+P7tDSiLA1VwUHmYxt8OatM5UUjs
gqe8QG11b/g4ZmI/3hbFVGagmeZC1tXx6yCUjxbLFH3FlNvNGSJzpSnjVM9mBH+LmaIARqW50d+a
RZEk7higMf3eJ8elu2DSOuPAJWybK1RkwHEHG/MwKfMzeQAxeFE8X4+AugH3Ccgd2IvKc6OCZ48p
eCeK68wkYGdUXvQe7FPKoYHab7/aOzXbND8yCoY4Wx4O2AxPt4Ek8Ae2MI9kE+o8wJpOW+Tc+UAi
lnJ1YUEgvQ84TRWELmZ72UPavkB1oX/uk6y4VyxowRxwtoHy8i+jk6xhNRCRL0L5+TDsz6wO3RpC
7jRFiNLB9YSBIjD5p2yhuO5LYC1hOBUVIbymRDQT809yZAtfMnUzlaOWriuGqHeWPcDtCPoBMpcG
XQY8hcC1dvyejtbh9rMDF06TxWPlD9LrAyBoe18U4woA3crrJx3QyhevvN4/s36q+9QzOgYnPkps
Iyz0Nj+NC5GvykLOAv70LNedYFu0TfE/U0/YL/9pGj3Gqozsdq/G9fpurAWiEwD0YyvabpETVvdS
z8VoK1ByYWvcdoN1M0+17p0q3TiD/VWpO2LRKChOi14Mq/K2AhI5SAMWghDBnCl+qUbQ7FaJzr18
vw2TWTsKU1GGzwud3YUB1aNl3A58RVDHZQKwo4ptJHIUjOku3IORdBkFR3pCW+yHWKoD5Uu0Th8Q
drWaOC1XhpdG6T36ITHcDdXDZFics8n7v8aO28duDDZYqp2X86fsuq0zg/JoxIQXQYnZBPU7Jcb7
wwl9exQdkNIaubBoq0+sK1i54apayx7NV4bD5f7MtEgRAEMXRKwsnnfPoD/U1SRRm9ik22Jpi6zJ
wI1/oJemMAXgZ4QExKLWgMC+QgEbRnJyMHS3ATCTnu6MNe3pgVzTZdIlqbY9irBOFZwacKzn1JuP
rTE1S3gJe/ECAv5gqr8SapKLaIfoqXWwDQxjyCLNtMBueqOOqjhMurIb13ajdtQKnXcqa97rmbPb
YzKVTWRbhgCUzHcOJn6QqOo+NbWxOxx5CUF8EvLj27JXjz7fupND3HrnEkyOCB0yxMwvsciA0tcK
a/cnsxSRV6ohpqIsSYj2YPEiIRaW0SPha11lwVxAuXbIqzpqsPA21giPokBK4HoqewZ06aoHrrKW
KAFIgLA8JxVZLAseoIu2txGdqVOgWd+iZwBQ7XjempOpwOlqXLKOE1t89UHSW3Epl2zp2GHraj3n
R0I6V7eZl6AobycVcFSJMISrLWbiKmYHMhdvu6yM+b33Em+VVybzz6rtznK6EW5Bs4XIyJyvNIBe
k8jDZAzOaakT4SSnP2yz7byUEFcXljXhAmvmMa8znQr14ZXEZgxsAGEqYE9NHXv3r7+TSd8va3Ms
/3+cGydLivLY8WeVBFVqpF+v7VAUoiyyHmdLvDClebSxqcFXn4oHgjbC9cwpfyW/aeXUKXsylMK9
6bUr67mPUm9xvokHNOeqI5Kz+8+fDKN5wHJ47MVpPjhGKKp5yWwMDa7B4HD+RDQDeEzM+T02VsR2
MFAEOkoZasMUv7rPcdSN9Z0hRfNVzMOXmkd0RVd7NthntfR5WuJqcmvWGbinRtWQ3E34HMZ4lK30
ohXHpItBBvGBD+8WmSNucegKlm1z2Oh3vuNhNKUgIXRJfMz6k3324y+yWafOQDmcywuvdhfDsdhr
M7p8dT27P4/LVkbFshMJm5nf5/dU3pis60K9NtuYJrKVEcvktUBTKipcF04+2wAR9XYyVvL7+AX/
we4uSxNE3+HXi30vOOxQjZSiLQkDzAyt6kP5JKDz/gv7kWS1sdQvp9gpmOI5K4lVzVWoO3g3bRNO
G978+jrzw50jpgsTV/sdx3WUoTJHka0CgTdVKorY24KNizCE3mKoZYjgjCdsyRpSdJtMNcIKHO+i
DPZPcFKlo1X/SfS6voRulU60id2mMVN+p4SrUhr6h5NgxuwRnn5yZjHQfb8GRo8rGjgjXaZTk1MA
Tn1WMqfkjAoKQ5s9ib1ytNv5k66/tauuT7IjfmLTHWeV39vO+d9UpAUvn/pyWBMsXVzQ2xTEdAx7
hy6T2uTTtcx1WiPJyb4U5OC44qLRxP/shAz8/HikkHIzl3edcva8dn0rCMVFa6DVvAkUbcF2/JQY
S5DAQlK3OkAqv4jfLjgV/tNSuk0eU2+4bFMTXI+FoELg/YSehKc6nz2WO3eOxpQByaM0xD60nPGe
ZiEyFFkikhEiY5gv+C45ZVBYkW6cUjh6hgnMejw7gdYLbn10IR4RIFL9GdX531wXEgU7Zm2SRPnT
n5uCZnYAymrA6JzKr9s36jg3ya0sbsUcRLN240iXLyuUu2Naf8qkR7473elgd/+vhHOKG/mMezIM
OJqES5AqAdtOpleRRYpcWVtGLdTlJ/Lof6Klzk+2DgI2/PDXybcISaQhhGCIoicG6yrV2QrXOY0E
l8B1YOQRaV4Kf5g45O4fm3pVJx5fFL4YW0cgVpdFcv/X5rR5rqKiJFrSGbm0h2lX9j8Wxel/K0b0
GMz7hCuAKCtlZxuivu82R3OumHZtAjJ8+7IIPozGU1IdD4vcDgQlcggt8xZ8z0TbklqoH48IaZN3
/6L91li4EJW6w33b+7GLWWdCZbBkKmWE6fgY5vvFVGkRjZSKAchPaZlOkqs2T6IRtLjXWJaBkCjs
CHJgEDCpnO5JEWdWT4i8r5/4tLNe8ybchM+N62pVAtcqKFtYo5L2TnYa72kfOOUXxfDA56Oxe8ks
9m93mYWs2ITv8dJfsPR+Fh6T0Vc47kOP6nOUG0TPtNzk3B/K/ogKWDsE03DYG6GGrM4+IEczpKr4
tMbTk125g2tBzT2lypiA1Ki97kjbWCDN8KyuUljEwWuu6Gk1V6ZktWDl2OTu4Akfhd82RkU8ofYn
R8vJAW5YkzJvRYBRXEwJ1fW15iCvz9bOf6lBDKXo5zwABeRYesVn228bHUHptiwxHHCNeDUzspBi
HI8C49qPMmqDhazfOhkEyvQk6Sa8q91DLUJSpOM9FOjIDtUsj91TMqr8TpAyH+PySwVyiFHOzSNz
ENnXxkLq5cXPSWvfUjUC2J0U5cIHf9dmSdRB3XTMzaqMp6P2qOm4pPDUJsjlHa0sC/QcSyCQ7chT
pkj4EUDjycoL1bGdgyF7O5LICI30dBtUuE+FZezlnelHZpODD+V3e9BFgriCXsPGIAlkbuVBVHvv
saD4+D7uZZohbNVavm0OeKekqHikZ/B5G3wKiMznflbKDlxAss+a4+O7GGDIlzPD3vzIM9qeXNjG
4LqeqVig85glX3jkIgd9rc9FK3TXiSjW7KsoE3A12wEy95h8j+b2Hz21L5/eLSjGo90eXEjkzeoC
Fff/mEzrcaNlOwjuIQ32RyKhcsY3jUb1UwFxDABH1o1+zvSJ2tq+9D7U7ryB9D9f3ounE7Jr13Y8
Z3WyFtyQoMqvytxs2z1tO8GQIkKMdOdqew/Ats4Hjt5y16RQIWDPiPiXnnMXpY+cSgrwy6NygjIB
JJ7QwRvLoFj4NAWCC1Ci+oYr+9btMvNi+MO7nzjSu9fgXw60LJapKI2MzxExNwfX0dvWhInlExQY
bkZEPiid/+3H4tLJP+4ET9zwPj+FQYjDVIpRUZm+KSN/4uKW/j/uib5qvbOHgRzCYqOa67wBac3h
Me02LvS0h/+FM83QahAMy59FnM7HpRvg0E6ohuSqOCYzNkm3Fgu6hw9ERO1OpLyZkL8M0wt3rmxE
UlnYb7elOD0tT4BY1bMrB7Sxd/BxhE/xOm7d//WusWdqkfbX+EcWHoDRL8lL85o1IHmsNSg09Iug
20NO/9GrMEo0S+UMtnHbAnZNX2Ip/nwAIxJSXbuU3H8aTDcAw9GwHLsl34YM2BweE3tN46jV06qV
DtKC7nwMFiApzMeJBJ6VUwjtDD8+lYY5AlqIck0Sl0Ro0mFGoZ4yogOKKb739GCK9+czoHsl8YWg
Nodl+wiP6paWR87yitZOH4bxQJekOW2JwkHIG04DVcDoQ4RWQ8C0T9hEQaWTI7ToO+JrZDf+vL+s
lyY41HQE+P9wEuyqVwIloZHe/d2lmMjZqF8EaRasu14FtRti93ueIz5cWVzexK/YcVlVusQYPqkz
YBtq0YKWcuF6Lciaf0qY3eM/wkfeOrlrJCQa5knXlESDfSEqw3qrmB0ccVyCt1T7WZs0S+vFUoST
O8QldJKXm0TKU6ZDWiwpG6bJan48r8v4UJhheQysaXPJ3aNSzG7+EfoeA4lbgb9VMyD/hgPGUySR
cz/b8C7a/PFayHPS35Mm80JxAT5ASU6dV27dnJBWzbP6uA/JhbkaOXyT+TstTOqhEwjpcbW+BohX
Fg7s3934uGgnX8dUkBmSio+AhPVx9OX2y3/YXhVhGzYdPWMLTqEkHSi9Nozm3rUYYIKrR6u1Phjb
hKjcELpCv/Nb3tZFp2yrNTzIculHBL7STwqzL2lGf+es2ikRpWHMi3TUw1PH5jAxi5FDOt3OIbbO
6aiZ5G5oqJGnLIvSzVy/5B1oxG3OtYF5YunbpyYEgcHveKizLA8DFlh4ref5Qqpi5BbDqyjZXovm
aqho4SbJtgBJZiHOKxXmBPqRkX1TvK2j/sirWK/uRLZzTLZe1+AeWS10aw+Kl8kHEXjEmPI2VCuf
DRZLZI8iw4BHpBOw2EvjaUGT3SM8qKXusi8kvIzA/KVQ/1c8QkAtviL9tfjfjCDFBKIciZo4lcKG
bNJWITf92ezv3FlyE8G2CGMudoU34Vr1ihWj/C6E+MV5R4KjAOLlACAnPP0BNUeUlKl2dXMndNP1
SY36Nd+wxahVU0Nw1hmSEk5K/0/1wrl8CQBCPrNBUk+xKrGcs9cMqEALQMhGJXlmquOzVbNio/uA
9qBd+dFQI67uW9eurj1od5NSsG2wqPJcCqTFEqJXh1IO9TOcq2l12Vph0sFUqrA3Qncb0EMhRpRx
ixAgWy6+yKj1NF+pm5KynJxuLxvU/25HOBZYPySUyDrz47PaeEOvJjouTc1lW0UaQy/SVYGlqUzl
PCjoTWBsxBcYpmOfHGlbmNwdgeNDDBgTayCjMHpNOccQfYP/YdN6ZlCEuQffUuLBRiidj/SOZvIy
ERU5onX1OxWCSdO9Jk8WiYIHIQMUvjrfxtBAs4aTQ9GtNFujYVP8B4wysoUCBNHzDtJGo15cVJ9w
6w/u6YLbMwtqqEo6pyVkZMgsTOB0AUYvIFlYehI3sew6OGAHSM5r4uzw+NJ8rpjYlvmd52oNZmMP
oEWo4FXQjge/ne4w1LhtYPDaF02hdpnFm3neNp/lL4LU2vOlFII1L4+88Xi8ztBFMH1TuTupNx/P
W83JWzI9X0f1/QCuu1tC3V/NCR7OFoPLtyp22Ow4k0mw9875Rup35iZ8Xdnf3WJ4pBfoYSzjSiR7
Z/qNri1vRWsmvATTiuqkkRfCokaGwP+wanBE3txfCtdCkC1W5UDdeougeWXCrxuBTKDeH0Zrdhhm
J1ZkoNRmtDLV0DLNd8nL2t4K8t9cCzYHIvE2EqA2HrqQEIQoncQS3ol59UQysI3EehVE+3zp3Om4
BTryBXn3ahMOyS6Rr4iCSO/erWPAC/Q766ATEz+k1qGTJOaU9G7AoDR6kyJ1kUCfXmt/Z7ySWx2F
s7OSRCAWJphmG810Qz7gCoTrbsshV/qYd7W7Rlc2KB1oVyFgyCDIGbuvrBJFGeAzZVySb0tFHmD+
jf62nqy1BJskOdh2QPmy5RPOxHDgIgK4kXLrn7zjo22b5LCuN6eem5VqxH8KQvDNCFX8uJ9LT40O
L7u4voDgzv3XZBIgRRn/8KalcxLXVqioLNGi8YfjdalIL/7xE+6pHqsK9CE+WD4mYhcjMEB1xUg5
WgIXyKNAbP7XyvmfDqB4uzGsiM3Pvnhk79F1zIG4BRDAGIpRTsRkAl/Cx8vv0IRsjmkv5Jh8Ov/g
nwTaI32q3o+e7FCcn+He+zpUqWRqsTcZz7e8UCV+e3wJ0FSu3gvjMLHR1PKTffr5Sk6TooXczsH6
wbeYnSzsUJYyQSmvU9O40gOIv2betSY3SHh0E0iumvp9QXyidv5QnHp6uVTDQgJqHei51V64AM1C
Wr7uJj8L+4wbxQcwYVPUsq8mPv28LWwTzGA1xLsDvvGTVU6ck8R2VcLPNiewS4jE9XuDwyfBfu7u
+FGIIInqwYkwwhhWmFFJi3ERGVyi8G0BtiLYR2TyFCTQqA/WbWj6id+EsmmHPl/X0TB478tmERgO
9qhxXloQG2yvrapKEzgPh6ONnUgYiWfG910EYF1rJcd93O82lQ3qP9CSq2l/RsJiemUWiSzpnCUI
nFz6hCxC9uGK4ZJEZ7/xs+FdZd/upHx8PaAyjTmYtUuBuQ0tNoali9MHP9txCwIRIlI5KLLmv7es
kais46CfDNbHxLpDAKjN+ne6gjqVPV3Xb01uDiOe10aPym9QmuFZk5tK6Xp23kjEdzGzc54T6cKU
njF2rX2PIlq2tL0m9ghZtm3Eq4jidnSiTzgXSCpr6HQm5xnjkbsMqzvoQXas4/rR/0K0KhJnK0H4
7fbjk6s0n49LcjAjCOzHcN3rUqkUFa7qiukGHHnWYgn8wEEG55IOoRUw6bDP/Mz9tPRJvrqOWIlI
KdjiCSpsJjIv88Aihkl8XMD2jd9LMzVMf5BYfek9cL9PXC2i8ooDqY4Usd6i1UUkBh8XUAgV15B2
7UNsZb0xZpftSoM1oXHnzqbaL31JOEbyVslqxB03AfW/0e4CYzA5AY92xw+v3ai4wE88xE8s66s/
YEiQmmx5ByPEJPhj3DpnT1ErDfr9ddyIaZsEJi+ZBg/Og+9dacGhjCaaU+/3x530nIFMCNztmDbx
/QrcmetglMKUYEHStIVKolRMjG17zOaEGaQeeRBGXqAT03nHCVUVDgGzMBmuZoxXJMoKsf3hDie+
HdRXfhrHyyzBpU+MJGUFuK9/GFjkYqEi6TohuwENwOLMuRFWc4k6DXqdvWYHskISsgmDkSgBCGJ8
kRN8A7mWtqaDq2qT7jkzV6cL9Nw576HL/HkGGLmxUREtcKRPT4T3t0CQLRaf+aaSTNcNcyCSWIip
WdpzoyRAKhGelme4L8WfnIYU7lHoJrtpp2CQhFjL0Wr2CjuJ39Uyhd1mqawbxgBy/wGyKy+91c66
soIf5VzyHmJFzFwikZwaqVwPdRn2vPKxPNb0qd5Zh+t/HvyIZbeQbS52xS0CEnscwHqxh3jByjmO
3iZ6vt0IcGvr5HXe2rzKOTy2BGHbj1sMF6u9sDJkSDImiHwe1l5Z5WYG6+t0M9AyYKPpj9y46P+v
hDDR1iT8vNrTV55FnFbjQgI+kITEogCzk55gadbg59dczC+noW6oTUESC39ukax9IN79tPdHNO+A
Nr9KYFfMJqQG6RUHYCRDMbDZ20t7kZuw/PIbQ6HEDJtISC1XKShCfZiz0p0gL9Jp4DrtnB7+xYy0
v52LwgJ3st1IoCFsf3VxfIvP1U8nSP7BJrCbhKLD0PETLEdd7IW06+v85Y8w8oPrFHAqxbF0ulPY
Ffi4DiHul+ZiM0WUijL3Pgqaemaf/bMQ1lzGyhjAVELqUqsGnvdT7P+o6GpcQpLWCJ65NS2ctqyG
fI2IFU3BWxSXVbWNpytwlNUWjtmOL+KwyZZp0ybeZRQT/SWSji/0GEn1OYTD/Yu2q1gtO/kT/LOX
+dU0Si+As/shBQnLo9qKnBdlPcxb2gR8dSoM9r+ciaXCEvvxqOSe6wmzG2CI0WNkVTJi6bkR8sT3
oiBLktEVu0BgKd7u1yRC4ha6oLsMXbkJ9RI84ziAL8zGkcM9GKsPcjzUQD6W0DQqkayKyJyED82L
LdYVTqtHS9SnZSmSKzTfJs+nPtTDzorfeBr7lYdFlx1bmxxMfkiDROdymC5Ai2ru3t0KOnKPaea8
sUWOD3Gv53Iof+umWxuKUEgkl5ir3KRB/NDmBE4+mQuL4QhEl1oejTDk75Sj6dBJLm9mIsIbYmfg
qKZAcjZzUNX17CYM37ZaVgaDC+9T2D4FumRZLJzlNnYORDAXiTxf5Hows+E8BjzMOD95aQSuzXW8
Vq2N80YPSXr6EkRQcUCoG4Im71Q9T4O8djwANrUThcf/qllHo0oK2BcJllRcbsqqi+X7jy095VmC
v/3mtyBnVigbMUn/hR4kkymfTolKx3r1/ATooeW/aMo+gQRK02/AshCecy8F/6XlHkTNRSG+gVxd
egV76u7gfjCjQrNytQMiuieS2+Pj7Hxg53UHU4QsyGvH3kNWKjHdtFdGWyooHO7Fb2Ax36i7ErPg
TtbC21xWprcogh5wRswMcum5f2Q0FzIASr5bkKEXDlSV/Ge47bdaj4WRlfLc9rhWoq0TGop2heJz
XsPysJvgpTOWaQHUCUC/B1fJsFzZ2+Rx+zhT2caoYggsSHzUeGzgDYUDZZwHKF0ywN72whL8EpXF
5P8G3AYXorb9ZisnxbeThRgJaheglKaweYSPFlRbirDm7zoVtCwSAqOWsMbqlAcPSfvfUUY6iFID
d2gBbgfxOAEPpnqt50JCgGgAV1VmfrZlvbCioQo8P5vOQ1nGSQAa0R2HL585ZSpdxXjT+SeCJBLG
MeuwTlibnrNy6nAaUAAOXIhws5phefJyqS9MAmaPfJ/kgE7rnXbGCLJZClTP0M760W5zw3BT1dL+
vbiL96vhH8ynX21DCmtggW5es/CM5iaM1Ua2uYqlV3MG5gBbXhB+jKBlvRJZDnz0Fjy0MkfpDPnL
Ho0jvzWjToLuKG+l1mZroQLai/9u4ujihIgRqI8cABNQp47a7bYqhhDG2X6q2gwgn7LBHSML3HuO
SNBOpEau0Z4debvJNZOjZINzz4o+qwbGxxUxuun9zFibeRee3jFqM7HHG6y1HAyJNYSfWjaZVoHe
gTu/7cCTDVLviSB9jvqBBUIsdniGq1uXYwMrxbxu3m5BjVQ/7D5fxHod8E5UleNA4GE/vm4r5thw
nns5F036ja0ZM1xcOLHTgwV/QwNeia08HGbx44sAn0+Ez62DBAH6ReGG/47DecXz8cyNQA8URH4T
DFF2nHbNGhLRhTbpYP/iR8q5npQFsXYhUjjqvKnCGp+ZF/Ekkgacsolxd6wBrzFUKEX6x/Yl6CmO
7+8g4CyolvdfF91U2APGIDesiK2ZQpDuvU0nRf17BWbbJurxYqyyrEdyXPsFN9bFae+Ua+LwAIyd
FWxvBNyVbeNA2x+YwvhkJPOKMyf5qxrZ/NZ8eFhNpVL87zyA0CW0sPb9swztwRf5aDlY5OlYDpjr
b1YrwMPiylRjGWbEYHdjKRIYqmo358X3c/GyzaKURqNpDYHH7wgwkg6hlyxtwTR8GJG8FQMViCYw
pK9FNpzwKo7pePNPDI+7nR4IqniXOjBo80OXtZ8oNKqs4G6/BS5X2PMVdW7PslNSrrLq1fxEVhnJ
eN+MTQlbmmdkmdf7CUIRA0V1qcOND5jZE3h2eQ1zIJAZBgOnSmbv29T2+ccnZYUS8DgtTb6pzoEi
+X2VDuS1gdsdB7xDxnDIfKMwt1GOwAv6oPgoOoBHjJCBr+6jmu7f5siUt3z5vqVeV12jM0kZMOnJ
mI0WL6UuS3SiNYweuaa08oK6BPct40Qr72qPOcQob5tmzcrEvBFcOG4wlRaLaW7RmdzInfGZkb1E
0EivhI8li7jA5iVxf2CmNS8pT1VI7NfRbq7mZbk/RxI1bR1yMBoa5Z1/MjTwh4x93HRaxvk+Hdec
hsAQONDbtbcrfI/9XsEWWinZIgv8yLFFL/OoegrcoFqPIzd7Ilizpm8E/NW43uBMoZJu3xH2S38g
65bteOyVVLRAi9ffjBYG0pZwKa7w6pGZKHxTluzq6+FGWWX+oVyxvXf0SjxvTSkRGiyM3nMqXLhz
iFHn4th/upLtR+64oS3lNyvm5ttuesGWAQT9VPVXQtnDqQ289A7tJuhfmA+dpegrXjMdx8s9vzwE
NTe+uKOje1iALi3Y0GSlo7uWUMIPHCYMMFFeRS+6JGGKPsYKIZ0l1nCWMnrg3Qk6KXwuiSnEplmQ
Q8jakH8tUxQ0kbUiBj4ATMKCLK3y8GUDu5y4LtUWUwKZ9Wk4kYH0ZfSL0GXxcm7srckP1W5lMjDs
lNeTOqoKw/yOyN+4sH8bdXTrYC71CU/25PC9who8xpb1frEbJZYxChdJFnil5mjlfFrS9Fk/pZMS
OpMCm37rB/fvcJcJV3meAI1sMzeTZy7J5fiLy0JHscSmt+2kw5+AFzqIYXxjs5F50O7k3qSaS7/v
A7+lgWQLBPYAqW6NhhB8yqILf9fPn8aXIhWVOKZ2qqrLHxYFm7c4VEnUPGbpw/q0xZwZaMDucvqx
ZPHktELXNqV1MBOgUQoO+/K+7K765qp95Bm5xlSLMECpe/8S/hD4Ioht7oRF4vSv5bGb5VZQa3Cj
DBDbGoOzbPXTgOuT7dyKWQGNSiEmUIHUg8TVjS4aY13X4tbZsuiloiW8/fVTgU6ZHIQiwsRgAoyZ
rR7qKNw95Pg8aBHwDydM3pqa53owapun+JhQoV9hEANr1fpU4rSsbg3djdhkubHfH2b4Bn+gothI
CtDtCLVzrcLAEGQGZstevAocODapWL4TBZz74Euu0rKqPdTuGVA7ZoxACdWrKCdHYyXxN1+n/83d
lDP/XFQX3AWijazJaXRlpOzmJeWJLeMoGdDA1CtQ7mc/OP9zJDueZo6RG81eZQ9q2GFbLnTe73Nn
ewivvCNpNJhv+vHQv7uaRnpRSo88Hb/x+9DzofkYTURWA96L0Hanqa9yYo2eXU8JDNbidABAqQI7
7JV1NSxFSBZWX/2Nog1KFABw2HwOTHC/TqNrxFWdZRLAkF3VGeHW5F0rHsjaAkyJOd7YDJv+P327
4kkeMtYCQD9Hu2AOJwaQTZj/IEt80TBM2ASAJ58/0fjNennfgqlp70TqyvUcEEO8kPmNILYSiPx+
dc9T/1wGGd8Z5IcW9uPGQHcIqnCkVBcxcwazWF1KEY+seOSaKM5GXYrz1NArX9Ky8OuhhLN1a2hq
5qUFWSncUmZvLpLaL9R78pJNG/FeX2RcX6lP/DjNdyq9EDCEhjYju2WaTGTi+SlZ5/ZMZhoy7dQ5
xHuoAxUHoye3htalPbJA+PFqfLyO5UbFyPo/RuI+M6PSGSBZlMyK1AaUuqVxxAzD5WSP/CxDIsgI
oTAtsVpa7YqYnHPiklFCgNAiadY6ssLNLEexzVvPAacag3NHoNxEI6WcTR4C8KKzMAykp+Ac9iy/
l3KN735yHomwNBbniTK8vgCahQa5ln5AON8j3QHnWK8ULaK3M2Khhyhbui+VeyTXCpQ+1+44qu4f
QfrEo0RVDTeisAkeCkbR0LKJgn8gfbcgcIVFKXc3Nr/OiYWwxMwikMCmm0lRgrPpdqf4cl8Bm6fF
+NIY72Ex1UM8eh8FT9zFh+bDXYYAkdDHocHKv5u64Q6h4dWyHmTO7BrYgtJmrZuw/DNihWBzgHz6
zC22IQHePuAom1bM0U1lLBYs91XCSGOcH9QJXvuDoypeANycLnZWljLWdNen5zktZqoKMe2FZkrW
29G1H/RvnW7uIq3AhPi+mtPgYF5iUppxHd6BCENb/NI/i6D9JT9+kPRoncKWtCo5QxRJu63y4Hd0
rHc84FM+R68x6Qip2pC4uYvpda4ipDbUUiG2wrf0zDn61jT6zN+ht4vQZ0GJFYi2ji6qLA6ckQ3U
CYGEVwKnpFJZcYY9g0IBzfcjVVaIox1sQ1oIHoB6FasFRXeXZSV/I8FEEFpa1J0eWi+AV+8wC9qY
ZHotTYmMEc+vr6uJABp2KC8LrdRvIp2Z9bivZo9WD7/OWQhUQMmDzDG20wGPrSBz/sriWjaaX0lj
8vumXKNk9/rEKojHE6OG8Im19PLs/2vyljEAZcJQeJN+xS4DkJD1nSKOuvuWSWEGOckSGYyNhLFS
BVMEnbNFjIPj5eKspNWgLWd0ovi2oDbwNEq7TWpisg2FbIPqjOMmXI/DiQypxWsBynewwCrMiH4u
oP05JBBvt9GFeL/vVFBEEbviL76rT6jvrqVdjqxPc7tPmwhS49nHvS8TjdfDBBgHXG6aln1UgwEl
3wm+XeEjFCBSrzCIRTE9Uq3p5rjZN7nSR+jPj4IFT3GGWGyB5MdpzW8Cb+pRi02wDGEuZDE+ccQl
CKL24IzEbcD2UAMrsZsfV9AalmTNSU6o6D4H8/Tx7XuUUTEeamZ7wGdR6q8NpbjvRqFqzFGejOOO
tOanMGoas+sSeELWUeqz95jEletI7YTTjFrVfy96qrOJWB3E+YUyrcn/YVApiPK+4qHT200qbRl4
1K6HzQG1K3uYK25Van2dws6CTUAL55T00NsrMse4XnKD0p+CZKAHHEpkYBAzsy0WpfnXE5lgBdH8
KGwKQsfCscRw+zE2j0GtCdxBfeWKM9QHqIsD4q50wfWLo9eJfLzJZGXChm1+cszFS/gtLCHCtBNi
Fe7Q/re6eB/7HDtcu5NCtmbzeoUXKfyss9Rwvj4Ou0uuMxEcEMmPlLnx2C82p4XZfyB4a4D4pLwp
hD6a+vmyjpmtK13uzueNQivQiof4YBINFkpjCcB+K2AfrPz7kHQiD6XIWqGJ3Da2eXqNzpYXOKHM
K4RRN4ntoc3l5g1cRH0kG99N67MBRZyUswMUQwnBDCb2KDXNQjj4iz7x67V+4SUj4TeDj24dN8/g
8CLVzj1m26ZITsbOI5Jilg45veeZ0f1zgZMdXjQG76jN0rIO4GlpUEyc7aUPhEleGpDtFfacnZIa
XB6jmdVAupl3dVtjslb2F0WU4j4C+tUer4zvx4tHVhBK99Tx10hazBNJ7akrrK5v/8SD0fmrAjT/
KMCNJMW4PqaSHLY2PtNy0CvOI1W2MXlcmsnMzAIVM73iGdko8b8uGhyV5g/R84okz1dM0lYOaJ5W
qBm+y0rrJm+81VbBhc1VgElBKnvfKYC9gw46RXpTxLn7xjbhKpopNuWviuqCgKVDWggXPu4mwRpU
mMbYU+GIOHiUuQPc/56Y4G3yo5PZ3434j/fjXsfCHlOGlJBg774re+SZlUho2x+ygZ8Z9oExyrYk
Y1s58KSha/035rk1um040KsfmrJtzIK14FFhIUbE1F3gHuiKuGN75DZyg0K09uoldsOJZ+Ztn6A8
xsIFMPRE1f1IwGovofr25KBwRpQ2KcMmdrlUuQDztKc+9Q5SFuwjmGQVFPZY6Wcv/XxG9NRKCXuW
u0ovK4M0VWsf72Rw6w/Y+E4nIMZLr9VYjk88ALCjFpLloTWyW8y4G+5ozjxfvLZEP1zlMymwT+Sa
cJxxZMqS/wKA3rXcc0O2VhAxpos6NWnhi1bpFXFUPGUmRyZ/QuKOb3HLZgoZLYsuJc0WAsvUkiep
RcP9AzkL89RliIgxgb8sLXahXEGVNBI53JDaPSWZJ8cUqfrIAlXELH/5bzfAxFgkeH5cxZQqO0Q/
eWmTKzZsreoYStOtWP5VBxV/Jov0krK/3rAoQej6R+lZA4carxLxLeDif7WxUquYquAmxpWkw7Kv
yCriBeSUduaZvtWCGNPfFZnq3Ekd/0K++7NojzsOcBhsaW4MI8m5dOqinpEQVMLUNbDcYBz0sHPT
G9BNJ/NvNOrhlFN4sUHzhtI9dcElHWVbJ40Gu38LUSeGdUYiC2u+0bbTUie7yfuhN4Yvhyq6F+Uj
5Ulvob7+jtDQ0tfZf4j3dea/LnLGjQfMjIgmXOg1949LbE574gZm7QPRy8ghhiMdRQ+v6EV683hw
6+Au5YshmnC55VE+KcA29OAvTXlLGKlquN0TaJMgmLXJo+gXOoX4NFHBXAP0LEU2LYVfRZ39SJrG
8RTHDMYa7fOwmRgxXq3ZlBaOYdO6l0OOKG8gewspVATIBZwLNMHw5kujDzlz/CaMlAtHIs/ZxIBG
AXgbbCFt4izUQT5XybCi9FhRz5l8Mp0q07EpQcazszK8R9g1MHr3LvDYQGZf2PV0pg7uW71f4U1L
yl0u0W29Mqx0qW+KgJI9PYvbWNEpPL1yy9EhpWZnmLVTQVfzidDc9XvyhgGKdRN0YFkNXByv+HoU
M4U3/wmV1X9FczOjatY9QcDjdzF58OuFMKCjyJvMIfhfscSdwhoIvZqXbWUrA8Pm/7fbx85dxlYx
a9v01xzD63eeBMp+2Ep5FwHNk6NAssJ1x14FFUkb/Gfq7hBUaVfJhi38dQDvn8tzN0V1H5m5L5LS
UcQygZHpfgewEC5PeRxj4q3Muu1zzegQrYj96oq7BtJSoLvJf3wnvecMVGQq4JnZdGXPgRFlxtGU
Lw8ZpV56VRpWeaoA8JZqWqKNAbR7GUnRF3zIuFS8orgteVw5tHKbaDprEs8q4KaiYFBc76KIh/jt
V0DVeEX2eCCZc3jUPFDQReOn92242bWilR7idqygLaPO7HGIo1YvpsCfq7KBtOiZsq8bSeHXzzrY
qhm947Lx63BLbwxkFJppOmE4mayRHAiRPP2yf/8go3RqLF440NN4pBKHb2uumdp3HSW/UntTaxvn
eN3C2sDezntlsAbMrfKD1cSOaDDpXcnbqlKlr1QsPJnAMJPUrftysRxf412/ew1SRNPONHkqFDvT
0wLhyuqbWcJG6rg96UA+UlhKtgcqgZLIuB59KXNXVQdle81Q42+tKcbA1d8jvS1vzTrXumjjOjxZ
R6yfcXa8iVYG7R24QWhtiusIof7P6Ca4bLs1/q2CBI2DCWoFe+ld4SAxZVVILWF5cG1zo3uyQQN+
oSdLBlQkDT2uDTGrdV6kC+1jOYVPnojS6CvZgZ1MOlNezTizQqaTzjvw/+1SF3S9PfQPE9tnrDid
CrAeJed1yzfLJmJWjbXpvCUblyEAVc1TUz+i2ub8JfPBOgrvwZcZi1Ie4MoXjrVcu0TasI9DAbvh
pbs8e40movnLb5WAOtwSYmoKm7za1N7GkkUrp82rt1RivOqomMzQQ+w21ySAUiW2cFn/XjY7cPVS
k/QlmFT0soISMRlG+KzqtwfqCMDu7+pkhCvT+Ra0wU6/u6Vx8JIeUEw7jl7BNrNvjdqrtt7K8LAL
dLbExsL2buVXAfVkYj0MZortv16muUiGUOclV/79RutleF0qD3XXCJmlejoWtGM64aXSXIPfYzcg
sflIVJCnx8ruR7rwLkKA+zWH3edHKS3c4a64oQibgJGLEGlqcFMvaKb2IH9FGEgV1g9f9EsnxLKs
NxHerCy2Sy0cb3fsLYGqrq2NkNdx9I5sz0Ft/OO0FXDHcf1jhopwLe8b9u70hLamQip74P/sL89v
4cv4ODMgzBnlf2G/oOzZyzTYIVYg8qPiN+o1pDtrQ2UvtPMB3S/P7e2VunMgOZLQ+cjZu8s6ST0X
ffNsfnTHGpc0L2Votvr3UQI6mCR5wAhG97fZx7Dkq2G5UUdc/+6T/FCpmTEKtRo6SCikXR1IMxIn
ASSR5tCD4dvT/ClN1NElnMDdKfUgs+ZzFII8XjZEQVDfLfBOuR+QkiHejNimTZ0kyIo/aYzPPoK0
xHp8EQf/U++0f3aTz4xdSws7FpJFfl4QKAuzMUYtZUcXH3hzC5jBMA0K1PSzpVqjB464MSogvvtm
GiFPA1kKLNycDPjfZo3IOFgJYlrQzF5AbSKUsGEfZlNr9/2LMwTyG5AZYyvjYijaizACA6fckE2e
SBTrQiAauyTJnxOLSolVwvBEXoBfbsQu51lAnxcR4WZQm5OJfD4P+5dZCPj+Le3lDHaObp/A9y4d
tAJuqKfqCQ/il4Mk7E6ALVcs/R0Ys285QavBptIR5LC4bODH9RkZvPTbpKOKIJb4q+tpajGDGoB9
u0INAbpGbUKzYWT3Lj8Dbf10EGCZ7dOhK3tjkBFldGrQA9fozPvpzLR2gEjZgPNdK0u1mYUsGTj3
xorSGWMSh+tp4UVfD9garr+y7zrpw2xSxjDt8xxqkRFdu5q/TMv1wpqevkZd+ySvQhGn7jCnMBc/
/LAreahNjAEhIgXllEPU4Kh2hYiQcSeLbOhaA5iWzF08zt2uVLWbwYYGFhvWB2rwRBTop+0fn2qL
XzxPJo9xpsf9a2IxJHDtlcfJAOG09Q+2ge7Lzzn0j/GgbX8uJGz+v/EoIincMqUv9g2zCHBOBPbo
/hw9fbxywFL+hbPrlgtxqmJI+huMgNyUcZH56/3yaDzDbNZ2mPiBRGPiO+x9rTdufz7FjxcaLJzQ
G4ZZC+DVkJ8/S7E7kuN6FRrJgMEeY+IMdxrJAgDb+yqUjJjciPgkZdl0rK67cEMaOv2iSSjlONFU
HXn6fqB6DGmPBiN+bthRUxqo4n0xiP1nKZ2DVSnKOrF8Imi9lXnxrVCAwzRFh8kKzS+Yj5/3NS4A
9Z5+kDEQIZYfXV3KU0+8nIoJVHsEVOnNYhcyqITZ9He8ejpPnKmmARCcyoYX44B6GTsr2bn3PLym
v8r0eeJHkEeb+TZ2aqh+5OBPUFMsUdYW019o+YwXYx4pnPNC1hFnZsGJYXHFna3Y7VnGiMRvLt6a
2tbPM8UOltF1z0ZNRLWUVGsrQ2lF5tfeQkQQPZv+VppiGSXVgHgKYaZi9jxNdFXxXGHwtNpgLEvI
gN3KBoAMKlNJLmoE4v/0KYwlF5/AawwCfnibKk8rDbku63WU4O12zDeor8DUjI+CuqIJ63VA87Qi
yThjB15kwbICD9E5cLN8ltx7Fw6DgTS1eQbLuxWsk7eLTWk6dsqUEbj1Mv5MpXPXSFcIhoD8Rcub
3UB+HdRghTgqxNXvCDq5QFr9Jm6lbTqTK9/NAQipNFVmY7l8kH2nTDm0MGdyiTkQkL4NPq9ZNPHb
45r5qA0MpY4BB9VF2Zo8nUVIZ7fbt8Z8BJkHupMpUKggsn8lkraFN2z37BjH65NnCNfadzjytae7
fbNbj7ym0+YuY/Vhwo93kMkau8QNcKeUbg/9tVt+x1HVl6LK48uAmCYj7lgAnrUzOxb1br9nps9I
ZKVOQKJlcMjgtUV1bnivB4gLTon+13KNd5mNnh+EJ8ukzIcI4wXCg0f3cvK7E3kl6bv+fGfOEpWp
EkbRdpcWhCCKcRHoHHgcEBiaWRE2mXgY46CYN+c74wTJQxdQ5em5arHwgM6nWHWFhn3X7FeR2Cvk
hLDbfaMKnWNV5d6SE+dEf4ryKUcbSYHP5ZgpKd6hdj9SaBrN8G/kk/7NeE3gY3XlKhUdhXUr57sD
EYaIw3Z2ckPYRtqCOqcAgZjxDCElTz4GX6NcVxGuEBPFec4P/qn4oKsMJCWzRNLQPzKP06+Vqs2W
PAYpWo8TRbjPUO5z1JwkGlVQFuFA1qsqAfgwia44fuNz8q2svYH/YqfSQQmd+WnTeyDoRX9NieVf
O0aw9C7IWjD41sQCx/ToS/GKtMg5N7/SNfUQoSheXpr0ES8UU5UQKiNcWBvL60/9pTCpeybyjBcb
BqyL2URtq50vOF4UoWMdyfwdUJAMT7hvcO55yjG3BvnrngMWezAAxn8EBzTSADTxrrUd/2qtIKw3
Tkj3kXGtqCdXGUsdXJUkZMZZ7vGutUlnH/I28+bqVxlk9AI+uyX2TIhNILh//ir17eIA/nK8iSPc
BpZTzZ0jVl3HCE5EwW+1OXrSW4gLB25BUrWmjqJqyPXVsodRQBaqcEXqkpgJFijSd/93Q8cACidO
K89IsUj3hNTFLDK/KjH0No2/7ERlrcotsDCBko8kxjFskG4k6d5NgQpsCivF9g7+urWS/FP32hmR
0u5lXtVt6dGiMh/PdqTzNif1bW2dMcyYvnmdVLo1ASbyKPLXieuLpj8+as4aau50xjB9+yfEMZMm
RRFWb17crpQ19xV+8OAHn5Zm+xQrrXkywSbgJK8eigXYhEL61IDMYAPus+IP/7kP7plewJOSn9Gy
5Hu0RDuGRX/0Tiqo5PdNo9cTWwIy3T+Ph8nKEwa36yYjlc4T1ndUY7ubedXiXF76x8dPZwlxNdmn
5PqacoJgfmeX5fnLl2bCfaI+Ngj8p1tmLertndsOE7b0dNT3wG1G+CzoAaKvCFO7aCZGysFzotXF
g4h+jDcS2CWqXJWe3eS7D8NXG0XhpG0WwyGRNMzNbViJkDuMoEDOu3cE1UD6shzJsscEdRg3B2AL
mBuiT39i1RH7NYwmbmD/33D2YyJvKlgpn0jRyETR1nF/fyc09rSaAMtcsJWAz+7Pzwt+B9ka9z74
7FCp64f/rDs0Azgl70oayOk3X4Rhp3aEozzu+NY9YAtTqcIiGW6n1eKJcaqXKRAG6pC397PDfNCQ
qkbMEzX5t9OuSQuU8im0umfin43Hba9Tu3WU5XLYGKO2c50EjINEvJZ9JOl6gLL2CXICP7A6PeUw
HKd+dwar6G0FPKJTY6qsoaRfTwMPBlbaZ4Y5/VBLaYVrvg3r+Hl1xYjmPZ7bWEV9eNKndUTyaU/e
VqRKZqzCKmm/Hj+aesJo1vImoKNjSX4Q2scsvD1MXNBQ2AbPo9WDLz2EOQvD3r6IhtwqYdrRs633
betTJ3fLzPHJixQQvk/VHL5HfAm4kT6OeZezuteKB4ENhA9dYZ5WtVQkT4elsTTW6W7mYFB7+RmP
FK7OBvGVamgIhJcsmf3BlnFeLEoVei9yzoNAt6ZyWskm6L2GRWJwjz2e/3PNrPiKWrqDUGh//SnN
rtYv/ErSjjihCw94iq/jlYWAWlpoGkYz+MBq179RCV7lzCgzghT697ZAdPD4+n5oHkA38lMpfdsf
D5hlIU0ifBquQchNkfPVp759gJllxwcOmEGSoIsEHTZ36Z2PEX5gXXQFNmdHfZn8KqLB+IBcPq8p
D9o5u76yc9hvFRIoCKtPUfmLwAdV3O8W1gL1ih0cDjILTAycAWILw3MXGt71/YfitM6nG33ZwAYW
yZOI7gXFc6e2zpNFe+t0uiz8JhnMkQ8Zyn63H8myomvgo7ure9YvkSS3YTkWsaT1Dz3DGaqoyXvf
tOdYXXm/R5m4AiIO26WfXTROPLJMwBkW8woDcD7JDJB/+D2chMtBmaiLbB++dPgLdWU49rIOLe4R
oGpyvSTs2Deb/dpcdUo4y2QsRGQJFimc9GXJiHG3Ah2NHXXK4qjCiAHpQDw1Uc0+PzHnq0sIefee
n3ERbfBjZP86fL4au3fe8dStkcpQCgqRMCNYu0Xg0YsOiRdaLxYRP2ZMsttCPUOjDBunNPj3DCGv
AMaWVWX26s+/8sgkQsnV1ntBHZdl8TN0AyFKdLB9CFvAftxQQxrGDDeYY0VtBep19ucbqmlx3FyF
sq6/JifPmBqXltlF0VaF2dU/Li+NxSK1g9vvWUaBWr8kiFGYhsMhgqp6RmKWaxYRIINl8hTGZYL3
Gsv7oJnqkyGLvfWedbTw7xE1KK9Xf2tamE8gN+1led86B0DZ63lVtiYFrtouk8Gsxac8HBofEKCC
b0NO6MQsRggPEyRvL/QA9uV6gI66XsSz4EospmLX/f8la6drbxj9OLD72ub1g7N7/I11ETTi8J+K
q5xvG90QkUG9Kgnsp+EM/6bSxng3b79ypI9B/u5OySXQBE3ZDJ1mpw1Nw48RgcmDpvMP856mWZXW
stTx/HQBKHe4bx3Tvv1XmdUOdA8GN/6D2VBt/FYSFK/zP5CnFdlFmVg6t3CKx3NysGr84hMKuS1r
ZABUlhgWMS2ejPG8AxeK3nX5a0OzdlG5bn7H/xNsu26jUplywsg6Awkf6pB2/cY0oxvV3jR2zlzY
0JEkRvIrFdnoSm+4/p6Dj4j0Q1HRNOgIsGMEgZHNhTprk7FJLar6YjxKtLb755ufj6OJs0G163HG
QYtQnoO44/7mOyoJ10KG13JfFaEtsM0cs4KVo9/OR170nmv6pVhOe5yy9/I5d4mxTCNxBeRKrEyL
2orkehc808WaoXBO/13xPFeo5Ivs0fgNDTxjPVinuyNwKApcdcToODSBfJnokoRuFknm2oWzG6sn
1yYpdTlLRObT2/Cp/SdZozaQLuPOTTFBZqvarXnT1+lngggmpx0vZsHe8nqkr4THBvbulgKS6QI1
rAitNbFuyKtf5Pvy5BrEn0YVZYuaC6Wewn2cpww42UeG9vfZSzXYUkQ2cKRLL60nYWBBi1WOIqW9
C3e9u2p0SDxn+mQSkb7HW27tzHvSs1U2xWLzkpzNBy6gIaX20d/asQ0voezAmxURd3lzwNWnnqVg
c6zBWAm5lEuTFWv/g1BQL6mgFWPL115mD5gz73OrMhn1z2XIj2xTe4CZwdSr4hc4KCDkbBKJJ56M
nzr5pOoArfK4ljmRazPUO0KufHeQruqjBlbeyRvby2ysFwvYGnb7OgMQX/WLLvi9CT0Vo4IzDqsL
kdJwZI5cFMH7tTPZ7aMDf+1FvEPtOJo1TS7CitQuQytgoXCPSh3LII84iBDvDAQCgwQ2oL1hViwf
lv8kvD36k5DpzmgWw1iuqCbGbXWLuaRh6Zok1cBebmirIwmA21AzrtK+bRNb0WApVYGPbsw1hdfX
+X2cLlXUZ+bNB1xUZXVDSlQZdaMheuuOXwc+N4dG8mLyFh1MFZNWSJRTnAEUQIIqO0XkLDCy/B2W
R1bt+cvG/sY6GIA6+pFad0JZPkGRIqn/0jv756LHdtxN6uuzsotCEtWKUpbTTm3VjcbXPShoUNUc
YwT8Ws3RdTb0KbsVm23cWvNe4z/FQq6Vcy0F+sYIGAKtviNCIOsZruU0NJlz6m8TIH4L7ZJVqiMt
Dd/JYKK/7MRKE94TdTWyBzErFfGpYqCXTzobuajDx/Oj3qmw2cUS+9y7n8K3CqfCBwc+3ZuIiCBC
Ab6Nsd7PbyiA6xkzzEOgqC5PdjqkSNrH1Al3w+GgKXe/lalz0ozcNrPaGqNo7rrgui6H7NakHeFQ
BKnE6U8paWuzT6zhmRVt2RujjLGErsyFJ3ZHrVWK66NqbtjKN9XoMIyDRYM4LnX0nlBvXCD1j+t4
2qWE4m7mz2nWVnCVALkGFq7UAPb1lMHHGCGnNmJwyvAwHo2PXpQSgM3rz6gX/KVbXfusqRjMs0BC
CBlqkTmyh6uYzhcN7Eh1889kg0JDSxCejcBn5PRGsaWgIamvvQwapFKl1tw+ryjVBbeh2fosooiy
n7ulrtbIMyrEpZV+H+1H96aF2Mkw08o3gnCI9b0aC6DrDApYdNyaeMRVc2oFP0kdFk9MtoFC/xLh
R04WiPVyaDklnm2NYljyHZW5jTL5cJDzVdk6y5whTuHfbYgVc/w/+UgM0burdBLYp58chM3a7glK
8uvczQGkIENZHq3XpTKHBx6cU7WdZSSPKBGRdaXLcX+Mc6Jn5uz4r/chYk9Vk3ICLx7hERrioYkt
ga08+/cL0p7quLe4NwGT+qo49HsUOHOh9ULcorpWiHS3chtNjIY0oDeK1vbvJPVgDGTRoNq90h5t
BG859alZGHNHAUphRyq5485cqs+0bYReSq+RE79IUhV7OBssRCbfrv3S1hHWzIvdvRMEPL0Zq/Pj
da6xXy0Q51hQmfQW8WVuJ21NjkGGuuBA0n8U8jrjStLLn6sDpb0bjJDt5OoG5kmWKbeKVcteQntQ
RW5mO1WFNmMPS1Tx2M4kaN3FoTektdPj9cq//2YvoGnWUW9gPZ1yn7rtBZyjlIHRgnP5DQy/Kcr/
uC2BejVr2MyQ77SRYByePMngzyX+x79hU5VIuFLDw00Nr54U/ZchaRuzCBvK1j/xORXXquMgGdyI
R68Dd8lrCq6oI9B6eKA/+I3cI8CJGWQMNrdxqgkg4Fe/tW9A5DeUiHKeXI3L/u2wDTpAabh1moTH
ge/lb12JRXK3ftUGsuvUK5Q5HXhKyvBOpFXVZB0A7F+uLmzIwBf48v95o9TtJnzMzfP/mzkgYWiQ
kDWEVXJ2lT7LKp9B/vXvROHb3pYEcEq1NtEtdFa/2rusKfzDNKPQphOj3P87DgzL5e4SURh6sNPu
ibmZ8pusLViqEN31x+u2LEWFDbaMxbd8/Rq5aesXmfRW1Ijf3ebugGd89HVoHUp0QpI3zHDxharq
IYf4Qjl21D86qV6w93pIqmHikBaACpyiL6AMPHFRkq3KJYGEK+Uzzb31gBwE97a7ByxKX5Tz1LUi
aegiv+AqZRmMXIXGusTvNQktOF7uoGmNYyaeBxUue6ClvM3qKr23OX6+5ldZhol/zhTTpldMEebK
nUsAyFaKEk1RNPSb2ieoKmo6iF3N+2LTtTDzbpWFeKvDktlV9xnKHdZEQm81BdUetWTzEiZMaYuy
MvMcXsrK6qCusQipCbSP1fRxeNLvtXdRgV8ExyBw4uc/RoXfxU+38ISuA5RWgn/7ZGC7Qf56Tv5w
+Cstgis+VXEm2Jq3A5Wmza1dbXAV0uVfxtMoCh8t5cQ6v7gPQ3qGxKnZNxyleZW3jGYLtc30j4J3
6A/z4P38XaZR73JzmxLzCUu8I7pnHRJv+lnzDal4sZ4Z6rTdhUHCmqPHBxwKVZz0RcL8vVFNLuM4
3Xy+NvFod7LqGLaFq7FzjPrabHGsaNVGmIluRegnfsDsb5A/ozvMQtFaaVS5erV2epCnoYoUs5Jt
qBVtXas2kJgN9GpSnCajTiMeXOJDdEAYydallqTYChSc6ei0j9KJyIBRqGcHiSlb4p1aYRdzhydn
6h/fHpU506DukWdLojnuYC2LMzlZGpOdoF7NWmJ+4y1Lad8qGOGB3IDOFw+Wvlhq9HILcGg8yx4+
HhMuHlpzlW+BSWa+P2M2eSXjRxldk/aPzpMrx6rRuRY3lXyBOymN1GfiZDvPmIbkWUOaescWz0Wr
sJCnSBpYM4Nt82bEZ2FmYXkn15CDsGQZiTBsfCZLbqPRpKN1mZPPIhZPSMaPEVc6JdNTEevHRmfw
aL3fI8gTj2N3fERmBMpBE/B9qdplfbneH7mAcYwKU7LFcevN6Xk39ipzjInvnl5zIE9Gkvkv00tw
6TbyTE2oYit3rDKnJsoGlqiQthPEUAaAyYxFhNaPazTnfmoE3uSPaDJZVGAd9hVkiEKraIKbgvVw
JKJfhwtO8hs+qfWmOtLyMDrDFiUs3dj45K5Jjz2Pim67lj4IHdby3b+Lwbljp1kHNMLiVnZTkoMv
31T8jLpw37Nskro5a4CBM+YrBpOMe7WeLTHxxEaAyMRNkEDXBNPGfxUBdrl14vdxYxcaZT5Hk1cy
RlQ88wsgksMlgKA0yDXCAzt5emt4EVFaBr9zQvgqkHhsJ2bTAn5nyUyYDFniMEm71P7cfCn+MUV1
ryhARlrrQBs8qiumnW0ssRzS7zPG/cZENVIFbzeZkC0ui+sLXst5ouJ+rnDNsCpICkS5w8Nc6QnU
IAIEr4hOrmzpjH0T+l0N5KV4jEZcf7JB37z86+bNiBqlVF+U0ejRHT9+ZbqSfhGPpfmVbYCKfBtL
tClZuOkLDp+P/GHzxvqsrZhQPHHJMn4ZznXosqZ/eZYu5gNks6tvK6BR7X9mQFO2Lkc9R+PLJvCm
cqOjpXMUDvF53MmYGeH/tA0hV2rizF149k+QP3VkPMQyF7GMXY96Mz4Z+6q3pyW3m79m7mjZpOV3
VOBt4CYVbRo59QTKp7D30WLJSuWS2AdGnIsIhAuLIMw7lViHGF2GaNw6dUME0ge289cVLmbUVVK7
rQ7zDheAP85ludVmrF3IMoSw30UxgETXh+ohgx9RD9kDMKsYr8Hv4rnuqajqZxPDbZVo4fMLd8Tg
i9MPuUsYiTuohAtbgUgZcxi2j3ri7kQNGjqlrCeygL20Uy8TGlREOU3k01+lk3WMk8uAzm298/dK
GcjxR/vYaIjCuPbQDWlDRZCKgW4iqUmP4jqzLzsurpglPttDDKALR7bram8QHfpY2dll0rA3ruAY
paaejOhqpXNjGHvHnRIwPfHLtY+q2UXMxpt6nlcF4Q2NQnKG2JAzsNjTph0Cd8l87OKJKLk+K0+p
L8RbahZCqvgeqqmk9qXzE46UEQWWM8yqD6YmfMmwjtw4YVp4RxEmFezJqRyxvUCmRYbzzZqPawEW
P4tGE6FGIhxfO29I+21Sq+20JnY5trSqGA8C3hhTiHTvd+/kqUGltvs4UIG4fHLli15Eyamqywur
Xz4HOdIVp5/lc14xfJAYeOj5HPEwmfRKBq8bBlnRc5iiBFbHmks4V+sjoIw9gY3+2o6j2aYOCtL4
AbE5s2j5wQTeG28zMfpGMAchnP/SbSPjCBIPszdwVSQEDFGzMedL42mw3EVz25UNyo7O+O5JuFS0
HsDPhIY4UmB1si5chrn4nrOrFU51xgHbetvXBYKOVDhIAj1eKaNiJlM+1uZovRTu19WJucFcvQEo
muDbBTMJKoh7yK01BeP3uUT+ZDNOMtfxnlk59empu1LrC9Gi2gIn7+altlHomy3j3n198PBGyQYi
Kp9FvPZ1iXD2/6oWn68Hr37GsGV+sB9Q2i8nm7bVy3PGXBo7rmkxbnxkV6edj04hZ1eOl46+xfLa
17LPzO4PXufWg9eAZki7UKXv5FwWTSKUaBRyr+sG/Y2dL9HmWjZLuSz8u5hAYIcZnKXubgo0Lrr6
07nAFyvzHJkPCBocRGV4NBYOH7qzM88RtHuD6/RW/qGV6pYOlomLq/pT4eFeacdxqqzzFK52ZcKh
/w08JxIPNXsVLmRtbE8t3/fFoACBmILYv0vBQse1pM7j7urOekDS4qG5OUEZyFNwP4A6Of92lm11
LTb1TcL9BovwmJ43O4IjJebhKquesodO4e5S1vdOxTQpyWVGZXIVa46vN2huclKPb5t1DIVz7fcf
Qy1dbC84+87xzVj7TlZaezQAcN5Dw5Y44hPNyRkYOQ7SvD686f54Dgw4VlfyhrkT/mzCWCT/++9c
T8KSDRqATdXUlPTBAFhjMnEjjzQpviKd9X8ByMMkk29W8VaO7jYAFC8+eCUS++oHC08DRF/DR9TW
b16thT4RHpxThKSMOT1mVDUqCAE3osHPyZZNbuW9sjsKu019RrmKQoj89Zin5wLzI0VJPqSQIAJ4
+UQuMX4O0J+6K91306EhbOkIQqEReEAA+HU09DgJYb9HbEaz1gdbReoFiTWnfz3ANGeqpBNRRp4J
w+vfPu5RzWO9VLLZiZR1br6Iq95OGRkNAm1FBGYrLOH4qu4ryFOSzE1QTGeY3zRc9PfNrW3aMc3T
yQTFKU0BWbQZZfSELqs6IUQ4BonjVkEbaCTLarsEwtHJ5/lua/TfommW841MmOU2v9sO4DxoZeA5
maQD6g4s21G532/zoG+dT7IdC7yt+dcEsSadvN/Nz4tqzhKdR6LYDW7ZEobTQLhNbgYs+utNWdBU
SOb8zIPgvbug/58WRIiNwfH1tAv+Vjlkbv+7/SUud5b0rPDdQPCw+2OQ+YPHo0ZCkVJPcLy1fh4o
SU/daOpR0vmLhHoxzgLtBbXGZa3DN9hmkVgyd0VAH9yCD6fWC0fLj0YDP+0uPu/j9K7wPuP4+ybA
+ejIU6dJgLnj6HJlVj1RBp2hQXhQmx/+v/HQVtOvIL/iQIWG4UcELaLlWkmAzJWbtia0MwXsq20Y
sm4oXLVyY+c5zDeiY7VAznOjPqMXjD+C6A0qt6WrL8IIASYSqUSRhCkzeQalhQqLgf6d0tdIkLuO
Z0geonXiYMpHJDoQAidt3iQPILYyMhTMkEDodncLAu5DwrBpBhavIL+NS8QKpvCw8nhCKOyrQhvi
ffB0M+lv8c2dQodDSxUuTvNmBf20CBuW1/699QgtQaJ8TnOSN2I2WUE3woaSStxSXy7kB5z3nm5i
GAoiJrkY0N8bz33Jf335V5AtG9HnN48JfNtA5ndRmD7ti69ADyvJirX7TvUWPnINtGTMVwxHheyd
6CMbayx7q3dn/3syxr5JtvCZ6kaYYMvFsd/uHbWCmQVXv40M+9Q7okkQy5JIDnH6tCP+4grupK0J
hFjq0ihuC/yQPJ2QDIVX/XpwsAIXEfaXHisXT4iozrjU0mR56ioHEdxA1AA81l83kyG/ycPDTRhJ
5lgkJaGKXhMRZ3o9tZ7JgKblwpOUsYBBj6Rt/O1RNFo/UiLi19QNeHut6vhY+ubApnE1yDWIJgof
njU8e7Af9tybs3Qzk+F0cmgrTcIrVKYe5X2mgNdtyAJ8KScT+Vkqi7JwO9hPgT2fc+DAXRlIcaM0
Aghxlxsak4TCsxkD8xji1bWT5tteNE/VGchf7MPUOBcaz6vc2qLZe5CVqJ2H3n/u05LZbPlO/xZn
z4b/wMZVVvNxdCoMBTWADGHoG19FIii7z8WTZZz2O+YTWlf5darDp3AcbbTqML4l5xvREyuZlvt1
CNw92ScfUIh3ufpLJRRqslVuesfb5JF8QR9J9kLiq28ysqfgoNaAS3N4Ey9c5bgt+mCw6i1ak957
vWGHkgSgRUVAliCxc3zXa3T1dOtpqNW1eTyxrcGWj3YKvJsW+BbjQxWeol7SEfDhFsvnYuyTyxK0
7Yx1zJZGrLNIgOeeh/bwnivFMa6yINnKbOCst+gcq46bgBghjZf3gehIQpGQe0zRfX9+yFsrkmOE
wC2Au8JBK5i4w6qCO7VUaPLFpLe9G5+BeedLoMXqhwU1gS4zOdS/fJLppsc/50BiBHod8OSqgkbW
rXqtJtWKA3EJ6QcekBvx/Li0v08SccdbIokoGSxX40xQdLnV872NISep64Cg93fsmEzweXAIC07z
yIVMukSHhCmN8ASR9GRZXMJ0qA27YzxE6RUR6E7ZXo2Dz5TB67cr66p/QpieLwapjtwhkDRXnMwN
/x16W9eNjCE9hw6MLSsMzM/2SAVtEy+x1y9AB5ld+FN4/7RKJqFIfRaaB34DYjZKt8BPs1W2vJi2
McJ++IyVZn3ZYADyZQVFu9fB5NpCMIOcEPEuIkD/MH7w59jgOeol4VvdwgWUExuRyc2VWetNz4ST
O6gET8qBI++X02P4KxxGRV4/ctUWKnSKfPBxRdt1ZkFcmQHHEIFn1CuVDC0ASW73p8y44oTrvIqV
+yKxeHI2kY9kPJbkPKMwG6v6TD1W/oBTVZFBTXamoGKCO8FM3abgEMQ/0txeL2Y2UXsWvLY7O+Rc
kf35zpZzBCDqF1mSAnvPioySzIT3RR8rt0YO/HbfffWZt8dj9QWPJ63mz9LXbCsvS6AjiBv+JmiD
Ozfa56O5kGWbovjy0tojXFNYRMQtNTf5UodXAPVzDioni3fufdbERBZGVqiXPuJKLpGQmtYub/b7
gCi1pSgIM83X5WhAGsYtpfr0RJCQDxPtz5/rlhXDwau6XovPAb0iV4bmLr/+oCWufdNj7mv4yJij
+21/appim3rt0IcM/6C6aQb7/yjRSv5sjHmSMMNfi40/j2OU9eJQb40hyuseFfTC0rwlvRRi0XkN
5mnePTMcSvWHxE3gIdJqMOR29PZQxf+N1K2qd1ET9zQQaaNjuGVEv/Q1Bim8zVWsssdCbDv/VFKL
ufWsn+SIrDnnhlBqkCjGol3vNzK+zqAb8+C6EciTXeHJX9YiRmKi4AugtT1BOz94hVCpcAPfb3mN
wCbGP2fr8q3RSPwdSReUKax0jmtud6T3CRbHb63UdUcjFPReazQh4cNHauO35gZ2sdAx9/auooCY
iNIzFEXEuH/hJCJipSiwNdcO9VUfA+fr79RdUwXwaVEptshbbKW1A8QJ3LIRq4jb/igp1S+x5Be/
Es36CTsR6KTv+xBtjRI6CRr8dQttZSOeFs1L71rtbY2nAvhLCDOc/A+yOEET0tzOFkXpqhDHZpCd
XcNSKAm2cL0Zvc+HcHmMzdYse6Yo/d9lWTLF8cvbm69eOZ1dqP+sqr+yyQJZjNZ4TqCNlw4zRpU1
npwUgLoFN32OWmDl/SS6sWAukDnMj3+kpZ+BMGljE+Sv713Dq4dqOy8J+Y9G/xH7/XIxkTdJbTav
EUdUZOcoHzVvsHfHgG+e/Fx9AhFc1ZOnaCfa4M4NMQeHBCBCQfQ2CLH9VkKtxdYHc4wzkJgUeSRS
lbngJMI1dLB0R/JF38XS38cXMCyWLSEoQAwEIH34V5J2WKt5BLA6fp5qO993MFprleLX84Uyj9ki
5FBBaJZiDAccGSS1Y3gfMFNQpkMXzQEDmQBTSIuWILyhlCJrgI6bKNgLuizHnvT/fS3o0IwKbiQT
DsDxFNv8tcq4/YVmEfA1QMjQL4f0FnHgEmsY2NB3G+Uni8dJomY91XRIBCxj1dhDVuTDwjNkpL1D
s/iF3wkQHRBpeLhJRXfUhIjIvljP9T4bb59sEi+bF49pvbHl5PBCc6bOtqhri+ObGpwNLB4Sr/8k
bquAiJgfyWSjm4MpIXqaVDsTr87TUoHXyPnW5OUCI1xFUJruXdQgS/ifEoJkaUIKDGbF6xomQLSV
QIC9IA8WlCsn8Grov8MJr7UxazcElcKM7xMQtgELmNMpxJB6xycFVURsDFf37zL7fwp5iteCjMZD
ykMelIeEAQkCZK1uWEEMuJDUnRlZlIOArBiw2PzGiDa/csEEFuwQUxx4pVOWA+sS9nHE1eamTSXA
r0aS2zn4pWWdfrm6Y3pBy0WC2xVYtBWSsXAM1AlGrZA8RotYBwGFbD10fbmvA5F0dOyToI+WCns/
hT2mi7g6CQ0SeE2pMsg8bgizk287Rvf3JRbfUnKt1T3p87ltwJg/H/oZjJNXlrTvYYRDCLA+d4l0
H2nYxSRxSiFNxBFakP8vrO9M1J9fVLe+QFBOYz1su4ZWe7tKKnF2AA2qX2rdDqF3TE5AdhC8uObe
ObK7M2bUnMA5sQ6F23vTyB5ThD6pQ0sU4bt3GXt0eew9YAhp2+SLIkmuxzLgwoIeLEW21AE0Fho+
Dp11Vg8VParbaACRc579rt1J3dVwVDGt1kggftSGs9FkKvmlTQU/Ns4LFOaC4nZtzDpGOVjDaKlr
OGyfr53XkGebzQ9ge5S+UrHAVWIo0EI61bThO6g4yzK1LOLqrVYl1DENIoudYCvvmRvXrYrWNO92
nSqKvL2utcpJsDUXs5ybsOMBal9vbAq+jrqtDHNC/qo0yJq0Bjt0YHEOppKrnVGGv5k2mB3uu43/
g8n0Mt4Q698zc0VEMHIHpZK1bXmDr8JVEjxI5CK/9T0DXkcNVKLoqgO+uixC7qev9aPsUFx83j3N
KunbojH3oDkg9Ps2+jCCQfLjNxZ419np0GNFogbvQZPxqeApz/r5cZHytqW+G7Oa5NpIL+6pBRjt
x1IkootiJaV0FAexAJ0g+k0y24ntSASB9ZjfnBWGPmtqJPHSOK6GS6ArCULRAR1I3l24JE/CUAiv
i+PEEPcxEFa4M7TJ2PRgIKX2fv22hVRzmUCdFEXOtCkkQSpGCTbMJFg65wfFbSg27OfgguhEUwEy
iRt2xR0Hwoz0U6WoBS/lgMQWWl0FUZSg9D3TckvKp8WvnYuQbRAOjE3EBBQuRT+2XBF+Ltct9bt4
UcbhN7I+f3Ul2vGHVTLtSZltj7Zs6JYIkDy/C5BIqfjFlMYfX44owOBS2GVVQSV7cBS1cxsrRdeO
WtDkGAJxPBJVKQ5ECiAx6UKhs0HqnefzgKrac54vfJgWjBN8fNlzQJd3bYRkNCeiL6q/rKHyQeuY
YbBqPy1r8rjRabacf8J1L2odaqkL905W2SDIwenaGQmivKoCok4sZB0ILtK5YWHp9rFKh+o8wBN9
HI+TtiO8CLtAYjFSMafGhwx/XvpMesWxZwHWa9azmxY5qhUcexuKj2i01uwCDnWVOlg/SvFJCfvU
wvuhocqRD10prunJzOmYHzsUNZoQbu1Hn/+/JpxU264qrfcMSma+tqgT9At1bQeY1unjmO1XzjCY
3Ex8H/YxbcVhvw8rvdXvFVldsZFcvUNvjy0bGv6OT9VjMJnZKTEDERdQz02te7ku2osK+F+SJiW7
TwQgCqKU2WiL6lA58+kmQwFXu8iK4lS+q4nhda1fofV/XbR8MSX02ktJIZTxrQl2AnlJ7kT2O5Eq
Pi+KbO/EPBe1wjuesxPYQqGWxCnYciIOvD0cZUQ3ckyTm0MTXnOkMdn7Jjl7k2dk5LaVivZWod97
5okXe2pzQoW1owGpH/yyA/dgAJfnSUfR2P7H/KVp2xEBimMvBLdzEX8O/eG2vAdx4L0IDpOXByP5
Y8EW5okR3eQFlXyIhJ9tsfiXxqUqujo0VllAPTg1sJq4nJcVp9ddloDxLuKQqNHvctU1XUeFtQHk
liHt9LV8sMJBT5KnWjbgpANOLNmlIu1n221Ct0G+gGkUjIHATppyaZvw39UMMb4GXgKL6TMQHRfB
Ih5q2Ygug+U+vWX/kv9RLuJzilWFtTDHqG69M4+2ajzAj3VxJSppTWnh7NiJmaSl/ZFXgJZ0pjXk
PmPfZ2HXf7d/+4wlkjoo+ADH94HOO+T/zluh3jUp/240A6wYwBNfq1j0DCa2HT4kWtQD+TrAQkSH
HlPGZUglWRWuFl9u5PozFbPW59Ojw6VyBcJBuGKk5wZap9MEbQbQfJn0hPspqJ6GC+MzGvXSJHJd
COAfq96xqR8tj2+hJZdLjFywdKr5lRBtu+QA8IzpQPZXgIAsv9mb0Jc7SsqxUpuc6LPwiXWo6el8
8bEQZm3dEZVRdMPJLV4AmZXHVF8G8iOqdBZ8qr6Oz4Whlfniroo4zPH2oGf+iqeQQS/UdprvLYx7
HXS1KFqdvsph8z3qEd8JBGLbGlR88oiAJx7WNfAmZcjuhPlsBqKTUeaCOqa3JpHVJL8vlu932lUa
4yA5k0xBtJd9cQmtCzcSfaTUKtAD6phIEuH8Nld/vh9Lg8OQyWySR67B2ExxTIMKQW7wguJRry4e
We7VPevIyqQ1rPTvycmLrktWU4aWzz0m620tWl0WpaKmtTFnVxNLAoK008rd/Vco9Pubk6ArU5Fc
fk1GGUeypkUJxXnrH2okiv5D0xzBYGX6orZaB4LUjfFAnxSZ3jzqR9hFw63LYwEClRLA5SeCRIVp
xsbjzMK8lcWKBEj0CiuMkcAoJQ3T3pycksGFxm5N0T+sFba2B8sP7UvGVtr38dWFduRslLEQJQ7u
mDN2r+nFp7EIJkEol8ko68xmz+hoFJeXgYElbuwZ/ikBm85a5jP8JhUNb3J6Zm4PmyQZQXamT5Xw
e4V+Mbvs+cbhGkj+IjYpJqV0EA2SYAmxlWusyvlHIni+zm8RHYGfHWiLfaVd346GT4FtfVzuJLBi
wvT0WhfxFADI76Oj8j2rW7Aglj7QlBdFALLtDEs24IsYBVEZGlsAnafZ4ZS3MvRFWmrDEtxiqOyG
2Cu459umx3/ftxSAUteqGtMjYMO3I6an87izuNTVYUSXQsIrqElA6bwqZiuv/qr3eiLp8Em1oP0x
bMjclK5mJqwc1mhcXh54J8Og4WdLXZ64wEIsiYXioz/FYuzIzoLl5H/UGu3dyvHweB0tpqPfbHod
o0d3MNtkC+TF7RmoVT0o1vI9O+kefRWoh97WiM9M03SDsZg4g9lg93XaMx9cBODyrdP5qDrqgNpa
p+q6zXc0h2eg7xXztb+/q7e3sufIHfh1xJ5AW7EVa5XV3sYL+V3wnw4a4jcZYIzlcnKH6pqZQFPJ
Klrmh7PLqe5aPsvao8UyMW/9g1GMtaqgS2plxlqfClHrcQn9GgvWtEEd6wW3PRV3g2zbTRHaD+mr
p14Ymd9LjuYaROPiqIj/Q6IgqepKMSUWh+6Zx4A7U+Zg3arc+vFBC3XNE+AsGpnc/kemLB++N4vZ
2YCtZtohZz+6jomb2umeBMES5fu248qQMgjY2E28UCbc6NBeStS0uKThl8Xy7lTbgjPTke3ggJm6
o4A220VGVAjhZreEOPn3KPrFj3GR1x8qRkBkAxFmb7+2Qy0gdqX7xDWBEi5ftyouK/YSufGOzbXk
mrEstFpXtPkj3WMGzGLGP3puRhyLeom/eXuXNz+UCOoBHcimI8PrlJmZq8dbUW1IbsARFI1OsGZK
ShKN4glcjlO7bVfAr5eTuixlqrSjnyrU/H74bMST9ScsvHgRVSdH3C3cyhMbTIrP+MAW/61zM7SN
GoYS0eZGeTkWxlN+P7J8WISxEGKBS2CocWVdY6Ygr5dulTn/S1qZBe8Ei6Nk+usTHMmenStuZGie
TBUiiL0LtvQTltE53Kdq5zs9d0n+wNAoqTduKXvoRK3JbkqGUH1J3AwWvsMKGB9/I2eijsKOTLUg
wuIgnYDfKCM7XF5GYN7/AiS7c5UAYBJITDgzUdFAiROGiRgoNCiRM01vNrlP+1WCOIx9L0uispTq
zRD6ppYocoa36nGxgD9tiFcJse1BVaSBYyT8CHXECkQsfhTiM/10Ns3dXJUvNDKoIWD7Q2ULZvh9
XYwybv3Nwq9VLbIG/2gK7tYHjfG7cWjBZxc4o3lZfLy5wQjxsvCP8rwZOcxTWqh9xIXv3MLdnoZc
MlN3k8flQDEPfqGvNKlmbEVlx0L9i6+xhZhdUW0xYc+y6eVB6sc94P0k+wJksy+wUr/6U1Z0VND5
oNbfco6QTjq92trnpM6lMhp4bbGsbl+RfKe4jNOrK3z788P21gwm1T2RjxYJV4mGPIa47eWaNywa
l1gTWH4XAJmUO+Ls7o8nVhPq4NWro95EyfZylGOL4x1DBZcKobdDmv+XnFACtoC6q5U+OpcTiRxe
+V0/aKNvOvyuG/dYIw8PmsZ72Z07P8ZWEuQM6VuhYP89jRLAoLcPRX7oo+ZqRtReHh/h1wneQJji
03qlsI+3WWdhn1a+SODiUZsDtGf+QA8Tc3M+9lInJjHDgDFaHOJQjoj+aGGFHxZ+9LKcgwjoN/so
is/o/tMy6BK6vpwfYsUP67Pb01/D7qPlnh55lC2I5d5o/YCRp74e0su9oAI7InD7JGSnSGFasqsA
rCGCbKTcdLYTiBSu/V88rTerEz9qkqDTiVgd2rto29Pr7twXdM3Wg/h976DbHWMH60epp8V/aqT6
zffMYnCJbusgFialhi5eGk76RzMqSZPCktTmvW/Zo9vneCXGiL/4kuEEjMa6sIQiU+OfJ0cmZ6x9
8m11s60i2nCTCoMS+vCjom/tCKUm/URZw/zy3E+0IUSlV46VZae+ZxJ/VhrvwjboQD6xrmqBxY7X
3oRyg95atMXVi6rZCnp3BYCmn/bfM8EcijgXTG3/LJZ4OhVsNQKVXRNwSkO73MLRh1yiNFu+xIhh
qnN4gQ0n210NYEC1Q2WLbEHl7+q8vGOQs5DJfBE9hSeMXY+C1OyM0nOqcCDMPlnxpD/smcrFjHsj
FZlFiMtPRnPfe46BSDTR/x94Go3lx/DFs9aPxPJYGQFPBB1r1gvZP+eAsXSkIPPz/3iB6vZ97jGl
GWOlQKXtRuRIW7ceiM2Ir75lNhpnoSemJCCLCjqwRfWI845O091bBoYKVEdBHILT8sZkSae9xEEV
T69Hja9PX5KCVMkn6g/K8ZuYnHi6QqgeBE3vTyt1hmiYQtXwyqOexoYAGwCA9MX1TAm1pZMEc7YT
pIJzOoDiGB/98XPAWve7Ul1ZXK3wzadYkdpY9FT03OxYyXdPD15+t/WwK+OLzkQHUqkuqCqsDnsz
7lXaWBFHFsa6ZqmuH9aJmUTJIabZlMQ3oMRajr4XCD4yTrErtdH/KOJG69OxSTbYG0KFnJQP2+uk
RABZBOtVGQcj9DJxm1vKub0X3/UU0i7plvFbNgpE6sYInzLBLE44FwrXoBdjji+09Pcyyvn/CpzW
JBrt4y38zDeqsIJ1upvSN5VSWzDIEznVqjSVv0Sism8j6UWJ0zoD23anas/sXQo4y4IbyGJGn5nK
yOZ495HyIKdfoR77W6vkOTSGQdTxbRYwH337mtTxBaWpoMUppaurY7b9RXB/5iVX/OHbdwIjL2tY
N62xkX5q+CdEGemUad0aFbGXq2LH1RSSf+mWRNI8NrqqvkySeRCFAXYNhdpyqU6lUvktWle7B5mD
0bdMTqT6TsbjBM1MLDu3D+eD59NRvvC2UpggLL05OG8E2x/FYl8awt7v0Q/TZKBHR33peG4rVJK2
F8eki2KAKPzUOW0mucBDyc253S2/RcC8mfQq9zPHRm9v6tWE6LeZjCIhOMu+GofllxguohDiqwNO
/P6KYwVorOWmhTFQQ0vRSADnuCNoY4ONsfVYk/MU3jNQO0TRaTkC8R2elVxMJoypLmF+VihuUNta
20uEpHIhx8zR8nmvqvgeH3ZpYxP7Wm+RtLmN+90CNCiiebg+XVUEE4yHPB57w0hd459f4XCgYP5O
SNelImV/ImBtmwFYLeziJ03MjuM8zQfy3SathKU+Rny6vVA0mtGet0+/LBwro0R7fjsBAiotv3OH
Xum3XPp4Flqq4tioPZXS6E64RW/USnqfrRkUF4d5Y/pKAKbGXU1LGqj+kK3EG1P6QuvPtWkBllka
8BXjbXeNKA2Yvyaih5CT9jn6vBPojrhSs5DGoh+w61KtUQW1BwYXIN/2FTUJMRUifm/hFpKK7lt+
6bbxhN04jKqsM2XroPEzG4CwTlz4loYU6ufGpQSgEu3mmwRKS4cQw2fGLgVwI+FYBx+1njIQnkcq
92Qj9hftWbMvekbzBThoB4DC3XQZzT2lh6q1LfpPJixrelw5gZd0YBMq6zpEMLGiOBBVGJDnxPQr
oWvLLxNIsI1aDon4x7UIKq05PglD6aX5vbwip+ple8345JRxcx67xIyOugvX8ImHR0KKpWGyDkBb
+DnMr5EHsSFsFrWLjtnCOXsAvD7C6CiPE2w3UxN2WsGXAzmhvbMxRhJdwDm+eXc1j8BLzvHDaLQ1
zHFa1vHPrVYhHYwklYbj7DD1Tvmto78878RSJpMOSDLMlXL02rruPMTF2kV73xkZgv7fg5GIrquX
8UKFeWhpKu7JulbblKIXQ/Mz9cpcLLGhbpPUBGKcUnMDxsskp7YXdAVlwUX/ZdTJunrmLDJfxYH+
z2w2wykpJL39bgtSeTqjpyQlHbt0HoD34Wq7kNXb7yQZtTRMzMVrs5to60JEU8gkdeoXCiu9Iyb0
4kc4CoZeCjn03en5E9JqqOHWaOtCb2O2gcvXjPfyMB62B5hnnubVskuJhLVExvaG0h9uiu9gRoCV
fq/+h2XlyVli+fwmnOwA+z2lVky803mIwbeOyrIhYS5nTpNr8GUQmUpgUp7lnVw4kPf7R46889O/
OSGLiNMr9AMELIek0bRHQjp/9d/+3glqlxDLO0r5qEbtcxSd7v0/TwgQef9WtS5YLTNVbGcBqYWS
F1OWeJ8/OyoFIe+3fKugSvMYLdF4+92l4fsAy49DPIuvetYyOH5/4DGN9MtHjq3DsXwszbUrwjXX
MfeqNRD7QTEzz+DXyzfKzeC+27iKsVYplmOXzeiXoJRP5whlTx3qj1I9vgDS4qvcCoP13X6MvzUJ
NI8Nf6667ZOqsIyYzmwwCIQ0vApQYi94rD7F85oNM523QByifOX6T6DwsvmcVhHRJeuHzQaAEtmy
Yo2lj3Znv4JJxhw/qOVMJerSgD5p9tMdqvnnAYeW3hQ+eS1oAETMl0Rh4toSXUL/ykgMGOkUBeMM
C0Iv2z7mys+X13CQvKHM8MiBsSZbIpZ6jQHTvK1Npvmb3THdf/qIuGQhZ1bIp6deViAa6hBKb97a
TfSPDk6nvfiOa3QkK7nBQcjUaAUFGRYJDBePbQBwbl4FRkbNLFcjDBcJ7AuAWbEXc3hnX06NoD4F
myXUofNciTLE3i3ay+B30vPGcmbEilYPpyQDriDnkSyFHAnIxrACV+43A2p1RAcAxgaGK/XwB0pA
Vq4920UH9fZGi504KlrdJmpQ93J4LvLs7e/asNGaWTM2HFrgys646kjs05Ea1SzuTmlNASW1gvjD
rsNTytilDHD5WLYCKvAIVcH2pg7Edv9RzzIXZMFp5xjL31hjYcf5St9oOAIzygZbLQLEbPr1lKL1
fzg0epFWS71IR8ASGlOqhiX1SYLilfZr+mKB3KACHGMGkRkVwaOG/OU/6Z3nfSpigptud99ABpI0
ZTfgHkxPHF7jA1CPSA6LtkVWwsl8gRkehi7FpW0C/VsUi5JBjTmmro4pDUs6GOJcOfLKBw9k4wbb
dNXXn4yS3SuXVtpELKgEO3W03fCCFn64+Gyxc4N1btp2iXs9nRE6dJMTpKXGeUJ8NZ+rQ6QHxlKi
bGPSh+7Qah2xGF2zQbXPzCP7L9nRnPCh8KsvW9r+nOhGUXqedjHWF0WyyVmsYyUWPqc3ScfrZF0k
KcedDRRh7SO+M8xXbq/nUrDpelLonYQ8Y+wEeDzl9LIlPHPCPLZBcF6IIIvU3ZkmQj4mA5Flc5M+
tX4NyO0cRIrVnnx9jJaWLnYI2Qyu28KW4gcOsY3caSNspJ1I5BlsBs0rHJ5IdyX9lFih1UiuSAwM
FkQZIGsum0rOCkbf/gaY7fsLaEdLuaUS56Ku40KlZhe1/7J8+EBv15CQ0mNTQ/ENDmOCkbWwSeek
TtgZmA1nQ3EuNYbVlFdCkwx2Dy9BpgRcRUJ5KTM5gA6/QxBRlhxf4lM4uQjRtWLVHDSb9NmzkDJg
KXH1YZDyMtgxiKYtDUkIuHKYUKEUdMWSpQ3wzsZNALvj4OiQwf9msqAOIbwbvgeEHKg+wOIG/Jfz
B399Gv1YXjvZlfrD0jXWc0oID6irdFvMOZ/G6KOfmoCcoXiHTpKARG9TIvgw5ZHfaBbLfpRBX2M2
PrxlKzYVQvndw2JWrmvmsxrT/aqrTA2ipDjrsuZvJsJwgIkHaSKC96lYQ6nI17Ihp5rJ2p3Lw04I
OgbAyLy4oC661tQqx0AylF4Gs7rfrc9SKj24l5YZaE483xTmPO0xvd3/2Yw6tZDGclyalblye6Ma
NzZxUzBTRE9aR/9+74EPhlVNEZ0atLFLS5YPJwyGAYDxp6HqiBlPFVrMvGQhYtY58sJ58wmyLQbr
+J+D/O4cktJ9/Gt5qLJnYghuG6Jk+1JUxukSPqS+IEXt/SM9y9Mq5bciIEn/TL0B70JLhqwq1a79
RQtYE7A74SlrLlwL42ApFkguYS4t+kwlfV9fNOz5UUcu7z4D15UOkloH8Mv7t1nq0+ZPTCDMi9D5
UbYSLMlnbY3mU9F9HIh1th+/JLqyvFQIpq911PVleXwOLZyoUiqMekUnLP8mL6eiE8Ae0oD5Hjzw
30DiCotYXOnkPnZuEk+eTuo1vbchYamI9nu5jM1WeaLhh4AAxxGeuHYaJMSmF2qs1LgH+b5s0PXN
+kvvf80EXsU+3gYizZKseuy0Id/BU3PC13hjdWrB5Hc0wDxWeBrdDm2p0Vcv00y2wdE2DLkFIzhj
MmqURWZZd+nLjibcBmMab/eC4brUbRRPDtsMaBUG9ODzrzEk/u8QwNv9pzM7+iu/nKK2iwSpqRQh
y7elf0y7SaCWTEuUP6OdPCJ7HBveeSHU4YZiKVQW6N5klPjNzUY5gUrAGxOVILX6haq5Jo3MCgVf
OqHkklPiMljfH8RDoyMlPPBk/eKwgC2Xsd0j7GUsj86Ip+EIXJCO0XIpDslwIYLPYgO29arxZVU4
Z3S6e/1qrS/sMGHAugmkvyqFHWsMWTpN0MToniY86G7KT5kiBst18Ydx7dEMsNxE4SREpWE+3FCE
gx109TWpL845yw591zwG5nrLHGbHoF2et0Z5E6U9F+chOjLYTJjiNez1hyN1j329qLjtuT1QEb4L
kA8vFm7xhVOXOdahIHHVwPuOkUwfkZxTDAinLZeyzBfmB3MkA/9ydNrlmTeixY9NTuVInGJSbfLZ
6aNyY5mBK7qB2H9ew0TCtQqGgM7mY5V5EveuIcKZUsDqn7z+jrNy3JXs1t8QQvdIeL5axk8InrZM
DkQgT3mIxe05VoKtlyhReApQmcTP1uF1EestdpGoiNJFtAmuVOidMgUYUNQQ4RUzf6hKfPJiwp47
rrqhzQwLP/Vx4r33+L5YbYlfGh5Wwh+s0ZgghOwW7L8SEG2m75u158HqQyT/PrU3450xy+t4TBlH
2ufuZY+j5oR3pbvYReLBLtQ9Y4vTXfAQvYZ8R5PqAgMOcOuEMf6+f/hymEYC+MFQP9cg//xVktYR
ZiGRvwX4xD1hfw4nJ2vv4b5exARxFEGxnQdn8Sno58yOV7HJqrG8Lo547/x4Q0oM6rIj1KJSHzqm
G7K50dDnNmTmszgVZpMzEVzcpaNA0rduqVgGxvI5uWPzIec9TYKGMNVKXKBp1QG/3QNWxncka/7U
n9Qbu3FRBz8EC5ARTVv2H/tcqI8/mUZFJOqAZjm4cZ8rj4E46RdrQAVDV1U3nYmyNIKDih2jToYx
6Sjc2Xqy5ptGkQtYqTbSOiXcAF3CRHoZ08X08U5pBgJ1nYcx+u7j3k8ESoG1lReytjNVCsvgJ+4+
C1W74hWwUx6/vjIGtjVH/Sci4ixiyY3a+FQNNwRCyWTFKkrU+0K3DrwTiW+KSo6VAAlzyFT7cutM
JtyUWiYJcnwZyfx7Io4h7Yl70BNOVLL8hnJb5zIMHbUD6RC4yaSEtTqqcDmXTE9FXtVB9R+gBj8N
hv+JMhxa+8BTLtvvxvPTwPwaa54uvmv1TJTe6a/Y/6pZXRpr3U3bQfRR8aQW8ry6ZmDb/7Yrw9IB
CfgF490SF4mq3pGlF2vKxH1eGSqbOpoCgUXt2KPo7yvkWcrui4nc39aOqyW2OSB2Fko6Tw1zgNfa
YAuQT0vvClw4Alk6Acdvsik3THV7GzSwVVVVRjK78oGaF8SEbc1zrXjJ1zOFMPYKmyxFDJ2JfWfz
uvnmKAvaZn60Ht40grXd0uojdDsxqtlTVO88SYrVRGU3Kd+OU9XwSR7acDvdqk4ULnxUOVXKjnP9
Pjr9mJIXwne3uvMfZtQcjHJMRgnhXUxXVkfneS5XEtltojwltjOjnW2VGqHeWeez6A756lyVvJo/
o7VEN+iTAGMKgqhAZ6d3j1UpxfwSq/dPeGJVXODUQmOE74C2Jfym0LCP4aIFhZhQa+bz5cuU6EPb
y1VSeLUtEzyskgRBQKBZ7AmWo/OAObH4ulNcKgxGoLpnUemPx//aNRyQwea1SeQwKTjtbaedcQUr
savNGggmapjUEL+nm0NdCjPqCvt7VxNy2xhv5c6C+j7mui5DoXlqgRJgR5PEtz7JNsaW9mralR01
kJEhyCB831e0uGwO2B3MOuYSwvhvJ0PWCuK3/QaeaksedYz8xqr/teZBlJJ0Eq4VGM/+6m9/qm4/
PzRRWY0t1MOc8esC2yTIcc5HFoY6LxB0yLGx2935jRQVIrrGIy+ipAGUDojSY5wniX5aR1whPRLc
/7a4Wqne+xdCBABXD9/HCfwdbOKccMFuVekyLwiNvrlpVsMiE8zGEU89YL+kgm756J+RfilI7rkL
SG7fKU12CsZ/6QP/7RipAvzvoX3WxS6KhM/9xMr2rf1EJgqCT1Lrwj8Ao0wvZxkgdNK+YmbmIIHO
0vKJ4zajwc8hpqWkO+CHorCneuBuxoY0fxUKR99hFDQnGJW22BZU/uZiueZNxEFoxiAOa8qb6zKz
c6VuuzhCyGaJ1i4Pw+QZcYIS5iRB8u0YKwsABNPCXaCid1n9wxwLfiCST1KVQBAIU7HhjTQqDepk
42DGoyEPO5VO0wfcJfcKKkrY0chl7D5UUeaWHsSlpHvy0bjop11GKof5c2QiYMOHOYf2MN6glG9i
YsMWqzgHAc0skZYOTtjLBoVHQG8TaNf+SBtGDJjk+oitX+eDXb/IdXi6ksjOLJWaqh+4LKguz96j
GkBEoBZrBinZonWJelczKcA+zwpT6Fgw2O+qEUsc61V9Qeh/1lSM7t2uj1DGAX6lcePQXERPEROf
aVDqVHY22tk5QgcATeQV3BH7w2Gvlv+LsxQcVbz7r8rSH4jwVhlr3D82cEhd8dFBZc9tw7U8/XBt
reQi/8ssxM/vYudFh2V/qYm0h1T2HCU8u/vVf7M62Z/yfnQGwkjv5IibZQTGBdAlztjlp0zvWzcv
zwfg8l0wcMbqSv8XwNA5IWC3cLVdtdRYVUMLMJv6B+u+XogGON3xqxaBLNbFvoKIG+yth8zlntj8
pVoJmKBhRe58Zu0nAl1tlvGnyI1PY5DPnjr5p5237lBgELahGcBguo/p1gApd6fO3v9lurzEUDOM
whgrqdx3qN14E80ZQiihcHMeehCK9pqDuPsFYFIvyVU5GH1VpDik94bbKdHBunHYDiZFjfkor7uX
b3e1kKJ25JiQoJi6UavXULsOo4okYq2M6AtzPsy8nDBcKXEFICaLI9Z6qr/Pu8wFLFgyKMCaThWQ
fJNdvozATRP0LYw9Wx0gnbiClVJpXrLLvt94fZF6+QN02uus0r0lNrahf4Lni9Tfyd7yrVIQMxo2
ZJoQE2hIjne3S7tKUWSc7JTHl2OAU3jSc8boZtrP7uTTlW5ar5WPlqG90nF0ErnNVX46JXBxnq7J
BT+he1M7a90Ta8Y5RDTK77/mNHUEDc+g7uDUZ0VmzHSKn2BkxB+vqPHkByxejIIVqGnPJf9irvBo
PQncylVpbX11W0+Q9rwYR4vi5/DoAnKZD71sdV+NNn8/UFEHJvsrLVCA+ESdpvE1Z0MhMpgXT1pL
JWAWvCjwoHfXqrwILYGmaxnkGYrRx4fAw6SuHP3m6QWJV0uMneZIAQypRnFUq0erBFps8e8D+geg
nGJKe/Cdyj2BUDCNnS42pzG2apjqu/H/HuLg4ORwbqSD5ZK6PCGOZVNB60Xy/OfiYvNUXSAzgPj1
R+KHez0JsYpRwE+Z7iLeBT9cvJmdjYgpEWTl9RyMPdpTFpYspTtfui3QSLguGzfeYNIDSx1vQ+dN
VXaGson+y5dMG5ousx7O7dyqejkb+JGn2cYg7Upj2cq7KHe8BwirayAqHzHIEa6DnvndkDvM+mHp
a56JmdDRBaQKK6GD/bEYTBpyihuyk/2jHbw8BZ7j+bVqCY8Y7z5U0fXBBzgnOSjldljC8uoVpwPM
WbF/MLcHx/IxqYnIv40rrdbPcIVtA78ikUzl4stq9fsn1y6J4EUyUh4aIjsKcH/zUzEVRed0pZi0
sd9MWpysfov2RV8n0zYvM3pLL1UhHT9tlmT5qQtv3YpeiuY2KAYrc+W8IYY76v+D76/SV/4PX5RO
1Pibd1bgfwKLKyDiSuM3wQV0e5pHFf+MzMmLXpaZxd15bBlYnR+GKcdAAZf1culGrNI81YNMYmGx
7F5v6FpU6SFaRuXbQFWn/Y+in1GWYkg1jP4VCDPIJTruBEj2YSYd4F6CIUrdS+Twi4v7EPwbgQ1d
8ZKMpdaKJ1qqSo6NcdHQwiBh1Ahfp3qZAemkpR1LQkbxfR01DjEcQ/chq9uDs7YMyh35GlXseQMi
wluHyD+1632f2rt9XNvHJ+H6BpBRgrJFMcalCS/UUt+7hn1Ri+2hb9U41/tPpFxhBFNgGvr6C7Z0
uQXPawWLyDX7K4CMuO47zj5Q+eTKzyjNVgSsP3yB8IjJCKWQSlpcK64VJGjT4ToL9hMB2y6TFAqa
z9zvigj911MsmyyITz0EFEVjXh0oKmzz3poeUmc0ByX1J6OF14Wq7RaBXGWVTXp8RtZuJ3TQD1Od
uLzWvEvTARWuYAH1D8z07sivRLec1RW9TJMH+3MsgRslayNrh+WTtDa9+VY4ocw0/g82yArH1lvD
HoBHUzBu3gFFQnjzrZoiukHVlPiwlijnUcyVoZgZ4x85P8PoNSeXHwSIwYQkExruGEZbG0K/pbZs
trPowLmUgzKmwKEAezkdy+R+GX5hPmMDlv8d49DwsHctCPICKOi1fp9/s4XeKtioauqjLjQXjHgm
oRmGYD0ghtgdmuSJkTZijnECzJaKa9SiZ3o+18kdDwwrRKyB86Hp9hokKWwpA2JxrridVGVuDAJS
8wJsT8BN6jzj2zigBghjXsHCX4Ec4R7/4jkFRf4lFjuH3i5TmYSkIRBSMakDWavTOcjC9JG4e9NS
PiWjtNy3Qy4jUxGmJXGQBeSkRB2UT8lw51qVztp/er9bzMLpm4vTMIuHq1vmUE+/G9uQWJ39cCgi
Ut42Ouei6OsTdJHOxhw6/wAs7sYPXaGaAoiQNqcIxAByyWirlVwrs53v4V7SCvGULvyeYNigvc+U
FUWdpuHaH3feFEWzxNLV0dZ57hg5IZERkytKEu3YWLoj25qsdesuFLOKowCFc4xe2Ydo9FKO5h64
0fjhk5owb7X1q5p21V4hSAuDZotwozlPF0q4tZ18nMEms3aIjmEHPdRs0Xy2Z4u5zw+jy7aaVDMm
lpLCy25ofegy4S7AzfTrugFWbWvW9kUo1GaqxUfpMJwAnuUTr3/79jePfgOYuvYfYfwy7VkXXJUX
8MRcu3uji4tsAVeUhYT33TuLYR5nZ0cEhUsVs2ihKJIh39+B3NJdW61ri4inK0ZLzYIOUrsTVI/B
RkH9lDbVBN2luJsajGivFSxzToeCE+06w33hRCnr/EmZdK7n5Okh67iZY+rT10Q24IlyDpma0iQW
3BBEdDxhVKQ4PUSjf1h1xYG+Pnk6ueFuJXDpb2+SpqpOXrBXGzDLg9l4ID1Uk9OmyAehS5CFPUO8
gaezBPjxBqkxMjuvtaJVdaBLfusqMDMUFN6yqws6zI75IvgElS/A9/+bhTR4B74PoIJW6rXmRYDy
r7Zt90tMamWm/b9Rrz6NOu2MAld2sYxJ2mMtLYI1QvbzfUcTcmnT3MX9Xi3Q0qemwFbL93sqeYOE
+inTVVfvEnee8bgo3InG7KMp52Wrj1mDpRRcgFq228RZFLiiwDDPWfsSYB5PnMulmaigmUtYBa5S
0ZZKPeeEiBRNRJ5hlXNWgGlkm8x7KAHjnbn3ZeOgWpdiXF9Hked9tUFxRpbNY9s8mLI72ryvdgFu
lXK4crPtDuuptXvgxe1TgXwdy1YM4UCnIRhcerYLkQQPUHcZqXbc40c/wC+yvvAQyu8o8QNc4V9q
h4vp+H7HjAjKs2UmikwrQJtIjbB3RWhkvMpmKkd3Tzer2x0fTRM5m5KWfLE9QDmeVymyhcu70A4x
Oq/IaaOzkeyqc+206Vh2WLSM0N3zb9tcKq9BcdIbe/1pjkL1Nga8D6iFnZVpHhF2Ef3hiwUKpJmC
FrrQE0m8hCq3LoFjbIjpncoAE8Nzew8gv1vfPp51QVr6gP9kKKQMwB8U31qSV9sfh10E6JXXfM/Y
jLTIaTtKDo0dRXOd2wb44uy5hZkVHhNVNyiG92co3drWY6ptiKr2qIuFmFlc49m3S6Xzolfj0Y8f
7s3stl6hkfrm2TvlIRsULdGu2wztxmmuAFVSBJ6oe3Nm51ZOMRpIUmfWQ0xJk5oW8gcUFnMBbY4V
qk5fBVJALzCoHyTIJHreRVVfRKE+mC8UVat47RLHReRZbIBR6K/3ETGMEdHoBadRclW2UXBUc5EI
1A8rbSXA0Zw0m2avmXkcd1mf8NOwOZdGW+okl1z0DwRp7cTlkg54yldDdbr+V98s+dlhkhnYBhwq
ip0SLuTPfpwFog3XvJ77JUjsJhbGcJewmvgAnprn2ZGzUdH9JnI3SPY6mfzT1SbKjLRjcuyyhFLQ
GwWJoe1K3hRdqGhFpKsqLDFReTHF0nVGFHdN2xDhZL/QGftdOvMEACdxZrAx7VTUni93Xwk8uQMS
+xZzc1YYGO/ffOeg5QE1KFxkRtaGCUdRWD80Z8M4pVaCv3kiUhMJH6fLCw5okvyIC8cOtmeuUwOd
RhxTWSQ7pLmPi8LzlUmFwOMyw2AF3t+T0UqEN7LfcJ/CsoGoYCbUfME+IafxzYcKzc/LFYpgXy4z
HKnMPjp0b/FGWMvyEAHcYn4BINOmICv5AqCth3IHH3axHX2nuqrht8d8OJKxSGzNeJh5B0kdLWcA
TAY9OtorYCQaXVBniC3fTXvtJDlKMN+Mhr4a4L3exqBT+263mc2s/KIZEGAjjQ7aa/G8x1pAdeET
yNkDfuDpNu6nc9NPfJ4JGTVQCxoR8MdUNB5xfhfS5dmhYoduMxQQZwYZa9QfTLLS9H5Lr5+zUxMj
7kKX2V0cmscVh7JPwpSTTxJj5lXNcTF6KP5JwB8FnNpzKyJMThJHtybutWZ1D0LilLMdZL242tJo
Nbjp67J2mYrbtZ+7dPpxudOLQ0vQey/qkbaL0JMtKKkS2Bt5HQ2BTZ1SI6WIbTdZudbLIKwDUcMl
sqdzO8u/t2OjC9TxMC2hh7Oss/ig8F55e474Xm2yCX50ZjrO5VKZmYzKpMQQsN8TABTBCRQFAy99
Pqe0Ea06EBZtit3jurHYusdZoGc8peqjKq+LDaIaU6uNwrY8mGBNqJMj0mTd8ER+7L7ulOX8zJWp
wDaQIAGbpYlCOK6pSw5CsDcyUlOxM3WoL1afLGLZYPQQaQS2ZFIOdEMCNWPDlFWxkJJeqLzJw32b
cf9IDRNtsPMUV9zWt8l9zy4JqVfJtUU9UfuxA/F4qnC5lDPBRv3qiVvpAcGNQjtAT9l9ilLiIPzv
1mm84iGuBbk3rgTFjeb1nt8mQ8kr+3TttaETwNZAMauR15zzd4M4eBi6vVifDw7gwQT/ktJGEeGB
TbSYuPt/QMP7+95D3lA0SC8L+F/by9fWIiE4OaLoS3wGotWceUr3azj27mYFDQnd0mbd31xPeuOX
+s+rckukS/82oUoO1w+3mcNBC+OpxkpR14RphrjxS9J+IBTuqvrobMeS1HlLSClGpRyiHCdeUXcT
K2FxzEg6TYK+z+rjzkwwhMshx9BewISwpKaFAUnwd4dk9GtLctZV5F4Gr+XwlvOS6p8DrWOBtex5
ijzEaxzRyke2ffmKwYh2uQukBdNyt93QODzx2iGLSngoLrUdzaYe4n1OCCtynvsc8JUbzlG3sEQ7
O5o40gAG6mYEF71h/IuvDox4SS7A/MSD/L1CbqSKWxssRPNVS48UQgBqXdqsFNWNXsHYq49lY+FF
YmEGQpFj9TuC0zgXn5ROv0ERSGyboP+3N3rYwqV1NumoYWOCU1z8Ty71yAKgIqbqffoQqp99r6t/
mvUdVfFCc+CC1fiIoNicDknukUZwc7yrXbSB89yi/eZPBXiju+tRIK57I+S1URaGT2ZK9UPioKmb
AB0y5U3izupbHb/efR+FNbgx1lqi9drMPKu1dL/iXuiCaXHXguP24KUfWZUB40b5JMMQYJS4R8lO
6ScHElH/UnwgafjG19j8WNDuy3fqLp4h4Gqp/dzV84uytz7j77AztAXoMkW5+e/cw+vvdncp9riR
ykBBtIaLV6lXZ/q0nJnVtBMbN73AJpIIp60CZhmEeEQ84f0rRdPYo7Grsh2VVlfdpP6f9EUybtSf
bEZPJqK0WrSMTA3gwLhnZOfpYLusDGCyf14Pc37mB5//ZpE47FM7rKgqlC3XxwRSJPlq/nRg3dGY
kgZTYWETi5uwXW8C4PVwcT5HZywPTmlYYOdLtEDzKfgFazXU10i4ovnmzc+esaEFMkoam1pGqu0b
3x/VySuH4iqov+tsw0HqqfDTbaLLOwaIv7/aRZE/lkeQhsikeTRB7T/1UtaDRKmoI+HLD6tdGMIl
GdV7oDx7uLkCYdabCEzx4y9V6jGEAYXss/PM/OpWj5GeXAsI9TaIYOPkWHXj0tHx2GH3VvNaPNc2
up/vrva9PA7VbQ4anayEqWDtxn9UE3lIjH89Liahlp1BuSKTLNhLbIhvUEKBrsiMvGOf4+b1IWfi
URD68LdqkN/3nnOgGaOz8mzNUsmDzEkPcf9AunH3kiijJQ5e42zBI0vTx2BTd5TJlB2pG7zfC/Xj
xwthRmazUcJLXIaSa3q4hLRkXVQ/QuXFj23INVaN1C5ABHx52xhwG6QpmNvlJnntKjz3WKPTC2ae
6G4N7O97xIsBPIPO5FtyO4g369XzZDWvA04/QUAYUqe4wpytZ+I4uBVvgm9JhS6c0n3BR71f9kzX
9jLlHgkRkg8sXK/u0HqEfLIHu+dNxn3qUkf4lP6RcIofuJFVGtPDJJeEyYjXJ8OsBSuK6ifDyV+i
2hKVdOFNEdnIdXtf9xu7UOtBbmJ+L6NyEgFp3TGiO/u5ZNggbA9PPd6itYo7/pOOcAJ0ErjkB0EV
zjyrTBYmVO9xyf6nzNbxfzv/S386aLZhgHUYdsiyCrC/PPQ15+bhs7cBCsQYr1s6yjLj8F/UIuxp
2Mr6TiA2QaycQZKGbPp4wAr16v7UTEwPpnXm7r9PE+vNQ4x6EC4AooZOd7avAMYIR7bhvhGmcf90
xU7zfdfAYOkaquuvUocanuwKmTQJKRH8uH0itgLNNp60St1+rxOe0enQSdzyJIp+R599AQsPTP2i
y3Pss6RJuIKQAsCSz/S9Fj+yTWlLWg6CvuNmbX4rDvwvbxr8J/v5AkVK/uB8l+rALbNoCKngXuoU
e2LV13b3Gf9SiEOCA/G14hgm4EVE6g9V5N576b5Ld+3BDwKKdhglObAGbRMKsMwD7PcDH8oTBRC0
ujlLAPyFuGc8U280piGzt9YvPoYKvk4YqzVHpYpDgn9Lmc3qR3j38G59Z+2SCP9r0BN8Rjrbsr64
5OhE+U9DLxDWgwjfoz6mKwZxuAmJX5lDKODGxe3cSGzJ8Lx7N/vVaxdWmxRAO/895ej/Mkg1zL2d
Esrm1lmaEJ3inFaYcpbbVAEiVVjSPv8wlBf7HdEUdgfzkDaKTUt9IbS3BEPIYagDx1BaG9CEoR8g
cLnIeb443hMMXgt1m+Osw2JhZtgR58q+6jVuIj2pjW2evP7pATW2i91Teo3yF0n1ul5WqWQD5UHC
uXJSHTR10+U57deW1eUKs3XLsFgKMn79w6xxpKVg0xvF3Ge3rXodR6xgzFyYsBF3Fn8Lv7PbOJYq
FsWxYe7vNL9eThcn5MqE5q2H/BRz3MWwo9mJlozujS233FTCfPA6lyqrrf2vzilPEQCDQgRRewZd
PiM2lWq3DyWQKeOB1GTTMmK8XP+DH37V1J3lxGit5TG1vhJt7ihtgrl9bnarzrVch9G5Vmbwm9fi
5u988WsrQBiWSdo7/2SsoncGlATkcmB8RPEKH70JxrY/wZMit9NdaxTL3CThvLhtneqG6qxeqXT2
ExSocZM6NELSFG/oRwClTSZ7J59luH0ioG6ARIJZ61ZhXqOCs5WCfVNkKi+Gg8jgX5pQuR79t971
jAU8ShOLHEdsJSI+Bmmq/cDx5ROw3TncGk0AZxBUmuNzFgEDJN3Iz8Etaf8g2gX8YlCwSzko6pzL
S1VG2wruUAuoa1Cm68ke4eBCBirubXQJ5wD7dwUvRu8SYmGGW5zOCUlp9huga5lOLLPRn2VZnRvF
/foABCBUKU6FD2tCsAQAsnyI0KnXCIjoYAlP3+hLLXZmWZll+IoB3RlGUssizWKO4c22YXdM3FFr
VdL96Czez7UYRycX7+F/+z8vz2+skkMDV3vC/3ImZdpADmoEGN4tF1uRnaio4OpuaN9UnybHzKh1
Ph387aJ353rTcWbwuyB0LGE35R6th9OTEE9rdSfHfijWKGbLNHfRd9q15DvHkzOCvN3tw/K17Cdo
pSeydgNWwQcV+XT/xwav5IN0mTu/SssRfaq+utr+xs7E2OTkTJErAs3C5AJT7a7j8qQULcyEnM7x
GBhZqVfMmAlmJKYIbtYCinwsU3JiT0xjXXhpFMIBK4rZ5RxcxQd3tZGNT2zXdY+eAqP5DI9h6ANv
YDSglGMWXLrkZijoztImEA2D45yUusvxGtDP8fjuHZ8nJA9FknMl3j678u0fDbOqDWCEeIiWLOHv
Aybx143Fv3v5DpnemV3H5OTGn0p/iq4/BGmIt73yk/nfOonuLuf7/WzNR4qn8dYmoOCTehzes2HL
gDkt9rit1ZfhXTgbuY203JSNmns24OZXDH0dgNv5wibO1AKlFK1Y/frVjp7I+Kml3essnx/c6P65
7+RUo6QKHBRAYi3U4sNsC32+1/4x3OowhqQGJ/dfeyenCPA4b2+JKW/bnKYNTDwQoRyg16fFzMId
e1jeb0WMzoFhLMBl6GLeUia8rpr3rrr7tW/xGToJKbHE518z0sZINFt0oWEGyQ6GZ9t2xNY05nVz
jeZXSoJLj096CAX0mr5xxgh0S6fjMarTbBkr8lJOCq3AqXHzZrt8b8aAWiEYuP6PzyPieZ8hClOm
+BA/fc2AnKfkXOoOJJn1TUqZQlVQbOjjhBgejJYW3qNZQ+zdGLnOONVbs1FZkU0f5j6dop2/KXPF
0H4yVFTw8kt3fc+2sQqgUX5+dESfACC2ltTYmWigqZ7y8kE449AcHHtJ24l23WYaATFRFa8Nv39v
9Ud8ZTGDPI2cPonup5Ca+xfDHfB9KSxD4l9dTYhjksmiJm3fNJVX2akNefyf0XJzOay71PPRGHVn
J1z2MAGKNxpmUDC8JArWKzcgV2h3lNzdjwAIzW+C0ERxrCzhWmwc/ptk18HAgGmFl7lIAXuQfA5E
ajsi3nQO/ntzMlEQZh+PRfHIP578oeUT9foqOekIAVZLTZ+T//S1gUZ6uECWcT1UJaJPKLEMsibD
YRb8ymIxkCO/ztMxoqOhaFa8hx2PCtDvAz7Dxi455QIjW/uQSeld9G4+sZHc1lP3ICBLS1hHnWmj
u/uaVkjGfKCCemsPsLmlqamp57fA6hQmNfArf3DAJbAO8UjPEH/8eE83GfZlo+xFyncN6Ctyg8vD
Jq7pfbvgD22dbJDx8MPBe2Iw8i2woAGg8HRJxAR9/ixcvn0xYgZ9iNwLJKGe1tdtYqI7braPf948
ecDoMSJkNd0YlwHV8i7kVQducM7PvEi0aCGV61nADUd5BBoPwEN/5uYs3MNrrYeQX+oLpW6odWQi
gviLc5ohMf/0L4TyKGJpk+IpmrfxqiawUHT/AHD3kwWW1glEiNoPunASLVxKorm98BQBMCWi9oem
S/AFSfrrIk2nptWj0rka07usXHrL/INGr3BVmjYjD8O9owhzOAtMW/Z6fXqD8zlJaeWGp+ymlLkM
GP3esMVdx2qJ/S/mQ3boCVADNt28+MbFdNg9x4nTJsiaCAYVqsGjPOaxxskw20sVg+zEee5gWImG
LlZFnakhab1yAV6wm1HDbsCrDf+TGNV0HHxS6FVQbZM+mq36gn1UA/R2zezjQyGydpmzls2TnpO+
L+RsaPtnVYJ3+3/KdrXKoFibGCq6fr9Hj8+jJPn6UDb6pWUuWYjfwM0Mjvi8uPf79u/QUnDnb2Wg
w104a/dNbDzAsSfVX3rbwIuZ4RK+KYbgLcP1XOxAujibloI01HB1E5WsTciY7jbNCzYM4EAFleKm
g/bevzFzRHvq0CgQou1oPmZ0D7Cuobc0yweQHezMYH7aJl4/I2Z/Fn8PrIDdw3tLgvasiui/WmZs
3d6LsLqe/1itS5UfmxzIAqvQxjO4UyTlmPybNK7vs8oP4b77rAEdH4TxxkKvDiGaARDT91+MGQQ0
debazVWvVAZ5l+Re3LsXdT+zjnDynxFWPgLaee1EXYRMLZ7EYEM6yoMgejnFzfIl3hi2dlDs56Cj
PjV8cBvq3DwRsB2VOVE4jOR/0IU9Tw+fYjiB1QSagcuB3HHancW0l/p71Tw5p4Z9ZBh+yyXm37Gk
JDumbAyl1bPlqwWrpSgIC+Y722mKBfAMX+YLcaOEc7/F1F74SLtbLEFAj2nAXq0EDsktRaLXRC0q
perFTA8yY3MxsBkutAotIYCQEPqbxWRABn88br6RjjT5bhQuLI2+yZYJG01gB1nTfB6hxdd7oK0n
MSVNg1Hh4yL81Gr/4zf0rkanbHf6uUS7BvZOlGG+SrLiUZzgLUXDjqTrOSERKnw+9r5Wa/SZYRWD
Br14h27hhe8eiYpUOkdllAt4e0PgN3yR2tilMxWQjE4vmoy89k8663DaaRCMYRM7dQaAHt0l8j4b
5gVVgi1EFC01KqaDJZqmZWYojmE2RHpSXsEg/Le0uQpkIs9QOlQtSAKBfHuB3um2Fa0lHVmEsNr2
+RcfPV+XKq/WinooFZmDOK6Rf3QoY8Ay9tZHAyDsBopKiXVN2/sfe0iY9m52FK4E5X6D0gSF+X4v
zUgQxliGLwMR4/9grG3vfFiP1DJyrnncMeTOjPyIoLGiZMoQum8l21vyRZdNhmdVbOVh3Oif3Yvk
0Yv/drkWnudKwNKWNLVg6EMatpFpRqZFxtNXzj4iAglhkmZ9Z9FmChCpSKtzEgpQwOgjTgw7RqBH
0s3iilDVKmy2Wa0yXjR4IyCjHU3pW10kqbQ16/X8IFvAXh7mpaNopQvZUqu4UbESpLDwQWPuDIQ/
ItzYC/Gtt0dPFvc1m9tjvVXXLfitkyhbLjH0tWKCcMI9sj4JS4MSwGc3nuaL6LgQoiMlXHpSkDAW
K71ZIFTkiy+TO+AGfzIYQ+kH2TdWmpa8+V+pms8MKX1InHi+yZy2NoTUhfVePtrx6gZZ9c95hvYP
OgeSf76PugYIkE/PPhSN5AULueMqHGoLAv/0nzQFCEMWapf7CErbe5kA1P06aLQlR6udKDnvhFf9
XvCUK3EGZp23myiYbLZvCklaX1pzh62n002c0nr1aktsyEzm3AqYXYSpiDQeFPxQ4NTQ3yZpmZbW
75HaIzbNt5cO9g/2urArIRrKyZeRt7CnLcxA5HbWfGBLiYNsQ7OP4NoxqkhrMXy8ElvhYaFJkFn8
8BnpmBAQHYdsNh+HsD0r5v0qGGYGSs0b/KX5AINfpzSE/Eo+uqrL2JJm3NPmJXivz8RgDeRQk5H6
6F9AUc0Znxf9fwygnln+b6ZwrOcMW9gRF0hIZp2Bp0gqz4nmqKfodiEPMkmI7ZGd2Wf2oNl/OCRn
X4w4gWrLTrkHY73aIhYHvwEgRxjrhQ4MwOkVFfhxHV9A4PbwoLd2QLUYjuACt30sYVx1YIhlvwHX
M1YA6E/jIEmttoDvCF9goNZMd5lsEdAf2lqntSM33QsvgTqZ2Oev4kpGGAWV0tmfbqYpQqkvtzsa
FYgePJNsKrXApRrfLk8GPdPajWQrLnLndVBWYpNW4z3JKblZNm34zPTOv8v+HPC8FMLHTbxRU1pP
hl9CDz8Zh5vXl7GdAmpSb9fDk3pcCCZcszTqiyiwK4PcIUaPyXw40bZJcDYglkSQPpPfAxSZ64RG
Flkr4fzV6ngIef1mctXavXMmID+gDLT2STIXLO/j7t2LcGdBPj+4Wu4h8hClwIUlTyL0F+aa77IB
KpegMmkPTCIsia7XqDvYVwgqqSxJXMGD08FiJzQplUA3TTVXOgo+Ok0SmPsAwLTEO7ZNS+XrKX0k
kz5Zr5OvCScgdw0UkKa7jMsIknBOQ2sxgB8SBCTq7seDOJNbPjb+5UiqlWn34JRovBoY/nfYKcLx
bM7f2yyJYrzipUaTGBqWVEj3YFOhTX+5OBXGPlDZAiw1dwPXhWkK8p/Dh3Kjr2/Oe/N4b/ZJOXJz
8QhKcr65UGIpbljTpnCMDYbk7DhF+cZvLWK+Z/ucY7DsHbb+oMND0lQDYfIMKcASZFRM9coWAFSz
w7D4mWbVovyiMHjQAaZEjTg/ItZrjQ+S22Jvcgnx2Vijpru6skAfZKey/jCUtapIe9/0Qt77tAfi
MYmIFeiweSvL30x7GhV2UnuwIBafPOMj92QFpMgBsuLnXgQCXeTg6drvq3LiQZ8dj6TDOW+9+47a
3db2Igb0I85mYxuSB0/psEh5aLqLOterDrsemJ99+KkRLu5BRTHshxBBmYsPCmGPY+EMvxaIXvGq
yI7ZOmYdNNZ5spdCazwm1KvRb/h11OTJ9TPFttbmHDrKmbCWbvUt3nf/+DTuGwWWvJzSrgKwCq0K
GjkPDNrGd5W1ygaLLDWSXSfdCJ/hF4ViPm4hFIOREp+NA0i+UN8LEM0c/ES8pb5sEW2on35aWcbI
qgde9jINTQxW+15nhRoJq+ypqL5kZeVE8erxy4lXUh4jY3BDRz0gnmtzkJVvSjZ2YfdY/9SNSUIW
jSItY52W1N9bsvrK1nm/yiJofEt9yjwPADCmTpMMkmto7iGAHahh/C47THL+s+NZF5QTWjVDTcNq
qxfX2WTQxBktNPQZUjgfro7yhRdhpIZsK3KV2PrkDbPdP36k+OCzxsA2TkhwKOfFbqI2bQA3jhDY
1TQ346QHsxomMoreoBHbr+egZjm7L7SHa47fyBkilL57nhVLVy5+W0MsYjtvF9M71IbWtZYCb0E1
vLXrAYJw3G4OOP667C23L0w7xEeg+HULOguU8cvwaTsPLg0swQqeXBqLjQRkKcl4jtf3Qv5vnbYh
JRqeyWAhTqbVovmBgT+W9gzqmfQ/8YSo2ugT2CiXNK4DmgmCr2gAaCu1n1ZW4MKuGY6c4S1DUQgJ
so/WuUdI1Y09Pxst/csasqN1a+9oCXtMsZLIVnCOWvKCPiToAYa4R8CYp0mFNUBFeOoTW8igDEsR
M+g9YJax+1QvRUV59ghf+hMDFZg9ffb+A7PmtWn1Xg6cwGP5lY8mXF5N3d5Jy6R2pLELT7e2ob9b
1BKkIsjDLgiMpR3mMzsjwGd0atxQ/gVYsWVol9Yd1Wp3gZB3XVXHAoGPzALtsapAqTiGhVE3UXvW
nfTzNlzdpZMcky3TeKnTD35sKiXZHi01SbhDMaFVPNfujGOMBW1i9tSTQH9nUNwXk4Fepa9wY6fA
rHaxjBSAkHtcypWL+HvgzongLjjC0FxKaOVgA497X4QSt71fSRMhecSEAKLQ8ysw+LMpPGi3dz1l
yfDp+x89OF1E1qEdTK6cEONEFkEHKm5VQgs6HXpGiDcZihBGodaamWdOWJ0crz6Zj0xjHzaO8tl9
gCVYP37JfGwNYCBOOBSwTh/vhxIoWDfd1x48uSYFZhph/bKk8AFE0Ll9BqZbLa6nPDM162UOYawj
5iEAP9h3stR2+OLfYwc9uvgZpPsOdqaW8a6tS52CQkal/917Fc5+4j18SqCwrx+BYycMhIyN57t/
lhRN/WGoyMiZK1Te1RJ1np9fXZBSsH/hdOQznwUMy0/gR8VNMmSYsQ0QJpBH2NyE2zQL6byz+MDa
Pxbo6Xc4prYGNOVOlwFX6SzWBd4AZ0Pl76fltco8D5FvDupFjpCFM8j3/1D8HsT9IyJvAM1N5gkX
eEGGjBNPX2TcXDlH5ObsVWcauIMzhLNjnVCzunNc07AH41wtzgrozu77IhaeoMwavSNSuGkcpsoJ
2wszmX6UxRoe90sc3Rw651ev0xpARTfS19ltsSDyyb+GF7S+MEANcsuZG965CC31JPfZMaMbZzid
sW1tnXKEL0H1QYbY99YsYkA/dXSGRumaJxzuwucavtRp4rd2C4q25H2UAFchw8ltn/b+QHTktuLY
sLQN+1OtLQxLlJ7Z6KwiMC34e/4qWglk5rh63+hBMj+MN0lPr+CPzmoKivYeuYHdazQ+XCIJWMC0
OErm8JjVgOPEvtwm9x7c5zX/eJrKha84O66qHhtfWUCdLIy03q77I/gAezjWWRANelGvA2/+nYK6
57q1qCw280GiMP+iwafT3td24Yph9bHKezQehiNFImuEXPGAZRGfqCgDqRxnpmZXJ/oQyWHGPCtc
IIYsQujpW8Kdrwy92wFB0DNMG0Li0/FsygFCOZECrQ+tmCPN/KIwI80RXpXvh6T5epel0qxMLii0
GhAJQC61r3UK7omax6/sxZC3vOmKuvWn6OCH4OhsWJjp6sskLTSKkiBT+awB6W9XWv6vvyTuCQDZ
OzO92zg3dl+O8+26Q5vV3UMiEquI75dBwv74Oq5kgakDQdCDf/XF+fxeVp43maFd+BxxScZdNA5/
gmMIp4IksOCs9nuscDBGxNO8AZH6BLfVphOi+z0rMKDxWdawqJYuCdwVgmWT2oqDN+Wb39rWHfvk
gzEwfuXX51NZE1LbdGBGX30luJj6qdUzuNWmLZ82j0fAPR+HQ0cK77jO0QoXUkeKLkYQQXDHbWmU
/+8tObPjgOfuen0izOrxkgDFVbNsxzFdLusgycCyWonpX7qtG1mbFCAK+Y5bhbzWSQmTnmIsXupg
Nveg3ObYj2zieYXmneCi0EL9gMw70ro0Srzu5wwZqxVRgX89s6BedYHD2zGfEn5dXN5TVkGqXMU9
nztY7jBkiGvsVweZwrL48dUxdYFMLxSxebwx8M/czP1xxAzWnA9doclUafXk5ifhpKfF+0KWbVjw
WXTFsjTWaRx22SKgrqkHS1GeDKzixvHWpU96gIBv1feCfQIt4yZtbjFFI39J3qWSHX7ymPxwRSh0
i5MvYaAbTANQA3AbHtVM0GZMT2PrpHw6dCmjWEVq05/HlWDGf7v/gPC+428SFNHiprKehuF+rBD9
pkMHh1bGsnbxbF023L8pg3hZND7TD2fHe0CbDFy5k/d49JnRy8JpVPtGEPb+aHKcDJfnIanvIRnX
qT8/0jCmGDb2cBvlt5AXNVrSl028rxFga7ApBrsNOUWy8mnYLLmVt7FBMUnd3QbR6lvzYE4oB9zm
RkJaJPcS83MZhkLOaQEFbATrQLxGwU2RoG/TM7nUXl122cFWQefT4oaCmsAz6hNvBR8hEi7aMskY
gbG0z3uEIWSGGKHeEpdKak2BcrtD6dhSKysdaZbJx5Thg6o7AneQFW1lgUBTDghbmcQVyhhMiTmL
2BPnpJkdpQDOUTyOOX+4dwIV1Y7MhH22NHFWzU4cuXEZ3978iLL92vB3qaAm7qFAn4Q0lMAd32QL
nlH9/zUcFVRHWMjmq54LqulmJ6B0ana0j1HwFQCgXIU8vSyw95ngSiw9RF84o8TGh+W+UG7Cu36J
a0qTZIsT+3qVbed5qRBS5ypnoMfz1g7x86wOQ+qTSEINAi0bM89GeQKmF5yKy0SsLXF0EY09rnsF
5i/5WDice1ItGyw11ZK2V09lJLAD5U4Xj3nGHMRPKlmt4wUXJcPo6I3fNTmpISoE2Ep0KAFvaVyR
9Hr9FmLaLDV9xtQT6ko5JysY+9IScdixr4QuTv0MfllwSoauZrnWJcOKT7VYobaLpRC4uQOCX9el
BDH85Ux5IAgAEjzUJh4LN/2fcfwfqbOGqyPIZiCH7rR95OrQvZzKhwxNoczeufuWsvo0Kjj4q738
e9+Zg+1XKY17fXQl4AVHulkWTZvikeVFqze/IouVNLShvAN7KNkqN61/dCeLPbTWig+FRsnoYGFB
oxxbWsR90emzpwVXw18C0Pf56J+KDiv3zDg+4rrIjDvRW73Hjz7DY4Dc4ZrFg4q9Y/7fBeTn0iwk
9znxr0iE+Wd9JGQFObNuGK7vndUzUcRfOcwtfJNZrWwz+3yx+cR9cA4RbhuhQuqhQ4ycyhJYNbtR
J0QAoop9dXWoY2aAb72hjCSCzOvjCuKxG+WzH9tMOeOje7XyEzANtgV9vFFX/JHQQIDgaGtC00Si
gltUCllTwBX2nze/M0Lnrqfs45SXvSmtDrqu+RUVNZRezx1zmfrOhI5sC8r5eu9fUfniZJr5kDNI
+ph9INPsNkLzZC1Qzce86d/UDMaNHId9xsPl4NvohQzOhsiQq0hcdXgqp8n6H2VxhP8sL9WNsETp
O+TF4lOOo5qYXbDDbieVbZKBj9ElgmnH231o/q0mxZsMLDLbkNFShUrlWeLU/GNHgv72px2rJL8z
C7hbrgE2aYACSQFm/R95KgVH0hogMgkJ4F4Ygf7uZLAZ4w5zajlhLZJeJ9neTpVt643huii4rpsJ
DYIvCDsF+vQR6aSSQe23cFVq4EgBKoqDaZUHtmxmvuQJxFop8F+SvkJ72bQgnjPvanMoCAx/Nch2
Tz8hjF5rlu7rGAd3b4Ehmao6uz7H9tk0SQh/XtMhjuvNAZS9YHSTsMaV8vCFEtYOiKf5K84CFoZj
/W6ZSKwMWYEu8m1E8CdSiNijBguvwKmYRvKagxvi6TrEWFPEUU2on4UAMgUYXbBAGmPyveUEQ3JX
BSw6QAansNm0oNiSJ5voqcZJW1aIUJuf+R6p1hR3jvP6nHMhdaGM6yiUH3Yf1n2HFdIVMgGVuS5I
IGeSueQa4Ey2uRYs7OMyK4MM9Q1aZGgQmpsxW/oE52oAnFeljjPBmN7f7iD+AXPEvw2H6qbo6Hlp
gPmZcyqZkLtvyJF4s1sTVmoyk9TT+J55hWpZn6PcDD1cwNw7/SsmB61jcyckIRaxOM0xNWHdigdO
1GKn9EVR1WUHMpTvi5yvODBLJdN1OKE/fkCkXivAS1d4vkV1RGIS/RQfB6ZS7Xv70SdfLq4en2Fp
UQCAYs6XtmehQ4Gm54pZcMDLBE1rOWXesI/XWvlC2BcJxB3eN/yaHhZugWSRulXkSOsV05cprxde
HxDhCf1s6IYtj2gvsRV58yf+i9hcwtG5Zgj9ygrHmcAqgHmFq9SslgoiDgskEk/FQHB/Z45s8VGO
c6YXuRwOOgFqnn+i19U8pwaHWxJ1XGaYrJ5QONPCr/v0dl7GdzhZfef1ZVQGNwllpHRl5c8i6Vbe
1XjFOpKa/rEc+NbSnfoOzCHAsuYDLPM7CYC0AXGA9IrF/vOb4waHajQFsrjQH444k9Xfr1jp8p7v
MIYtYM09V0ePIg9ctpzERVJEBShW0kruSO6X7aS4ianH9LHdHYpgnYaNWypNVUMck5/oKGubb10D
hmWuttkev3TDXzr3zkPSRcVo5Unyws7/uS9dXBzWldsKVqYg2ngTvTLNapbDLexul2odOAktP7xX
MIOR63FPBL+qwifPFAIB+QGM9+H9CNYIXnJOMd04eyVXpvlQZ0TsmWC+1rLKKz1JHy+fAGYh/Fwk
l/ppQKgphFHDV01BAxGlb/7hUzDgO5kDQSz9GooVN8DoSqksxHtkZ5JoKC+/tz5J+JizGjklQlo/
fPdZU1zTklFrjvvjem7MAhT6FAPAWNiTpoee0+nTqMRU7gsCdsoCxDcTvywcWfhewOXCkc0D0AiG
ReeF8CG+E2+i+ejS0hy9yOBHDFvoeYXmLmOmGgCzFv7wCu0vhVToe+y2K76RX02iW79c1eBs9lRI
UqG30ghhK1nS+Tdg+ERvqRF5F9XBzg/Q+HhQVgKAVQU6C9oJqOZKWdtKgQrvzN2+M9bz3+juY8Jl
Q2JnAt7VqUk4HvJ6MsNOpkW6eLHdkon3f4CfNVHtcZfqyCSp4pDzg5AK7TAUz7QvTszyXkVLQThO
gaj7b7WgmNiuk0FPl4ydBMPIyDPyqhoXiObCh68wTIrwejIrSEbE0H5YHiQMsMZVm7yzN3Bzu3XU
VBX0rlVOBUi5JD4g+af52NSxjT4qrIzIijqVK2u/LhCFjat2J+/ze+u8/hSw5ubEhCMJ788q9yUB
W+P8vloX3O3DaAFx8lqxg7gIqdXAcAZuTcYRUaQ/g5UnDAKaiPz39jNkmQJo0QZJwQisOT7EK0fS
C9ZdPoIZO4G2DbBfEoLRi4c2rbgWfrHj5cNLBhgONin3kP7pLZvcR0/cswiSi4Bzi5PZYVRK0iKx
SBH3lfh8SFL67ukheUB9LzByqokGr1eE09GzpqsMTu9OcvSAjP9Sc81dneH0oQJMUyz7+D5Ohb5O
dx7zdAB2lsxou3kKbogwXKTEtXPqTzqKoC1ryJhrkXNt5Zt3FV5ZuLWleZBzTKDPCNcn27BNN9rF
dLnqj7HY3/hiaa1jY6j1H7sZDtpXv5x08lF3cnQdnyhZSFuVxW3mmxIWrxLpUF1sPHcPaHFcB8ct
aiah0wYs9BA0/ftd5yqQ/QdohKs2gIf/C3k7Gcv1UgS3wrVmGrJAndQbYTpqxPQqAZgVrpM/05f5
8pOBLsU1jbrOyIsKTYJOmz/3sOK/uVs9X+p7CvEY+hnadRKm9k36K0N2lPw5UNXSk3u7AzhHQOvD
9ev/y+MjDBkMn6m9KveaOq0xfnQVG8ieJrL0c8QsjDymLlCnSdoFom+BTQIL/Pk3OWLblFf3+tmN
ISty8Kot9NIb8EkNTwsLjdVRK36nnYtXu0BxxE2K4+JEfxWDV9+3nEX3W+aTlHxrIC257XG3cn0x
RGLvwu6WX4uw6GjxQe12PHmGsDQzsz/D5xl3omvddEpBSFD3M4wiYLWWYIGl8sM1xsmvXzpxGziS
gHPfR2tcKceYtmzqLaT0Zq/wBqRVPBWT7wgCyYltFsZmQvwpUEOIjo7UjhvFYnj/0EXVOFLtNFpj
n7YlxNhJ2XD/xHZvRQ3V/Q/pePiBto0JecvxeqGpRC1njpjI3t3Z3qonJyHXYzYd1tlbxcu5WhmR
OuciggvHMpiHWO41+ipokylLYRK/v8HPAwa52f6Lg5RksXydntn0FPuWbqUsDmUg2fMRSpdZxRDx
XchpvlHySw9jAjyitUC9plK99oFaoKJIaawGz74MPHKQJ0B8cvy+udA8/QGbGHvIUNA79LgdLqd9
TAwyyB/XYtCAFOYiZEHYZehuULTq6QhzeDsQqD7yBn2qmtIeTsKTuHZ0/bchCHJYQYJ8AVR0pKnm
mPT5MKD4BW0m6MHAI/FhLpZRa0xbiFfcHxsU2nH9nWxMkbW6BP3OaxfHYQN2GcRym6Vn6HPuri5V
Nf//DMHc7qolBFnZJ+DDdqNALkbPNYuVzQYZ1grfYg4tJE364hNLJkPJPKTb7zmJ9MEudyMvMZSr
i0YcEH9D2m5J/8O8s3DL8TlwTqx56omWXUNLSacYCteBNXUzkEqdE8qWvMkQheepmNSGfZJQVcpU
B7y+2alJFKaQaZfRwDcfQEAWGeDvuvj93Pl7mvNmd7J4ReJpDfbqvAg8DPiKuECI6kzkQEKJ/mSM
d0StfcvQ0jDL/zaG/kUns5YkrE6F0/Tg+XG3LA834NDMWGGqheRMM7UBQ23pePvwdEezmakUmTdN
1b4jfcWAJQ/h1g7YSsMSWCS9uY9bnFPrxPvmaPT8w/yzRITafyKX8/XXwVIlFaJFgza0e2DFFTLt
LeICv1Az7ChZWnKhsPn0J4dyTomSU8t22hG8Xjc4Ia/h1JkD5+QmYFBE+IHH0K9J+OhwjnByGCKF
dwz8c1AEzttB3gaL0yGF+qVi6c3XkSljKSBALKTGER2NC/gn9g1O2Q497codRzPWI+oTT7eSG4O4
aVNxSLkJGCZwEIm50Vny0DwUrZr6doQmMqWaoZss+w5BTt9ZmfROcvGWzHgslPdIsl/x84xWFDW5
tlJL1hr8ucbUF241IB800mzHS1RPkU6ndDZcLjYaaKdMot82rCkYZUKL79xsQ2I7TXeA2wtIjHOF
n6+z2td6Z82GmZ/fBe1e7nGUQ8sDT4XuzLvCj55fIjHefXx8pAyH9GycfMDq9On9z5PPFlesG+it
4QuBDQlRfltXm9Baqh6FhFlsh83zZ20v1qJvVvVxbRPuPDFPK7XWizeUZzb1wVR7BcOMSeXNvP9Z
nEBgmNbiHsfssB9ybJujmqGKGYYiBkrxU7xSZqm7L8fmyQqo/i524CPFyIR8kOm/j5NSKvG18zC/
937bS3y2C6lzAYXgy4fVuoem8AiES/ta1TrNXxqejv9N2/pmQKTBL+ceL0CRIzqwoeyE2YDA9+N/
Fiu47CbAFIwQXPvu5pwsVNq26XsROKdMMkpuvdeVXwCzyS/uDvF2o8M3Wjef1FCLONfXz0ABxB2F
JUEU1nKMMH/GpSONKVVS3DukhUtIEejqkbVE840gInCnA/ZHGM4LrEI4UVzCD0IauLuETA1FzXfo
zRn8Fp5h2CPxOljuIoyHWkhiduz3C9ORbpVszu79GG6cv0RLsnTc5BoNovHaJT67lytscqzGvc8h
2nI1yyah/UFFJTID6IiAbaYz+cLLWxO7oAe+vjPeVeVJV4/QnKDVUlJRu38NE17T/LvBKt4aTNwO
rILJplUDoj6zKCVTYzRoxGlPaOKOr+HTBjY3UT74S+JwgQWkxRfbDlaFZNwW2TEVqHvxO3Y3A4CW
B9mVaMzHhi8HjXoThETStR4EgBHXqkjiG9FCddv0atLt7SWH0dhB3X+65WJiMvyHsWFbNxZd2YnV
zl+S5PCYMG7/FMzR3xnATWZz3InpP9ZdjgrwZuGr07N9nUMVcyEuh0hSaQaMJm3ibPQuBlwCLX8+
i8KJdmeLeploKkOKVVNEBvOJjWPIYs99dSc01YHVwli9vT+LnQFZVSh04j8tR6ORNrwrkRnWQZ6K
pp2ki5eityPRj2ezgLnLqRnlAsmfXf7XfUlO7OQumjofHq5NVptrHCRJkPBu9ltyzARswMPaf4bS
UmnQ4N4wHV27pjW66QNN23lHXe7oDS0x32x9zoNgIypJNLXeohe5YrLFxvtbmJ+DEDy6kO3Fy1NE
y/Z0P+gJjPoMMxwMo0oEehuLF/q/gT2fs5Z+nthK4WY/lizby9DQk10ZcgAeOCTI710gC3J8x1PS
7qVW23MwLxpsIuvcSLez35vYM/e4LVWUcdXY2uSQ3r8/RaqESJj9bx9HHBW5c5e+wMcOten3wYvs
N5MSGcWt4sBt65ydxtmikENFzJfrKi9TCZoj96EMDK7bDG/MBx2/oc1uIEa0K8P1jhrtobEgg9zV
UsTLepJqI1aYBTI1feX+x5NjZyE17sO4hg/eXZVg+LBUxgb2p+bQAvXAKlueOvbFDE/PaqB0/dCq
K6LGkMuwkal06T9r7r6KUe0GKWsSfK1fQnLUL3l852+VCVdm2XaO2UZZOBxtN6k7y7PNfznXRSok
DttzWXUev+DsQf2diIFC6jb8ti2L+XY3fbglN/lFo0PebLX7RAkZ2gKwTYqIXLm1nnUvwNTJrigE
JL1BkuNVJeWS9NrM3+DIq81d3uyOLR7DFEN1d5rVA6zM/Qp6J7wMpiUD5+Wp7i/Oyj0CmpvAAijy
Pn6afqjh6OAuApDxEAY40XyUUKAcQPENIs4Cn+6zsjhH6qIhJEYUUCLTUs1bhKN/0l/KQqbYJuci
q5TXgxdXdfGBFZ92UCOcMBsLve0YmZ2qEEMCg0LuUS57r4/8P9K5YiDgMlSxlHEoO7ymE9zA7wz+
qhCCXhhY6TCklcLQ2MBYCKuH6optkIMLZl0y3u3Kd72Zb9MR/4tKhxwfT84G/AZKEpJOYvmoffWK
eDdE2hJ3vAskyVxfAYb5vuibHiwNZEgR0TltjiBQ6VYgTqFNed1BAoDEFpbqcIOFAYVQzOMhDn03
xGF/I3mYZeVOyK2B54E/dOHYA9qMgnpg5jeJjTA2rusTNC4XCbnRqJUoH0429mP+u+0wePjfSPVY
q1Z6UqViRlPZq5erpsCCFEZQmrzw51ROc4/1Zv39ZMNV2xoPKqP6hrEC6NHmo7f3a1nN5C2mZT4e
OsEiCDkbxUQ2sPeO5V720I5r4qBOoe70OA+4Ft4YNQHjZKV/9QokeLNSWhCRSaJMsDpfWMSk+qeu
KLHMOWO9VHJgmoEkWJHJQR6uGDeyR5KXJBfLq2uU9K0bOiTtdQGD2jfj4hN/mZEsK+7rZECM54fM
OpKT+DVbvMlzWhGlD2OmsThbRmKGxnXh/Ezy5NbNZvar1hAHLJQxW3Ot9p8ig/s5dtExH5XQmGN2
9mTq6rj/qeCfm2+AUpywtkjUirzgGerjOA+FkR65BOXUoGShYZNezbI3DqUdy4Lycbbp8lwQ4yx9
UPbxZSMeqjK598lBP5u5ERRyxOKs/LWSlt0iAkZpEzKhg1LHrVOgmejtoe5ij884mfoBpZQhidng
YxBGmPGIV9TU7trnI2oxW1NsgoJI3v3LvtpghWqu6uajmTMquGXzS7wnYilWOWCtmkK5JQBZWRsf
1KMHUIr646Ovy1XbFbDhKSuNj0VkO5k9BWEiubIk/05dDxZL3gj0XQ9esoclH354tMaCGCPOCAuH
CGfWIPEAeNrejdn9nOBM28eFU6TY7EdEct9UpuJ2aCKQw81dl0X1ygx0WO39DgVHLYAI13vGzATc
wahMxv3gr/rQVAx7e+te+L0oq3twTX4IOPHEhF4UlEarWzOxXBx0GB6PriRJrkhh0Cwy3JHZytqC
LYozSjAo+dhyJlS/Xe4wHgCdq7J6txUlW0l0oO50JPJWJR9qE7qyKaYQyNHmLZ1GYRxBqTxppG6W
nYChuKLZ72qD5OXBgmS+CIIhB8VP38Rua0GUKWEOtd4CV/wLVdZZyXvSYbIvU6KVWWyeMe1ML5Xw
k4CbgGZvScLnkXEG5KOnJvtLdaBpJU1vwhNYFgPTTOB7Ow+aA/MbF1kBXQ4GJe/HEM9HPsQZ9D/1
3ntOWchuQBHrbLdjGbWxt40tzdGJP9+0Vv8D4RRDANo0K4+wl5O72CnZUNviojKhTnadOAcuy2Fg
4/8yuk+iwQMcfvCnlzNGKx0dUrV+fl1ELSmHGNHcW3cOu3p6eL1/UajtD/sYPROsFSflOcxXlMip
BScv5Vnc+1gmjh7SK7xRgnt10lHhW5gU8yRYgEqXGUq/qEOIP6BqkKXqe5bNunKWUER0hoTbmNyt
SWPMFlP9pflffb5B4ZP4NXd7EhDSWHhWmECsnfQAi3xy7Ql0+xShSEu1Xi+b4/tbg2KGeMGkLGn0
+sHFTn3sUUmojc9ZIBUvzduqqDU5Qkt83LLiVEGaTDxhkKAzWh0uD6ghwUT1tkVip/FTUP9xHiO3
e0uua7BhKnvmFTWQMKxODnLEoDCYpM/0dLCPhf4OUwFgxXwqLF8zWMbjDxZg908rURvwXmBq/kyu
n/REsIxWAoE7tn+eRH1kWiaMlOcF60+ZxDJxPczjCkWjP+o9RqEgHlCDglMgyksic34Us+YSbE/E
O/JxcDuQ1zfMZU6NYksUsXYE35bCy/0kBhKVsLL0s1mVYJQg3ikeQak0iDSwGF/WyXEZ13o8B4bn
ATBOWHKvPO7pekF6+VakvOZDwPcM/prg2r498nMq8H5yB+RhhN0unmCqMlTnAYJGposiy5iei6Iy
ONNldz0G0HuJhooNHOjAaTkKqSpkmwiL1uXHUmC76v3XWEr1V6dzfNBoEjBMDRtnD6YLVRJB3kk5
T5hIK7fJmRess/wjmeI0IzVqR5RrPRjRjXVD4sF1jxPkUaBf4mOjO1XgLyVA/cS0vJ0jStqY4dxT
omvWaE3M/n/2uUpblOoNf5u64EzG/Oc479Hcbc0aC8q3EOZjpVUTM3vFYPG3Y1ThZ57Dn+dkm8v7
pP/7A9/qVTykvd6qw4IIkhSaFno9imCrUElx/KPQeLVdkVxfydpP6ih5B70Ej/Xh417/cvpmTNkz
z8QOunBmFEO/vtE93DQwFUm4Vadsksw4h1g3B9gJkCLUxiG8Nc471IOzdN5Ohqlni0qrXt2aUZ6D
UKffko2sfPK8rodRpwfbv9TDlBdWvA2kqOm/iberlk0dSgPiW2xusQ6g2/SNiLFa41j6cxtgbQJx
CPrImSROO5mN7S2JSUMaBof3JFiR4KVVpYC3kirqv7lOEZgR/frvzTW4yTlFdobOCa3qo9kgJt8w
KwUZ08x+lHX8BXRWPrPBypTFRc5MZW5PdnC1pKjRhWDSoJSLkUrhuAt5mG6NylhGKtFdQxpgp117
513D6InfhqrkpY+LEOad/uEDFMsxiOzL+AToJ5dnumpybM2ZjpB7kAdgGRWlQQefw8Gra5LRtJj3
xMM5EZ2GuKRBS0dNFZqGcRhOPfUiDUHGCQcIwN2aEL8YPbDZhsyrKlk5qxCaRxiSBPfoxkIBWCSU
0kFf6pex55Xsno3PVLEJRFAkhCwIuHzcT4/qS6ywQ9URezdD7e1bSZe4sf9zOnt0n6jtpvlWFKtS
0MMDUEBxPk+ss4lBABDusEsP6NvdKILfhfvKycECxuI25kczgPaNVHk8wxlqVqF8eCzzg82os+dp
bUkFFu1h+LFGIwv8aYPLp5R4BgQIs+j7PRPCUlVh8vc4r3S3apg58g7IdB4tDTYjtu7AjtlFsbTx
tNc9PthHxjbTxnp8dfCQZrb9eeyAeGEgAFOOodLaXWEj6Hy+/6jndsx5FsrDNi8zICMV+sRyu4yn
oBNXAD7sRANBTAmyWMV9eO4Smdzcwy6+r8HYC4JzFLO1wIZrpYx959d4M+BjgHtMKd8ZNJg3YLW9
kRGRO67jjlNdy4aDFhzWR6lmUbUcRCNIny1KP1vz88YTLpNLNsAn5vvVNxkTHwZgDAD5WzTJQk1X
M9AKq91/QtrJ8WrLWRBl8+ZCpRrK517EnHWDFDzRVCn0hEt53Mm/FXEJPKTnHE/nMtFqDVbikI5f
NwWmfWxBTq88rSyfGTYes94tAQbG67sVkYcASJ7pBkmQPYIKs4lilpQLFM9+vbw/JNL/JX0BpKuA
Htfh7Tr4KC2XTjx4euG1xZE1YeVWslN84gqEVNiXR16QoS8SKw7zi3bpYTZrfPW9g1OHmxZlGzqS
WGOHYhbfmsrWMsClJCs1yM/QXNb/WXIi9d4zQWPUabS17EhGYGhZhrsa/d0bey0TlM9uXnr8EWFR
nCZb0KwOplOlE5FjmpaUptkfIinwuQPPL2tPIjAmtEVqsJGG0qPqgfJ3IcBpwwTg4lZl9aKJ/cBn
P00JWjFmmSy/EbblhA2XP0nu3PtKIEN8xcW6dNTy6QdEXocQZO66QX8yUqu9dM4Q/o+2Oj7mjLI5
PAWH22uSwTlbCHQSf6rxFstcLrLPL5clD31Ox1z2Cxo9oAjw29xEYg50z0XhkbhJgey3oXd/duRi
9uy3J54MC0YacgopHBg7WqsKxRJC/2njWAe+JgfSW+UwmBdakfz8EcJoeOnlqgpEYsDHAvQyh2Sv
KqtivR1qAWOxpLjreXCuYzSQQngM96JGnL32qYaT6XACAqTZ9wTVgAY+91EN6nSOcua+MIKaCOdQ
HZtaNotOPoQmeKURsCj5kuju/vucxOngVMICxVd9R9VY+2NqWoaKBR6918XhiPJHtTWnGFAXBe4v
D4yBelBUsaJWm4NEaoMd2qMXVlHuJNAdwQPWdFiKDqpieLDzSVR2Q5wr4xhCBusU7v4xqBZ1bOql
dHVaWWLxHegIXgnOwGhSFGbE+VTVK/+suJ+h7q23GzxQ3kQL9nRwFiLObK8NFpcGgi6wXIn062JQ
Cz/J1bgb2XRECX15wWrczMbEdV/PicXZRb3rSg5eU4YbSx9SyqlBeK1LkWAKC81CqVkKXcKd7Dp5
m6rGgUxsQoupl0Jl/6GfbJz0XHHI/t7MwHj+9w2GWyWFMFd8T2DUeOrXCBOgpTviZyu0oC/dtRNH
5C1Kv9OYRhHfQNhf8tGLicfSKNvOgTg5G2U40yXiW1CMVtUyAUTZ2WYRkLQWcGuPy5UJ26magfxY
vkOGD1nCR5mjAwB9j6wndi0ExKQF30m1tj3y35OkiSsL4WfmHNufChKF5Qf+R6AnWz5SFz4NJwp5
B+LvQugCbspjutTVn8P+U8EIrbty2l47CtpPsFX447ta+pu7i6dk4axxdU5+H9opQLtPRJosozgM
8OfwH21nHLdVO8h0jOiGNly/DTYl2BI0UPJAFHooLjs13XukZFWSU4Ke/LqPqBndtS/k3zOo+EEv
SvW3TVvGrfVWBUAuAX2svA27o72v03vPQfoooRar2ZuMO9/Ij6RH74+u4+DL4+qTYu0S/Jh9MiiY
Bf44eFNJGiUvJ8kZetzr3IglAW/q+3APnFAsyiPFDs4FKa9HK9etHG8XtHoUZbFTgiQ+bJwPxJg6
+fYrEpZEJeRq38arNVdseOuG8u0MQgY8/LhaoMghCZ0hc01czl/SaDDKg6m/iK8w9p6PFJw035eJ
5ZJpke26pohdIlisfyAWpOWTFTH12GrJgz+QLXTrZC9DVS7PhwqXoIwMgjhF4MMZm/FiMVufYoiy
i9E8ZGJMnuTzmzTnq2wo7PxaghB1zy9m8B1kVls+O6OCZwBi52k2XF0F9/SEIuUbb8H+1Q2bWmPZ
75IT4I5Vu+zhZvLqSKDRvsWERZcMw95J5fLfr3NcU/kEH4dLHIg/YcKOaQLaV9HMRKXDkWvYoCZZ
HnluJEV3sQDC/d1oDyqMZuV1HKAd7tTleQpLSG1bawoHWob7EdREEsN/RG45/E7wPRSb/cp6FcIb
kZkgkkQPCIaKC0s4EL4FjzOSscwXCxgSZs7GGqqvAaJ9tegLRdbk0AaZGJty+eqgOYq1Om84viwu
O5EadeWMS0NJCcIReMd2geUIbrfF4JbegQA8MqXmzM6baaMz3kJB2Qd0B7Jf3YL7o5O+Knvk9AWk
bByDUCh9NowgqLgdgJxWUzgP3nkleahK/q4/CX08BBFAQe3RXRhmMD7XxWHDUjalEkF8chs8W30j
0J+FWrbGyTioxsK60QAPIb43QIiSiKoBkR7Oewj3a6kyQGpwr33Jrn8EIBEOn4y9XXELooJja2HY
2OKOz7XC9K4UU7bh1arkArUW8Cjkbo26aMywJl2+VGaVTsg6jAtcAC8YiXKldWXNRA36wHTG+MoV
0HSTggPB38q/4BRmIDckySMQTJv48F6zxXZEcom+4szkkc7T7viU41EUluvIny+uFthPr+9cdxTU
oLeAOIId4Iz30/pqAZYiO/q+pbGRNKYg3+NFFeL3EUHsCSuj/vRHyLN51+FQYYB3GPLEtMOmt8I6
cYlRHhERlFJUPIy0ZOM4oW9l+3lp02WeH8zPHLPWXNxJMtn/V0zeayflZrQpiE9MCsMzQcmGSIGf
RiDAhHy2fBZJdVnyUnw/k7Kxktz3UnyWIl98CGUKC4n6fCFT70gsvCnuqQchnaI9rL2s1pniUPEF
zcE728Q1sUUeZrX9oMkhZyW8gvSjb167fG1cWiZ6TtSp/ckzxZJltvg4NGyDibgSh2zSf/1rvW1N
MD/W8D3X8InoYY1Yt7xka5EN2JI5xht1eJYZXMgPh4P2sNnckuU6De3v6m4DMGwI/Vz69Asai+82
DEtOS0YbhuGKFpoYFeUsOFKtwQ3rqg7AEts+Ds4u/EXUGS6gJq89ac20xAp+oV0ipRxZuhhwyW6C
0ygAQYChL0Zmk+MmN5BxxuBl2fJCbOChmlUSU6bRsxltgCSBz5ohBJB6P2/8VSLRoI9YjpgTReHK
Fc9ygMjdgFFRUWIhx07XtwzghKjMfvBG8/PUzxmKn0ctBicdSk2UV6UC2WIgDK5ItMltyOVIaaGC
eqh5jWIhAXeG20EdwFaqmym281VBUBEMlE8Qcr4dGTdFv87N1h507BGIKp4ZwJqUm+XqdzLoEaxy
EijyWYvo76zQXWGasiTEN4tPQJeAszMSxOAdT670o5mYHFNqQB/cw1meVuh2yRo41xmQYgEOO6rd
OMkuxqbhh1P4Z4/YsfVkDQ3Kb79mSok+qrQ3A+aEwujiFCgBgn+d0uvfBiqjoL8jlivX3VavLhpz
4OGBD0Qe+YA2Q4nOhFjH59WDVLqONxWxjdOMWNOZHvGZ0aeJ2UMXCkwJ8Y153aQ6ZL7Sts+K2Kqx
rz2TkYWJtwFy0P5XP7czIVJyQFV5pLyDD81pjfNCXRGX0xZyuj1+4XoIfe1jhWCJGi0Tx71U8B+m
MjY4sg8LVTCrSpvuuFGUCHhmLmx+eg2KzZVv+0nRxGXpTzucHYCI3CcOfcF4WEmtfpx3NCGYQfYW
wmyYjbG6YgqH5n7Q5aTszDN+hw/evXUX7xwFUb5gqP4/nN6olffLdlBQwc3qM+0qXDzLgQqZZzXE
jLY58jZpfs8MP//GTjF6paZW2gG0ZOvR09vQ+7rSIjCyueK/5sFYOpP2p3cpbuIo/dh9xvsIKl5R
4MrSDV1Yd+slDHeyyj9iRAq1sRg9QZij3GbMHgeGu6I5WX6xa5SR7XIU77qNV4rTiyCGzxGuvjlz
1Pfw9vQTlWE0DS2REvOTUWtwjX4pUUyMvYz3Kr0MVpMcKffgzPmPXAjHGhlz12qah2NbQd4SeCNs
RgEy9bYMS5I+drR2CH9P+0jvNPH3TEFs+QdShFYWjqR0xRpVTlv3QfW29CeAXTB/W9EoelGVa1m0
K201j58XIHB6q8GdFHeBkuv2yMy06aw7Zl5fWxERkJCf1n/kfFvRmfx74sF5jwBHHpOaFQEGGrGN
2gYaXnw+LDuinVe+uz19oszeh+bG2asNJmZMql/ieMVC0VzQfK/ZmzA+CpwG16O38G84cBv7qy78
yDrtVv7sozcMTVY9boyUwfGWHfopALVozdRBb59+iPOFzrXbPuFTnoBRlXU6c9TE7j4vQQTcjcz+
WtowGlLEYPCeeUg2Tb9Dg50uUXjJ+NSPcuNBsqE/Mfpv88MpiJYp9j6C5FF2JUJW1mObsMmYY5/C
Jti7Jf//CXkGbD6M1eEGxoC9tabcj4WemL3skD3BdH+He/LkwAFmCKdvzhNPfckTTU4DDWBENc8D
herHgn5jMmWMTO5LksH69kZ6EZ579NKOCkebmBZflayqlmtOEBNEJS7xPro4W+JAt9u/6ghUnfLl
wqRWgsyjoLKGYVvsRs/4eUwCBpVtho/2pu4OXgmfSOFHqn6QrJUYfbVrVoONSW/S5Iae4sUHCoYl
H/qEHRA6Kzag32sEUJ82GIwjNBgAu1y5f2H3HoB28frD6DAkYkNRGDxPXUWPs/ifVLp2EXZ993sF
wRZ2HBZrSjWbFxFsvDtKBLWYXuSQzaVLAq3GGcupIFHZKfi8Cz38b/31Ywu3//5oSNGQNn7HoeSu
IlqWMx6efvzvwfwaZ7iaeZXaSNpnjo1QmXn/BqWTd4tBlb5mKvcbGvAQz6UoZkksZ8qRMSu5YiGv
lMv05J2Mbum0Bxd5hJEasSIpt1KFlxSlh2cXMKViIg/XtvJo4054/gynWM2rOY8qnyTEYXpIjcju
ZuljhzuP9u0oqQfMNEcofIOvG7qxEWJjY96piLOKPwCVyMwRYab1JARp+zNDuo2KYTJ+J2wobb1p
gQOgyHneWM3JpM2pyo17VmOa/HImkzxW/PydgIudd+eTgsTitLCpY/PmlnUdPW1l/d5qnz1uDNjy
nePB4GN801/IxwnQjEOfdnrfCtDlfLLw1SUVE+80Uubw2eBCTkEU8mjf2Zuvh7ZkCgcOitev7PCL
Ci95et1QsVTiWOdLi30TCNXQRNKHyu5DygGwo3QC2RDV6V8IhEJrp27xV3J9LzUwp7VqeCU62IGk
cii7wTbA1y3dq4MiFH6mIIbDnRu+RgU9ul+VBZ5Psm+RfYH1PLxmyEZlfkL/ryJ1JsFKi2dg3/HX
NHxKFWcJczE9ONvru2y8RjlAetZTJvAIE4PdHxjWAjplW4jPTGiL3IB+ksI/SU/7HRWRvdc/1uAI
WC2ObU0p5TsrTokgdEvjXY8MGS140jPS7OOGg9/gfJKdQ8TCvLyEXt9nIooSXVNY2eQf1di56wp8
sTOtuzFGSpbWDWwBrPLUDK3i+C98pocnPQUKArkeV45QHlY2d8groWyKKosCYfUbsg0KX/mOChc5
nw2QoxEkulFFSXLmsAmGv5gBqH3dOs4XQVVJEJsUfVpWOt34VA7awfd35GYa1Hrpu6ETX8Qlyj6K
Or2jMUrCoR8dqgydQK/SPkhJBkbhhdP03ko3rwxcefR0bMXvH88Is4LCuL9PtL7lZuPL304hV71o
snBAhE2Hhg0I61AlYkdZknstGvv/NZPVnJGCcIuv1Pdg4j6bhCNkUOVXXYGor65apQJDd4EeldFj
Qi++sSlDWPZAvGdUI1Ko59SmQaPUQDelK4lW9QR1zb6Lu9FRRbMiLBRriPDwX5Y4/mHtUGrHGlgF
1a8BxYs6x22VS1oMfokBIp6P9/kt5G0US8sZl9brXWD8Mi/vaQlxZr9aHT0yw1C+E/aJrCVcMZjR
TctHJkZUh3Ek2ENR/nugTkc7PIxbmytV1QxEVZtAHlVza0v6uJJ5U51QGLsJPTrA4Fufnq5GZXbb
U9qOjpJreW95Dkwq+K9vubPyNj68rWw/3rh5ojV3xRkoMvLnKt/Vcfo42b4NyOokBbNQULhEIvl8
D9JMuxL4ZT//PdSw+wxksqwHBTTSqsLEMabm3fUJJ2b5cgffj99AM35PRQZKA8U5XWmsDKy35X8B
EucIiQl01cc13XpVQLqTq/a1A27tsGSk67YNJkmxw7cmBJ/WypDzMBfXVEvA4JPj49wTzP7F2BDo
78ESNg9rj8DwyMD3Mgg9uotsCbqES89OASFtxfDfVpLsn5m2PjoSINZnFMG8MiTEDUkSvPkgvNi0
tChM69M9G8+qfxTFmbr5yG9Ti/u2wcJKAx5ILutv9UazuOli+pzNIebBIKXtDfLZ6xYf3u2hzs4K
VHrKxe0gyrYKOnwJhgVLiVPyELlHup/W8xTtONkZCbZNn5MOSqo8la29pH3RCKjI+3QG4wknFpoS
LC2mRCnmQsSaGL3ZfBLh80JD+zov4mNa8hJrW9CQ9rSXznrgxKcAsCNmE7Xf4figGIoroLhSc/OX
+ONKyFax+liBXmNBCBSCd7qgWFD2VU8UY6atG0s97azhd4f8AE/L1uaYEsnDDVNma1SK6Az20Do9
SafcKEdwBmEiV2ztIrkGJNM2qAYVW7Hd1OwpiYrDd939HkchPBqLy0rU3Zw2hlFU6vx8oPhen1DU
pgHisxeZfHV5PIgfBex46BZy20iI/U0MMFSj4w34bdQi2AF5hiqRaYTM85hbuT7jzwklz7zqxsQA
cGRFQraoEx08bmYWbpuYyp7JJUecfinLmVmiUjP+ovPGQU9qoi+5CZu//PmgJx4mO8/CpPGKADxB
FRCZdG1s0/R0JzCrMt5yuhis+YDQl4bVJk5zt/n8DsQ/xkurRS/Gm4pSmZ/vE5055DcL+Tr3i/pp
QvoqXgiLw4rLmsC8ZUGOklERg3sdjSvAOG7ox2XCukmkCnoooStO1FatgnALE7/lJmWUDMM1dNno
v70YSD03YRiJU0oAnxablqMCFkeahhA1dBOCrk3YqIfa0zZc1KxMQt/4WQoGydm3GurJt8QSMx2+
w5x7Mv9ORrVR91AAduYXYFS2UTM2Tl0z3fHAWGNIWse82XIekYf7wogBkFyCY4UAQcAIFPP7WJJB
4HUbSeofC9z36mIbHAhJjkahqhMQ5ZCQj9A3gmJMWTWdRknHyoI9FTHTMOh2V+Pk1y6wZMXQ6hoS
t9VZbrocD9WYIE+xJ07ov1KGrw17zpWlHCKLrJ+T9TdQr1MTRpAb44yBT9qJGTyFA4r8TQ3x3UoB
tRaD76B0gd4YVcjwPP+lUg8hAXiq8NnbRkxKjAvNZi4OoXOywfuGYMF3uXpggnrvWB5sWiVajIsq
BGix9IK+0/RvNt1r4/RgnyAofShhpeRbuNiNQvneEtWOq01hPeFOfsLJF9YVobNBojrO68ZpwuML
2UADpUCjee6EDN2Ed+aVr63dMODCAbFtNO7+nlULApMZyRmY1bsMyuuUH3/ene/RzDtx9P5PETqI
x1X+i/VED4rm1PxqR8R/nwP95bKWeaxESJc3my5wMs+wdxVE/MrIdkIJBqkVeNvu+hBZgeb9oMDT
K33UJnF9wA2b3lrGidsnKZr1cNwQBsfZRxdE2Kg3VKzZWArImcSHP+n7oqG+SiNiAepHoptqa/MG
yABjn2KxS3fonL4pTxv16uscpSyLZhyZEJ18SBjMl9ZuM0XyclhzMqYPozJLblNXP2dI0Zi59GED
/H4q8/nse3i0Sw6cdQdtT7hTvHcOJicF0x27B9QtvWSs2hLjp/5VJV1TisVEvzNtBMF+wGJBgUu7
6SRtMYx3BQJsj6O5XiPQxGoA1RMboQNs6y2hQ/fW8cqPtCUpOW62F5TlPgU0etJ5UxpbOISu2xAo
E9Tlu/LsoU/0bOwhROxUP4aDddcGUy3pU47KEhiTEoRndw7RI58scvXMfeuCF3MTS0AS6bNDpslp
Ea8clENN+VQb5IGo2QKNa2n65lPbMkTQgBn+74Kfu7XbioqAbmp5th6DntvZ35NlWNhZPWDcZ/vj
fqx0Lr9apJfmveNYBvlPZnX2P1ZZL6K+KqgsXgiUeex885xWk3QFFI7UwxlAmVp197PUoWlcyHkC
CtUaRzxLFQTau+23Tvi/ZNPxW6Dc203/h1LUJ7cVGs3oOnqA6KUV8+Dte2ncI7BMelK7zjyN4i4E
XyFM6MdVt96EZgGzGjuYrUpLGwdZDedvM3FYX1enH+s2oA/JK4LsO6YdxH+gNCh5Nuek1cFdYD6R
F9BHCnyc/AP24MFKllylCiOi+buLQN7wjF7tGByl80uK4LO1+pwEAEabw+zTARBXnmVUFaBfxkoD
j5VmXvQgLwbX7Nfh5vrBRxTp2iqTIvrpep4k0zAzsJ3EOwBd1bDncz8cqYcCL999J8/GTI+TdzdZ
v8XlK6YcF1LikgD08iH1dsDpKdMxdvL1Qhx53r3ydwjwWTNTLjFuHRh068BjBc5EbiToz7767XEo
PUcIXM79WYbrw7r7qpuH83+3uz1+k6SW8jWwxdisemsucWoqFTB20LXp88XnAZXTnF7arWCF6V2l
BOmJm2dd2g/5jI0P2nNMqcjjV4ygKP5IwpYNGX4GEe6bKBe72o7BxU8ecXnTjrR11vlGz9LJFe9K
BgCw9/IAf+536e69WKSB4ve7kNkEdmTNjF8rygtIe3qXRNBWjQJKEXh59D6ivC+7zfwjKDKVnCrP
YwDzFbO1C5gwH3LK1X5tMBVpVGRFzt1vlkujbocZZOysMEZI7bae5IkEL5GuP9AAmmGR+6I3wqw3
zLIHcXLEoaVxi8fqqDUBOK1rH2hrpr8uZ4944F9rjJa/l55R2qlFLtydSMVmS/ibSes3e9Ivgyez
Hn0/cqoEODDIi92STroYbZpUmg/7xLXitYg/JkdJ9O4OwWO3FrApkInKmpNZZwkH1WVTw4qv2185
zrpxdAn/hdD2ekN6mUnG3YLOSqsu0Ae4WJxNf4Xr0NE+xGo7lX0Sbl1OI9PyM+mTBKCMhmuR+eAr
2x8a9ZvxPkuvvjQWqKF4OIOBOdTQH9y/jJtgYV/IxZmnM8fhtvobTvbQFdiN4de0KI79ZCt7OF3I
0YaOhCp+IW+ifnQvxDepiwoOMTvZfWt8T+QCmWX29+CM46BGhxinUdalpQMkmAZuJrpLQwhUTHgA
Us9jnp6nApkPUJNUsoikjfx5Gk8Qr+R5tTZJqHF1Q5u757zpUL15b6fJZDoFfnX3hE+QBCj/oIqn
PUhRTPDd1oe0BV0WzR+xWh9zKPl6Fi7rap0PoPlvUCOay3CkDHvGBVdhgj4kWUcQjFaGZK7+KvPz
AFhVOQrWTv8AI6/KufYf97XzxID0Jg+I5+H+zWSJJNfl3qDeqpWeYbvPvYddy4N62JTiifdFYmJk
+fdCajan2P4Vk2pU36d3JMF3jo8vZQE9WWLInSm/RK0pOYXGtUrRndI24H/mY6fLldcbulnIJCi4
OntPrsbLEkK3HnwdPR2dNI3l6wbV0HC6lTtybLxCbfYwQQhtMdMwv65WjotA67Z/O9bEz8R7QFzQ
2AdXJNYI/sUMd81GVgRfnEfKr7ra3RYctNz5FTpNe2MTAs2g+kk5/p7r9uxbQBJsmly+K40JfvAI
3HSCEP6tBY0IHCitkpEkRt7be4o7HpROrMtaYaE7C+boYhy7Gcgd32CeZ1VRU1KvUTGN1ubdRGFH
uab1j3+kLIj5MnmPnyg8jdB5Vr/PHzbWnExm2F5NvfaswREmKuvfNgSBwMf3enWtV0XNYexF5JG0
GtZfEjdZAJWVoeHs28wToiqSCNkzmW3o+uxDFIEV16z+k7H2mJjhjYEqcy26hH1AjMUnxis3UabD
AbE0xpmUliYRQYT7NqA8EPo8ouBns4kIN6PWKdrBOsjDa4Iky2um18q5Gncf1q2FcWhQ7gJPKKS/
jNgOLF+VgUQsOpUU+VQvihADlL+/axYagHQf4QHDexH7UuLGLozKKf2l+Hk5iXaPg56I4ruzv5Bg
43Y+qb9oiRzQ5hi/Qw8oqtW2+jC+KwpovoaCZs1b0miJ53K5sSFkkY1zRPhIgyIuCipZa2mwJZI4
zh4si9KNA6JPnGKblz7ctR7vmGYcjUvoK95zeme8HkB/BSMcgWtK2DJ7tB/21cvVK6PAKfx9PJNG
ywvlpi38mw9GjfEFFib/ncW/x5LHq1d22pAReAcHYocZ3fCkRODMcP63owVkCIdEHhAwcu6hGVq2
2B0DESo9dSdtCSzmOjaLGOeEMkFnmyqyre1YoyLyPTa3aS/d9Jr736boj0G9Wdsgj8C7oIt/aaQ3
MiK3MK6IjtkKQMj8uxex3URC2W5mxda9lcVyUqzxDSUMeUixYTCp2xKVtKnc6zfo44ZfF7z1wK3m
YZOte6FpfaRCNRavWIGlPLooe41eXp9IMcvyDcrQTsN/mNmGvX2DEUvOmqzFfr0FRN2ka987OUd2
JaDzrg319dKtnEN+5jdd2/cYF90OuIVFZjpXvyIOuRPnESpK+LNZkSKQb9h8LnP+0pLYnBu69nnJ
XJRoqTkWyEOrThK/67iSii9HV2Z47pu2BCsm+OGzMrQnDwW8DZwsAhUxyNHJ8c1xk96rQ28WjYRT
J3VJ4xV2YIzpXhKF1KMXz5S9Afy6REbAdHAzur7/HjXjegGGGELVsJA5cJWH6QcTIXY27D/AGFEc
NJkxWD830aOirsqJPFWBcxQFNi7Q8Mn2NGMnmYimj1hU0QwOe6k7bMQhUjzWRPkOn4z7tzEJtHGi
l6StAUL3ArqLFUChveBlhEMtpiV+hO83d2qewh3bdcbj2yfuA9o1Ue2s/rvT8aAmfld6HtPi9YCY
+HBD8dgI8sHgOT23jtvkwLNM8JYqeDItkZsb1g34O9uSmp93FwoGf/D8IPar35ZBy/WoC2bRwVot
8yebPi0u0k1B6ZsOr+k+unenOo8sfT0x6bvn4wTaTmXG3DAX70fzOnVoOt3BET1TZYi/FngktvJf
IT4lmqfN3tgCdsr4shxMziUapuCHW1m0/JkArdd7GIVYcekOkaHcPyz74HUWFX300tImmVeQ7os4
TCUWkx/YIEnOTBl6+eTN9FaMLAkUZ1+WmEKPoBscV8AJakVRQlN2AQsL10OBXFA0l6xh2bAw+o/o
I2HX+eooNLIiya8FogiTQTBhpM+xTiOSVeu49kz5IjECkNsAyKn5KlML0ewRwI6JlAs+snyn9TWn
6uyDD7qP3Y9mVGlDaLL49GWWWZmd3fWOUMeXsfKbuVygl6r3KsP0mzGFtrP8aOvSVKT/Ltme9YqE
J6p7otYZRoZ+y1eLyqDTiTWeKxK2qHIb595M8aNowp7UbJE+H+MFJeRdcsYaFb61vHraPK8cwQu0
GYQdoTRzkhF5uH+cRGdllhhHmNcyulAGaDOOcS4xN5YW766oc+YJ2O/vsW6V4y7UZ7NISBqBhtqm
o3M83ONB5eePwqquCBS3ZppE/R/pht32jKVhj4eXDglAaMBvkF6dVwLyJQpm2/gu79Z5ZFxq7jjg
uidTJa1A8SUmyhVd8touXu+cgY0BrNACrC/RFTKFrNs0D1oRW2JLCCscqhiM4P/1Gg0oxHyAoeaL
J/SmsNivftf+N4HWWbZnll1UG55CtWVqUztSp2phbsBtcXGj+8uleVPJ/ps+X5ElB8E1YweGtGG1
S1blJFQPfAm/nYw6pjJd4YAXNZmtDxz22TfPdkbKp0WUijUfM5f60kLetEAtp5xyJVIT/zTHdFyy
NJFQpHGY3ddAc9oI5Qo2HvhhHdDLbdbJqnG/SjFNdKBZzV7+DGb2LHKD3xSwYRnpn7Ih0NcWJO9u
nSnmp3AdLBdMZx4b2ezs4pzdFJwE3YjVscc0YGDUxkEPtHH1/sv7PPqHEHYIhoyCyPTe/V/YOLtb
VIxWkT8VwMR2Vy+i7J/WSizvpEfw+RRNd7TcPieLV083KWfn5BwGdVMqnFIxYeFboW7WhRUO6j85
xCN53l+DshpygdviA8aNzoOJW5cWQj2S3jt2n5Vm0K9qbX5ZxMtNHFie7txWbSD0je6vBD2jrUww
3Hy1e1ndykO7EHA/WLx0gAY8Q7Up0/xhJyY2ouFFywrOkiOz27yGfvWUNjbOtiHFKCNC8o4NbanG
dyC8crag7lipk2ATo1j7O1gplBwG3Ao0oHkFk1MgDgSl/y+4jdBFOE/8MV63UM6Pplt7P3dDSPFn
ETRNNA2UEzl7JqMIJASlUwkADuqKx1BV05zYNWiBt9mOmxVkSdXjnY7AxA4K6EGF32A8d+aGf/wB
eArakqtcoOa6avn0Z/3hi8HwzrKdWMIIniejxdx9Eqf5AXG9nBDV0C1djkQTC2sICxOCF3SJJq56
OooOxAQ3/ngC78UXw4r/PSMpJqts1BswpQxdfpi2+SG6xZptJ2JYCR4sY7yGvNXbLgBBwj7st8Gw
9JLXLzCank07y3wYNswr4FwSwGHiIOO2cZKDosabY4qRES+z9rIlCqhl4SjHzimpWWzpBZu0zY0y
Cf2Ki3AWC7VULH/6uCp1oJ2/hXc+Cm563cbGCUju/DA4ScNlYzbKZlHde8ciccFuI3YgqcDGZqZI
9X0VvQS3u7giE2btHEfr5kd7kcmlF72qeD4IFO3mo3kC9yMGoAJn/tF97sedOeHpI6K2HO5TwfY3
EZdd9ua1+gqZ0mO2hYXgK34bAytGSgn3qMKd+3fk9KEKjs9ekhk9qmcQnYbGfxf00KaWV7qorZlM
3XI9NnI0GTGRa5B/mCIPZeTLLY/R0nXWsgx6bh9mMm9FC07LMkgy74ku16JPZtQgV0pSJO1Ym6uu
oK3KOXv+bcXe1W9mOFXQFkRkzEV+3TUQYUWvj6GjNVa7xetjMzjvWLA6ltAwiqDUS09iXYd/3Uu+
/xS43RfVjCsucVBkWYfuLy/BMzr/1grcvMUDp3Jd2YBbZnIGS91fQOIxaCWrTh0s/ShQSVD9fuMb
ke2f5iFbX38RGjQkOkLTfmG4me4ZO8CVeRYnXnJnzLrbmcuJSOnu3lccnoBfhxjlguV24zj1BihJ
NQFHXshDl7SGaqAhq5TlIFX1uwrZtaOlyNuCd2zVe6e9PNgoFfAxnxSoJ1ZIw0BHfmCSwrLmZxE4
uu6HySG4BkZalcK6GRlDGectk7cM6FwSsi7EQFZuenXEpm7yjkhVlXrFkprb45hSVtl7QLcHotXq
1tIr3Qn/1wHuBYy2aKsKJrPKNpBTpv994t/zkFe24GWDrOC6sZEkrsKSuS4kBg3eiAKNP5sZ3RbQ
sG5zeTC/PvR6GMM7pCUYQwgnOoJu85IEuUeNFJlwWhjmtujsVRS/pyIQ4ooPn7ZL/6cHsIZkxMhC
8uDl4Q66OQ4IdTSJel9ABusN+b1qY5Hn9xPekCB3pj+yd638RB+NNsW3RbRuQtDDbOHpmrBj6VZN
gVE1fkHwz1FhM4c3dnf4GJFNSUu7IYIrGN37tQBKw/6w6o/YLDk5okzBjbGf8EflBRMe4FXhFb2P
/KWvjUU9wmiRTydKSKPnMPlgNv9zVQD9Ln85xyrMdKlB1SnqiNBQWwp8aUO6IcOlTXcxs/NrajPB
TjFOQ8uuB/YOA7OXa3iWjdqwrv8a+dPMPh88pDTLS88jNFEbYnmgEj0UHDhurPVD/FrOBz+QEGM8
DPT4PYawX0EME1YxDSVmWVwhYrOImc3JHFW2L/ue0CKsxSbU3WdCZsFa+dCsHe51JfZuiPJ4bHiH
yKwjVpx0VlICzQPZfHVmBgDMGQeAKVjiVQkb9uT9LELxlJfm5qpTXyK/bxi4TyAc3NH87fbkjuJa
a+mTqOS51o4+yMuQOfdIjj22cUAz7W/SYXrbCfMbutKMyiSvAa065SuHqKNhDlf5MbBMVXILYdgw
eZhAssU4KUlleF2GAiEu2a84tG0hwdc4lGZtVupDzck4xBG903nrz5KojJrJTf06ULNhi7Jw9/vy
fjd73oxJpRLCAo/P58QGQ17PXps7MMyuk2Ozu+vgEm4SBS1RjHtKWDs3i13rHvZpbGWIMnHxT+m1
ObAx/eFYl11YzUBaGnnklJ1jGWRJRT1B7Gw3HagcDRSTT1umdlw57n9Gho+YKD7xp/WJyFtC7s5/
glEa848EMJXstyPruG3eC2aFdYlEd76aNnsfcqqpsy0B4qiwkNXAliKWPDmTIrJFgUgM74zYg0Pk
L23TVVNnrppox+0jDxvi0zzU1sxVwLD+gqdhvRZdqPMznROP1s0PNAg7AsPsC9Ch1JZ5AHzQt/BH
C2Bl2Fl6c/iFYZqZqVcR9ugvQyx6wWo7GCiEIH68ZbFOS4bactBqEaL9NgbJesRP+3MpqKgUbSCb
xE2qiRmbTpMIVoCyKSU3P0qu8L2q/WnT6IhecQTNpw60FfdNVvnz2BV6sVDnbdjU6JxFLwyD4vDZ
ggiQvOorZteWyYy/YdciVTjiN+Ycbw43iOXIv89N8DPH/xTvhuZYlyFlYOo9hZcm2jwWu4UZH80F
YFMTpuVifVGuQQfClGywmGS5mO3NXVh8hcBCwOYDAVxHgrzuXqwir879XmB76D6J2UIlQ+ApyMLX
8Gvd6CFVEQkEFMADPilGd6CmPZg/o0h+72h0czgz9PsP1XAQdbXMOtkdEu533SZlN4I9Ov5K+Jh2
svQ6nLAye+3LAElDb1C+6PwqjC86276ESHAKky8sK4fCP7TUb4ppGMwaemKXMvTPgFOYh/u2zzhf
An7UjORu5n9kj3+Cv3yFc19ai34qhWGLD1d5mfR3nGzb2OcaJxFwKh+YiI3FQ6rALo1OdAE0z1rZ
6vyr0AzXP8jbp9WxB4zXqz1JBNxOIPaRlGsOPmW7BcWXDXbCMpMUZ/lxa5Ts/DBp2gnLferUnajP
LxQqUy36G4WyIFYmnswNAU/4vpSVYeWG5y0X+tKIooz+7WnyFTbmI3+si6ix0Ijh0SMjRChlVeY1
SZqp8gWEbPI64EZny+q9FYlX1FD+2umHuXDBHgDu6fdWnripFd3o5ix12woSrBUe68DBL2moFo+D
mv2FM9Gqgqo1flGuXYDESNG4c9t25SkVOpmBLL4nuW1Ng1XTmCWfSfTV0s5iAu610EEEAlsp0qRj
wkRA5G889WwjRnOtxAsv7Ib7mN/JC8dtoj36pPMi7yFboQv7IU/5VvhR5MC2IgzHQDSLTDlLNvoz
Plo54YkoRknFjBi4iW0tNoUc70lhlR528+zwa4AaV1URRVgmsqXONdKBS6FdULbQ5GkucHbSX1kr
twmCRRZQY4W5JjOzw2tR//yvZug+aYV+tnHrBgEdAkfG6yrD0Tz7Fa0Z12LEi12MuR24IQ7Ibsge
6M3WEvjSYo9DIuflN9JumXOyBygWwmlKbI8vqgWaRRjjCE17BBhB37anRJKyb3+xVsB/QkGBGVNe
4jZvLtKQXaUaD5dO8Irwd1NT94aDEv583jRK+oZ2YEufnVZiRj2MqZ8GunfoSVtAgjaHXUNgnQOM
J0qvfIdZvZWvFrN+Kr9NnLNOhh+LrjXt36VyJWom+tkksgc5p5KpbbS7u3U1Q7uiEmb40QtySA5s
xTZBPHESgPsDXmoFzl1+nxthoiyP17mRg8Rh6BJ83bb+cyaAGxmk0erFyiUp7GgRF2+t5HnMQdwE
WNlW/GhD09Gb/Jo+k0w2z+8LmExT7vkEccnl/hHZBM3aXqEbMYmow0OfUSmaswoFTI3es3QnUJzR
eFffhyBxQY5wfRWTQZbVTNdKbRfrYllFumJxb5gndNxCLbXqDka+GrP2Cg/2Ahr8AA3r3wD739tN
Lr0ymZBHtCqy5XaGpJITQLn6Ia9dwLT47lqrWirKtFDfailL2N1sQNH+WpMu8zHyas6ilaDbmMBt
ZZ0E9tgStr5AuN9gOIY1d+dopCSwyXp5HPgNecJYo/kWtAAT2eazRQ7NptcQ4buOgdbtW3de1rZs
arHwBumakMqr8QPk4TmsXDUFpqBvaBB0Sm7/JxSzvGU3oL2Vxr+TWjYzxje3jionbOrkxTP7F0EP
dEuNC/5eQhkpZabQQwpCd1lY0MzseKK8aosztuf2XtpMUDITnI8MhJ2viG3EfIy+aLIAYIVR6efT
YApMZ66QqIgQp8uKGCRley6OO82dgQu2d8OW//JV7wLkKl2DIE3RyQTXWkbRGIYCBxc4aRRW0jDg
pRCH6VlnBHI3yxSpL6IS2hmHSV37I+xjq5Nyh8phaeQZiNDfL0MvPDOPkoFqnRlAsGWxxFowFPb7
ePcREgf2u86dJz2g+95tqFju16gn1vmIjHJ1zwdSm5SnXDYb03jUNuHZWiJVDTDDFWkq92J5HBVH
Yh8Igb/Cmt04sm4DrZXIGFBXhIvb9qnP113xYb/hAcSMEgNDlT9HDzbxS8Sc9Jatqhq6kl99Y/ff
GtEePsvOwdbSS6m8k89YEm3D6uPYp6Gb/WiKx0+uxnegp8WNN9/i1BTcbMmSaTkLas33kL0a1uSD
Kmfd+Nd+JyKt+/2dH1+wwHMVRNS3hHDvCSBBC3LBo5rQvEpQRuJh19MH9Fq9bG0mNlxr5O3ivoG1
KebykMWBhvRCoXmapPSbm3ueMsp9dKNh1DUtNeV0XYrSR50w4P49jaBt7/zX8FsU9EHhsZzt9bFl
2KMtRihTfblR0367yD/qqdIN5bdkFoP5eT/XZvC8lk40fObktmGHzeZ4XkhJ+U8X4+24Szr/Cvyw
pq2cvgXCmDocB04WnOIAsOvJQJ/NeaYUKtDCyzPc3Enz8rOAUxtGCuRrAws2ZyzHKaWFED+RMq/A
EGgGUH0axl/kM7iuwfaHTHDfJaK2RqW1s3VFoV8236P4j4UuWuDfrz6Fks1HL7sLRtyhKNMumzpS
2v0gNO88iLdKfeq8/OTBU2HeJ9XFBxnCu55uuUCrmHatrUaswwVMEuKDopwFSVnLSNBQJvPT+gAF
Bkv44nw01sMwNJ+2lk+fz3J9Lj7DqFLb3o8qqRI1Z6A8RDeS/ccRZv3MOjVgBhebo6Q9gbOsbJMD
pGHlu6Zq3L5+A13JNeGR6DKvBobtT2uJy6iEQvqhvL8AJRQF9GDzJHHFPSeZDwlMAyGVNcJFwl8y
5TpHgLBErKfwoz2lIIl7ayHQ/h7crEOaogcB0eO+/RkhdGvkP1JYsH3BQVvqSDuoZSD9iXci0i2y
E5o2kbmXER3BWc0wNjp81ZCJqqC6yxe8u0TwS7ZDZ3OTYW5f/7G4YRP1UH5EpeJZTuCg9N3sUTQ/
SMiINm0SJNgqHUVaHcI6rULVs+JHxYI13MnFZE9umcDso/nxSUaAg80XUe8B4qADtR6uwfipSM1D
mOi/I+Up1upyde1cVOoMBXDjoRotdN5+m5JYi+FJlLIiBv75YekPXSEEeHQ6+JmxKPoL6/jjP4xt
c7tUVh3fAW91IunYqnYe7/G//3+BOlb1M0OtlnQvRYsctBvJ1nMlpNnV05Pnz8QYai1zHD9cnzFL
2dFnQxYuIEKEOFMMdItHG9+PzVP23qxLY+MhVkVAXG48KOb12wQgNfIub4DxcfDS4Ffkkk6+hOYZ
afyslIRLcnKn9APmIxgOOsuYkp0Wlrzn84g9nThqMZvnrhXW6d2eApQ5K5QDaqHItO+kqLSCTgA5
vircCHpAPKfCK0DhxvAbqkH/pBoEiudQ7+5FmUb1CVNBLL2HruND1Te2PHG+PKqG4ocfOrcNKlXi
wBGS+y7YPkhSDFBMB82ujxTbiAeAsjEBhkEnQQ607HuyLihUdYalro5v+k4rxjdIp5BpWvrnONSu
M8wimchyaYoVYcIkEyRltwNWq74hn2nRgxEmdh/aTt123B3818x6BlmA/BYwMQKLy7LihFSbtJy9
xCPyS3aU1PHbcoa3zCS7u3KOwWxxIIdp87zhGRyD8WJOhwZ3EZe7BzHoJO9EtY3jX2uNzzmu/osC
PoyfE8w4acjHbKcQWGjQJaGgUoqDCFxBHYHlESydBSJ/6MZ4IC9g1vX8SVMvuBlhpLmzeuaDx6YB
TwfARmkHpC6QS8S0Gi0tFmuDdXskZ2QZLI3aZegK5GAL3GS4HKYp9I0zvMwVGV1AMGuPn4HDIS31
ZVth7nX+57hQS6m4EPy+TTpG0b/2Mef1aC2wxG2uoF5UGQS2lTx7IdjD8pL8ep72UJPmYSdpiYpZ
3CEtIaAUD3nxtN6ufptJ4ubII3edliTxWvbhVREO3bi88Xl2kHSo+yPuLByqcGiJuIjcsgPOFxdq
NR7Cwq35Wqpm8OFka3zKQ+niqUG7VIQwwMU1IW2eM+4/DXn7lEt/DfTGbKDHQAsheRsld0K6Ak61
pCayG6wWI9/gk9uLPQmMegItnSMcUr/ouxnxLOzmGenmyxzxKeCGssaPFcW5lgoq+pTAow3qZXh8
MIPBtgb9aoiZXn6tlN0TMX43c9waKtScLoiPaFTlHKXgU+pYyyURmXmZinN2rgJSytE/3MSaqmBY
0BkRv3cZnPj2+S6moJ1Vapfis9Q2g3iChFuM3/+07afyVEaiBbaoIDx3anJBRr9d1p+EB9LGm7Hh
d1PuQ0xWM0GICn9UMDQQQBw64po08sK5Cb3K6nkMAM4syoF7gflIp3MV0tHusgYDo7VfsAypRqvG
Q1U4Qp2JoL4PuXO80Je/EtNwj0wD6x55qThgmd59nirLy0Anc0BB8fRIjWsr+1fK885QP5/1tVO8
+UaZYVoGk2f8Blam8N4REIcrscXwj1H5rra+1vyi85AU7N+S1iwX+Sig1L3qc5dmbt5lwEW0Ggxi
lc13EKTDMC0+Ee8pa0NVbo1gU+PGvRqdxi6t8S+4Q8cS9q/eLttW5W9+v+t9rDg9MwqpeZYoC34Y
egkdpHrSiJhPseXbjXcfkA5OGiWCy/msrRCndFuaM1K4Yqc3PwcIm5JvvX59aY74zYCQk73gDUik
+p2aCnO3LElqKgo++RzV0krzKwyxVfnccMsTP7T++qulXlApsRZFdZcPGcc38JuYCjAJkm8rEE9X
gzo072PqtnxjCwiYZs1ASDqIG83pGdezgZ/oerbGPkRosbjtYji+on4kF20QjfejBkhmFR9coVxR
NsR4YiwGN7Jr9xAOYG0WjA5B04cfOFjiIW12OH44fVbhrYk5TjiBhDRsf/fwKKT1S46KdP9RisD7
9HdUthhdJPJToNiNE9YjEDSXKexDWAAywa4u96bOzUDIGn1dyx/t4N9SdNbrdQlvG1/XjqcLWOQF
VEg/COezbiHlUcZPckGpYW1QvCr1OycN4+BkTQf4UEcIZFvCcQkXKmhU/vSR/cME3KawNzuKUslh
LJILQE4alEfQshR1CRkc1mLo5AKGFsBNyhY/tSCl6uGJ1fmmkFkFvSZdeIb5cHyVaUb9ZIslYZKv
J13Sxo61UTZRFCGgV6O6CMDrYfLaOyeKMiybyVSniOmjQkKURyBT11FIloWLpAO/jBHs4ct/sPQS
ZQBA7qDArzCZNtliNUMC6hXw3heGYokiwijgm0A7JNfWILgy2c8byfxKCYmdiE+PabODc592YCgm
q75VxlLrEFyndBtogcdNoK/UEZ7sMspdNCaqSuNqRG7rDcaDl0nIJ5/YqQm8nkXLxYGgXCawCgVR
7Im17y+/CeZ3hdWlt7O+3bh0bjZZTXyvm49ObKnHceMNLVnHtlDQL6hP/j8X8Dp0cyDLFYMFykb4
6mGO0C7/5r9LQKsG846aOimv5ADXsOlnCIYDVoFRQYH5cInV417A/PdCZVyJif4ydeRrPVbyCEG6
+wb8Df+W8boN8gq99lcQO1gzXIENSaWmGZ0D6Zau1otWtGd8G52A8oyjRAwCmi0os/6qSfTUeHFY
38H2Emvv2PBqnUza5Dv00rXlgEOyIpGxL3g9Mjij4dv6CSNdoCm4ijzpdG3E/igAsG4WUPp8oloP
9u5WvZzHHVeBbHRShoywsez6O7bS3RuDzlHLTChZrsZVzDOPMSFxe+kCPI9SOsxDg/SykZeAQ/bB
tXZGD67gjN27/sdf+hkj4TMgWh+4v1NQQmQmzwXDhpqJI6mhh5ucP6igh5rn4STVs7Fs5eFZ91kW
5nX+X6UB4bfpQkhFSXkZdSNb18CAobAy0mw+WTQQ2FhlQnDDbmM2o5LdP6kfjJOwQX4eQx0KyGHA
VDg2iizmOOwoJgED4QMqaYQ2msDtLU6SHeG25JHq/g6BvIEc/pcVzkSnviD/jnlj+BPGSorluDFX
Xi0XvgHt9HSnUgXTMVT1ZonFbPL6U73X9Xy9idcQ7J/9eBXAszKMWnAyMPwgHhszs5atSKg00JPQ
mptQo0vcL/bSJ8WbMiBz5PqYHy1r0/jsWC1b8Kt9DbV/L3RZ4rwuFFRuCYPgXuv6SB+95YAfa8cv
1eP77PxA4BNaY0udxj3MK3n3MndNlDzcYuoGdBoZp83uSZS1rBEoqzOZzPDRTResBYhUp6l2wSnS
b8/NR/7Sf9eCHrNqOWWjAmv8NG0snnYr9wG5+xzo8dh7Ba8C/8c0jflXjlG1PSJ/N4RiptNX9L4V
G2atkxza5APmDnxJjJ3BrP7rsE8BV3UzFoiXU+AjgDHgwY7t6Oa2MYfrLD2s7tqzWRSncbHAhD84
be1GTX3J3Tsw23FheIZ7LTu20F+8kd2pjYERdrYAMs8iYD0pYPP/oULfkTjV7dTLFBGiCtTxAGz0
iGQ3yO629JxN8pda/xGH7eC4TD/+21Sbj/JfcTnVpUJt7AHRiaPvTeFWcg8+hICjOwj52RwlUHr0
ToKAxeoaMhZ2SwSRCDuuwqtku6wyGD8n+OuxOc8ukvU6s+25HX/nZ9/UVSkkQs68qs43yd55lchB
xPyh/qmW1s6Q7b51hoFXozU1pqz5aLQ1in5OPw7n+chZICnvS5dnymrOeIJhzEX+ZjJLo60aoEZw
2rVGu7BBerwZ0mQdUQLeZCwEeD+SpNSzW+msQ5i9InzNC/0gsZo7fy77SgiaydSWLPk4tfNfOK3q
plnQZT5mNmjfuEqVX4P8DHEtzXhld9EKIevZM4/odU0uO8GmJEEaNRDwnpvc9EYsHWR0dHgxYzCs
+Db0ITg9vP956MDpnrMqDGTTaGd15HIQ1RKa6EJBhpBHPjKbyNXnQ3wl/VwObhBs8pInzZyvlQWS
cpo/xF4rclhnSqcY68f76OUG+V+8L1Uw/t8elxInxF0l5Uq2lsk1EO/R5ygtMfmeDfRp/PYC+Rm/
vaXKUWO0g66yeR2K8FzP+nQtv5xDRoJvcSExczgM55vut3Dka/ElSwBoR3CkeqxT3p8Zd8dghRkJ
1iGVZhSJbY2D+jN4iNMSND7LZ0trVc7j0Bi1xN5MnfJbzQBRzOfRzTV5OYgLi7GPHs/AWmH62C1S
v060r6szZoj1GaXV2OdGxxNXiPDxaiBvaHW0jEclVPNLhylSNOnHbOAGcWsX/nT2kkMoPUMCxc2q
w/CEBLQWqVLrvFhsXWnV/N/9V9AyOkdpS0O/DSjOgYzPxQ5O/Lrot996meazS4o882v0ySHDch+E
jZXYRZWmEy+0qsHk4K5lV/M4fJKuo8oFrYmXD5CvHBNG6TK/Yg4oCLQf+JfzeRsIU6cL2jCE6L5F
y95Xuml4kJ48ZtJtOoVRI/lBX5qXL6sFbb2AW5b0Sad7V+Tq0n69MRwLHaHHRlT+F7CJSCuYk/PK
055a9PTQtsld0zty4tBbqTFKrhu7l6xGkXzIfv5Qcky/mPs7x8zx1sNCV0614n/ir1TAgfVgluak
nKBxzrA6Dfb2Pl34XZ1k/uxaPf0cwKNsyvVNUGT7ZQ+CYFYSszf5SkBtqyRcWucK0hPiWrJzWPb9
EpLJewYtqALpDXIXCYIE/To4BTAy97qXT7fl1Qzb0oOnIjuGTM5C6ui3cShOp6Js5U/wUUaLTmXU
ueLcAyN5NEWP9P8E2jmM9VHc3+fosrvW+NzOQIgdmkQVe+SnHRcBxRleEtJhEbthuxfw+2xSFVc8
kFtEDu5fxtKG8jlSprFxfLPRRgwLjlKiekqNYOTub49lzpYpJnVKhFNgNJs0nHh6aaWyuN1P/Wdg
xmoeWmWuerE8AY/SAWXmkO4uPcScZe3Rm0Xq/bCLo5TatbU5jkCPtVc7862IuBnO+gXiJv4Xy8wI
1jsmQ54kEO4AQ/+JEIaR4jgwbeKZggG83mjQG9Z5ZMqszXhcQ7fe1CS8yDnLMSsYwWAN4tJjqUnM
wl3XYKQic4Zq6yPZ8tjGA4/P62voMuvYvf84q7jhqGvpS8RDfGY5md/ZU82nPkWSQ3dVD4VJouze
YVX4LFVyn/ttTK5lBpH6cHNLbmw907vxHuHQ6J+Ks15tMGpsWmjKdbuc/Y4WNwElF+DHqp0YprgS
JP6gQKq1AV3zUjGP+z3ga/blVqwsC0nUFD0QcHdzUsjbSC7eL1p+UeXs4sEDYl/Isij6ElqRDjgz
8zlYH7gzoeRsWKftxADTB6GnMKF9GeD1qoCKwDH3I8LQJ6GpkSDypEUVXpiPXFu5mFGW7yB3lota
Q+cdZZ2L0DfgNjrxilhSDUf3Xe7lRtq9cMEEVUh8ExQBT4mw33od6CBTaNNiARW2kmHpnuAXpDBC
oqFlEk+hSmUzIP9J770wsZYc5k08RUkEay1kDeAfpja39jdcVNJEIxX4SMOuYlW/0DZjoeiLdq5q
Zwe/kl+VGCmLfy1ihFZF3R131k1K7JZ+Y3B3OEfwY3udvdakYVrp/mAThtRrJl131mZvIgSUEioU
3qAlgAyfAe8iP9Gl/ZlPNS+J+bCtcayUVSBZN3Ajo318McTSFXnjy4ujic/LJp9eZictM0WHGL98
WvWiGTddmGaze81x1NVrBB17vBMB3yjsPrHffswEvZS+YzyrVrjYIQP2FMqouXgcQ8fFGrnnmh4t
U+LJ3gi1QD20KWERI2EQGjx3XfBTUYB1+ZDXW5cwQ1zlQUmIroPFLuzIGHJ7NiZSE4c5onAAzO+m
Ec2M+wyC5lFKW1/FUIR9WiG9AKq1OxgICCrVe8b+r/KEu7eHQDGJN6b5nY/d29/TmIfhlVN80zVf
r3Kd/RX0owTLJtrKOTewe6TgXQi5OGSq/z+v4pfamdB+d7wOT6n5JKy4DjZuEBgs8W8amGQ+mgfn
9AMTe4W4n7miktxKRIGq+vXjWhbjTrhAUwuOk0l+NArhC3cxvzlMPGy1sVBER3egn3Jwsn5G29dD
RpP6J65WkksHbPgkiJbn72qcGCC/MvBMqcrVJ3/Beq/EtnF1v8XALLkwG+XRRmHbvw2fypeS2i9W
eYQu1n+lJrd6jxD9QuiyJHriKr7t2DdCX2v/yP97s7mRStdS+9S7UT67JkqhoR8JPu/VCa7OiQhQ
ssNfCw8kcFbCjX6HKGWzr2tqXmbFaAMc4k/Ree/yQkFx3jHKeJau6cAg5HKyCJBMOkxFaGkFg4OX
EtsWXlAjzeqPb/+slrQad+f7M9pbUuubxAwxfoH8x97wo+S+ZzmJXkiN8hQ5fL7uLtO4EjQyaSTI
dhHgvx3uOYdKj9lDMFuHgdvwmC6/zFF8t9DGiFOnBIBKxSOtqRUGp1eHd5rxjPxRzQFw/9Ynh+lJ
mYVxWhPhKCPeoah1co6QCsNUh1zSUncrtBfh7bg7E5OiudRD6GwEQ34NWf7yDMQ5jATJ2HfEi8eJ
uhn1ljfEr7yceZ0OXGug4NrZ53SyfmziZ/TYGVoPos7N3AQg9Nn/pP42l8391CUTeN8SiE5is6er
AQycDVeps7UITAMmxCIacua5kefoaadQJB/5qyAv/LqyZS5zhlQ6NkpH44ZBtFZWzkE8cUxvkHyh
9UI/bVBQZwa+8Qi5MN0RWOoWkWpltualeLOZbP04BdeVC2VX9K38kVP59qCCK7EfMxMEzhQwOPy5
hNlxyCTa5BAQumlTX6PiJ5wk7RkzPUMXVebMmhDpGWuU74DGhRxnw+n+OwvAwve9Y5rbIRpKegIW
+PIY1/75dm00TFWmHC2uSArVNdBIwaQQ88iMeVuXz5Tu8XL/Nl7mbSkRNpS7EF+q2hW08Gj3PtcU
8t1qRgH16R8Jsbxbc1xWAZsB0nf35X3/Uzt44HYDXMV/NZVLXgljTBYp75QzqbM1OM8wlf6H0Lqh
9G0TtArqadcJbnyTM6BMQQ2wdZgQ4ku0igJ3NmPAZZ+LI9NVTedYPDF0MW4v2qx7Nd7WqXizLhd5
0bExlq+eOSoQufkDGHZ67C4RZu93nyNmhu83yx+JlzOfJli134dvP15+5kOyl3gUmyMvneicnlnu
Hi9X/ghprchscxWl1mqg3nZEj63ZdZXs6vB62LutWj1Ajad7TfrjZFgGWCcJ/6w/HCMF4RrAM2lY
E/VmpHO16zOt8mJgbjPIfl1aE6XSRGTwHkm4kmGRd6BhcZKCXybVuvlSCcCj2vDH4/+LsF8uWox4
8d99l++B+bZ/XWne4SYfUFM0OqNW8YIbYtMXxVYwJQRW3aVEvxpuErXbYQm0F3EyvLq1f88Wo9tC
yXr2rDWxel9K8cN+QSK5CL7iZptG1Q5OjUwVc1HXsesn90kh1KxRdeFGogSexM1dfltPlGatI+hE
ZAJe/4VNWxyLzo78ZjXNtZ63xo0Nt8kRTP1/VcB7lYGodcTSFvgWqwU+5GPZGX5ikbMwf8frKMXI
zBlxmmimetWLUkEA3iQNk1ypyMsrfqutVAx0kecxbSYVr3C3ZYTE0Zr9W6KoGtHluytCzWvcP3mJ
ObGx9jjDQJlM35xb7p5uFHBjg0T32eiQTgTYliG2oyB/7v1TnTmQbMzoM/Fr1nMf3bhNlIcFZYDJ
RoAUD+5pXkzEtqsgK2aMA3X5xT8u3KxNr2S+DMbg4ihSCItsUTGmo/6iN1ekyn1C76YIWURwKMcH
nedNWdbFAieAC8iwmUkEeCdTt2C5kyniUAl0rZNlV7U3nYXafDGvYhNsd9I38KEqP9Rzfefbl/ak
CNBwYyVh8ea+CLRUN+1lq9uhHc3VYsv4arBy+uPnQNDnCUQc/ZnO2jUwqw8DrfoT5PineNp2UB9U
e/H9cIFmdgtcRW9my36411nyn2sfLwr684jcfpdb5P6hpO5AXn1ml0KtINH6wgkb2XY2oGFGqOKU
sFynwGigEubMDuX9M04jHW7tMQwItm+TMhoJzHsR124RoU6Nj6h49xP9quS3DTIwpFngFEFdy48K
QCMDWrBwiCLCp7o3xYEnfgEeTLVcmKxvpXVLKhNpepbndI1Ig3PG2jVfA0pXNV6As+0fQhYOr02Y
iBRIWs55f3n2ATARlKsKezlmWfNf2TOvUFjG2SRXbn8Bt/7jnYx9WoXpEL8E4/QADUZKy9RvJcqi
V12fZxfFHGw7M3bsb6bWNe1NuyzEyR2XfhN8rZgfH2AaB6gtWUVYYsT16tIY6SATtYwcH/uBMw/e
KBJMLpmXzgEO9AHO2TRx30gacZ46Wg5DA+mhXbGP3NxWGmZdFewQlCjB0suZ3LkqqMnR0UiiXXEZ
Qun6zkTAFPrMAlk/xgoUj7v8CGIAxztKVqisjKqREjL2GKj9SeUmZzrFO0WYBhbPIwgtEBbG8Jg+
PGzAll7pAIaUhDy4A4WZnKrptwEtt+2tXobzGnYwGpgz00ATBvl056P2H3rpwwlBSNl+SsTXgijf
FTAyI0z8LHnnMcMJJHOSpHyqt+6R2WlkftEd5Oun8jUEbm3cWEafH0DOCG5RRFqfdE0gqi9QwdLS
kqS8D4NIcXr0JaJ5/bNXsx2SR7Pw5nEVv2oR22qvdj4xZ0qmca0NGk2OTkshWyrce3gOmw4aawJb
H4B4R6ZQa9Mki2Lg/yp0kh8CNfLdNfW/5ClspRj/0jGiQg/7BePCHgRor1BidMzndFw9GW/ey+CD
Hp+S0Xvpi8bNhA2CLfkZBjOj8ixMsBD1LwAO4G+CB97J9czwH59q3ZU3wFdU/Jo3m1PTgjoRhYha
KE6rzW58hgrq9vo+00NHXR9NCi6GMJkI6t0q8OxF+YANxrxezir0W0xRvjJ8jqhIUNWJe92NELIi
yntfPy5Mqrdpqj5dUhpdGpEzLkIa0OyZvNjlSqAw+P1hCigstu1M+/xbpTc7ag1d9TH2nUIVhJXb
pIZgjAcpIYufJ/bZ+MhHbdDCtp/MrKxe/GuTnit7AQHjWcyYBWxwxVn9ls2idFKXcWDZRq1ZVp7E
Xu1p59T3QutHevTxJ1dZY7QLpuUdiPP/Y1cogn/CqLiTaHB/X9rNjwLGvU3G8nnudInnJmoBg7jl
B4L5J83+9gB3r2YxBlSSV99At+MBEMIcv41BfQZZlk+cc2HjQpupjZ7XJUPopTAAHJEPdDa2z+T+
/DkK2ee8dy4gNLgshZQq4sEQ02qBDumvtcyikOLGoBRjt17Uj2Z20xgRfQ1zCgbWyOqlxD5eO5Ov
NLUhy/7aPKA9GuZ4TleBRPd/1BmF6eRWn8nMz4wab3ybDV02J9uCuldU+474SZUeSUbF6YA55gI4
bSo+AiKwRA1SZKutFMY6t02xmLQ0GvBRxz/mUbkolK2nzRh04utw/ZDv0koBPXFOH2w2FkdnZ22G
Q7N16TFTN1BODCwvxdS3IV8Z8fOMDEd+HhP23P7SV2XYTlps+I6GNvNc58z40CNqfTP9GJjyJlCi
JFVG5WRo6XLa5gGtVMCnSp4NC6ych/EeHzkHj6Fgs/NLUFC4qKQbrnTC9Ce1UlnyS/aivzxr6kzB
56ZHckGT0Wb2HvfUfz3PDPp7CcHBelUn1jDjiIfptNymJrfLSrL6WbkNbgCvBrBQ0S6XBI4MUq+F
yOVuNZdqxq3G1WkJYGsT360td2C4l3bl9LglISqKpGW9ZA8Q0S91QhkDpVUmdGy4AzDKrj4Lo0Nz
+AAT1rlKX+MCtTIPcbw1ioIc/jJlaN9EkCne3aeNTRemI7QER+tLiIJLMUhD92JreFrXmjUQMj/2
AzIWE4bbJ94dT2rH4kM4lK6PNetcGq83ORPEjunI0kHuxD+dAZiX00UWSavvNipSJYJ6p9XSWvA5
SIbPVkuhwMmCiaM6Tzoym63zHaHmi6++Me93IpHJPnEdKjgFFAvsuieHWK6JEE2FhLLaIVuz/ifm
iVbgY1cjHpRTnZ2BxvxwE+lYKQuAkN5f3eTeE6pnIx+U72GxPOcBlvNXZ0j0HZyrE8QD8PM9MGRj
dFf/f52I6uhkvRDVncAz/ny2aZNK/JFhchHcq72u0bjBuWpwnQvfUEJKmdWGfTNo5szPkCU1w0Dy
OMCBDEVoiWgxMZAgls/PC+ob+mjBubMxLTU6zR4cq2rZbwWr+GH7ysY2x+TVzAaZkPQz6c7rZnTV
ZgaXPdXxSTDHGcmL5bGiPjaUOZAU0aar/Phin9HjfoeirdhWApp99o9K8te1s0D8cvVJriJy19Pu
SXtbAkVECezbT3QNWsxrGJXH3DHp+/F3v8dSNPmBItY/mDDNdi8cxcrxiAp6nOP2Okn77J0LV/do
7F5ivdr2RYrdzrubqaQ4+yw6isS9CCkL8J4n3aM6s9P39tZSw/iwm/GpVIqUbjlnXN/zX+G0vqlu
4626Ck+pieho+oYg+6OWpLcsXIJCXhwp2tQ7OHUbv/jkj3lRm1G/7rNRh6x0nlnTH9IuNpGyeurv
dRqH61qDlpYiIpj3vubLwwiZI0ZHS8D551acSljm20mYSebz/B/X/pkppAjvSZfMj4YtVfwdWq9+
zC8I1sX4tTXY7dhJ8m0FlNXJ2A7aUTKavNSL9HugIsBWudWLdWdE6ml1I6wd1gjTffBp0/eO5on8
cHMPKSd+W8pjJ8r7FpOcA7NgE71WCryaAENaGFtYWufJv0JHui91KYyr2O/cjPP54bmDvqJxOCse
JeXHALjRz4+PoHoMlVtARHgHCNrxhA8hJ0hKvfAm0HDPQ8WTfFUqmG/ysJWivukWvAeXzJ9PgO9D
CXXyZ7MntMv4uCjHrUcfOONu8TBWXeQmzC+x2Ab00mQzKtsemERX41QisLYva7QS/wSR3REBOV9z
W0uZd7rrw8IFHEtJBZSud2Y9PlvnDbe03PF1G6XwJNJVZ/Ime2RX+fwpI9vhrXsHKUV9BjKcbAaV
KXwpXMOse1rxr88r0OQvIL/DQcN3ZXQRQMe2xMslYamGicM2XZgkR1XjDULEFBYy1yzo5OwPEjdM
vbqfmB925Gc5QDoULoP75i52tFgy6aNY4/8TP6pr7wg/jpWiA+HyzFu3zl6fWG7hh4vvzgk88wV+
TN3LRsmzAnsHfLbygjDUWYFZyP5qHvLiRn5DIZiwR0K6XqTC3ICMTngsqWCCG+woc9hU3Wq+SLdb
bgMFJCpI/DNuRqqFrpqhiPLg7Y/F7IUoNnrD3kdZSi1Eraz7WRH7aYDVjweT9Jssbp328UnlPgyy
UPK5hWHlTPujFJjox/j8J0JsalPifXFd7oLQEnnZFcB0NcZWPwH6F+bPudnbbnMHFoqCSjV//k9Z
xqx5ab6hFtxvgDdIQ5SVGpkDRA8fVaP4jG5LbENABgA8tQnvzgOY46gjb5qWlvkzGJaCCU9nF9z+
gGUdcC1mHmfxkGCYMpdbpx/pyqQXDhllGAFTLyOWrKEde1y8CSvBkxiLr6hi0rgLKq3loiKpNlsi
jQXiUpdA4BhbnKZk6IeDpFmVo3P539AhYA8tRgWkc4Uv0VfHMaSOMtnB7tIL/sSVwsF16ujlCIIb
dXzE6lDx5m5XK63oibEIYYzdEfHIxjtGWwBMK83QXaW1alpEYh71v4gaQGAqrGQluHX1Bcb3RV09
jlXDaGYNjfBKezl/+TvuhDd9nrFNS60aq4rhB85OOEJ0rra6ZDMcTBHiqhaBMRUGvJbf/K5Xbbmi
kuw/h0AN9Qjfi6Rr3HlGSQShSsZtVDCyW8G801Wz2ld/iOTXzP2rDOpx+kyvN+sV1JTHBypU+Eia
2xpz6juMdKaZTYAtXqpLvFNWMaK5PH6LiPDeCVT/E1noTBxcy6K331R1kYOxnRQHwmbbiCoTs3ej
Tts44qvrTDnp2/earUVqzpXhbDaS6S57mqRJkF0S4EayHaHJp2wfYFjf7J2KvmEolqbKguouUvaQ
k+NDoTh1Y5RojOiQGzMdeM/9/6kdjAlgI2/DmAJfVEZQOjlXdMO6ftMZyBXSPWb09KXIJp/wetyY
De4phfSjGlhBGEsYLkYycYf+XB5afZXaWTeOzLF6D5qL5KkE5GU9FDDROWLTt6lu1A5Vv2DtXl9y
2XDvWuDbEbpbn/wHi6GhVByn2IZc04aEBlVZ3ayMcb1ok+/Z9NmjbNyRwpsCrffxrvMS57SAsoiN
PjtmCbAFoS0NwuNvgxWhDcfWDAGyL/zdRFXMKG24OaO8QbKa2nW/pPq0QWHGg32sY+BdFyE+pULY
reSb4bJeLBYFUVupowzJtigqz8vNtmgO6v4Y9xekyMbLSohlMYk2uTHQ2mvlNWePaq4UX5FH4tGJ
EfjRpfy5BlJip7X/olPXc0PfJ1rkjWAPYcflo/IlMH46XpOi6Mnl49dy5hUrDs1QBqtvQATL2y4w
wL8O0/mi0Amg0jqgRdnGu5CdnLi9nK7UBQZ7ky7pgr0Aba5W9XKf/BxZ9eXr3T2yzs9ntdkzEKux
PP+yX5iRohN8/Q/lT0V0o6waC7VsqexDUe0+m6YO+O8hA/FmL2ZAJKu6BaQrWTvEXHrUYox80Lt0
9ZXMcr4RwEWsSlNYWPts0fhuaF7RYpxGbWdYby150/Z3R2JJc9nvT98qONPujQcnPrDEbM+Ln64C
iOnmcDahIA4i4kzUoeTO26c4oCHZTLH14cADsi2uXFnWXHee6dYh86gQ8Wpj8sgH++vD62GOd1Sy
3o3+XGb4zCWB9K6YYHfWnVUf+74xGRuR5/VevEOCyYUGM3V71jppI3AMYFsOnQ8ytCYHnWrom6My
AMV+gGNXuJx3hDvrR9AgtkxwiCOnXaXddVKdHV/WQK/ukl4Jzc7Fo40qff8z/vAtBZxkyD8x0CDi
ZUV+/AIA7NDxxc9o0xe0PHjvMGcK+LxjNdL+5ih4dbFxGRYFbXkoxh2mY46UiH1FWlGaSpUjZgn5
cfzJJjnwbSJap5HqZvZbnpT1ph4FKhlnMAqSencPR4xG5BSQLme/POibwepq6p96z5Cs8REP/wvc
8sYmRAYUGas5CkRSxOc99tD3UrRRrUrNZylG27Coy9S26n6wULbzbschbMWcguXKGjeHV0gL/ilL
yJQ/CYtbkFYWXxLYaNHzse9mO3RNE5Ii+kPC6QjBKkSVyCinqMH1VF637uZw/VSpjcE5LCluYlIW
Fm1k67SY/Hmjb2ftl14UIBTsWOkW/o7nu9HQWEoN0+vSj2qVbKWsrak40OTSzkgVKgZmorxyDWb8
kYH7rv53HnwjtR5uAph9H+j9iTnBHy+pepEjhKXgJN4KGCHsly1yBxcWBj2PZO/4nlEfqmTmrbtP
cKmDPqrn/SwICpa46Z7TyPQGArLg7eMPs+gXUx0ZLwJf8ID380CYuBJw41FqsBUfiWD6kCicO40c
uyUPT12489Jtpqa/vzncCb9kX7lIHCQ+US6WwYFeNl3+laD83fnSqpQ8nYE4iJzMYOH2tztqbW7q
VwaqPWRKo3bkpvaS3tifNlfaDQz6FQNwkRUq5qWSRsLPVtfx3Le9cYt71U+hvACvpl9XRzHuQU4X
69tuueOEB6+WulV6ksM0rr9Zvxm0kylubd4x8In/pf1UgH/S9s4E5q+ziQZphFJ2M+ilsEatUmrL
D7PqvsWTotbTnolbQHbQSNScylP1/94h9nDpm/LwLysv/gz2uH73Zbb3+zo6pOOj6vS2rB4pCEMC
QwCKw00ZfWHst0o1Um4UAUVPLPD7UwRgfUjOjMqbrTmjbMeJsdXZujQeprgZ6T68y3nWm5QdhKWw
QbACC4Ba1qqDqOCqL/N0lXKA/bHZwcOpqQq1KSvmgSIgxPy6AeDAsiPN86JXyMwF2un1GjO9iiMb
eLv4dVKjJgmgNdIzAVVmgPyHIhGq4z5Enm+lBB5NC9U7w/uC2H8hzVkoYva5VmnTeW2fsCQpU/LN
+hHBq3EbfYM4Vowy5jvOdjseb8wunatCdciyvL+tqMi+xJexBAfnHdIu1B+gbj+4d3HEAcy2MDSZ
XKsjnHrgncU1luQHSnlj+wfucMh5b7eRW76rMECBvfMxGjihT59PU2amT3RbUKpOC58yvCnNZsrr
SiZpoI4TeykPgnjgcf7h9WV9MY0BHfS62Nw+1rzFfpUn1EpslDsKbOc5aonCWNrzHg7+xSQmdmSb
wRvExvfjnRMKA+9OTTe0TJh+cEkbPf/W6AP6xq3/H4adpQJcqC6Ej+xVJRotzBbuFmomIgIq9lM5
toBCotWcZo/QS0hYXtoVcfQY3wooMyRpjdlI11Qbxb8pPaAs+4ru/lcXNByZ/OTCynxoZULnD14R
JRBfwapKVfSbUYZlwobP833jy2LsHJ5gLKN5vFZRiGABCt4LImI/3utV2eA4bxUo5gJK4GTDISZ9
lQL2T1z2rSJw0DlRn+OfAYIjqbQ0s+Tq3hxbp/a9SxZgg5YuFWCiweSJRqRzSnE3eMNBH656CIPw
2+F42NzkOJ9VOddUoJtmYof4IPCr1iDBfu0yHxkGcZ9VfqZTvpqJf9TJ7f5fJQ0SkQgzh38htQh0
pXG5+ShvPxsbMcwcLr807J1O8sf9bgH+Nojckrc2UUX9lOtC4HYYPq4VQYPpb37y6/+UBCtdGvAW
fTTc5vU1X8pfdlLt42Is94nr/xhHeO5AFqj1QPsp7liWnK8m92fIu8WHvTTV+6Tw68PIk8Xc3js0
D3MVzYdSD6Nr0GKk2osqOlgCktX0xyhXYKwt0lPaIJ+PX1C5XzweXyZnCHpdlZQtsMGfzp0e8oZZ
2DiVacdEtW6cfmxO2LMopmgSuO23AfohAjBZcBL0+CROwE98RlKh/hm96eQ/xlLlPM7/cWdj31yi
WpHXh+bUlvo8ltom1AEq3M+h5aNzORJQnk9AuY/9g/kfYGJAI0mboeZnPcc/3eFG5P4rpSY6BRSJ
pwOZ3HGpE/t9QDVArDIcXYal/XjKHvcjnvJhHy7CTYEuihZgoIWxQnvQQ6/cDGQe87Gnk3BnvBOA
JiibJ2vjXV6kwfCcRIq1LIRCwEQwraVxglY+LuQIRdh1pWy9eGjV76f8Ff5fzQSBrcjySxGrTPXI
pmeVyC5VK5++8pkmKM2VW7g4AEA4Jac48slTOU85nt3yKth0YAV8+bG4oDEOkywhN+6BqXCyFpiG
a9l2fJd1GgEe6OMqqThZDikj/ezCtqb9gPRN27/LEqRTmjHLej8hft50EC+RuMrUT0cQK4qGyqM6
asMaxVE69aGvlKYNwhMlfBcMdsux9HUdAQZsAfD9Zdj3e+Yt58t1EY4ll5eMIfBl73QAjXpaEQLB
xoNsPhMlLNZH9HoX1LM31lk6+S86ZBA/8Y7Pz+EOFALwtB8SiaPyGJEf1f4jq1w2vqqxlW4fC9Ui
4fUOTkJKW1jGRuNiiGXxcKy6rBg5Uw8KAMhdzYYEySSTOXa1neFcRe+DUflFUzpuorW+5gq9Z/us
XySJuUlOSDaw4FHyfm+a4djQ3AD860acZE7i4NaYWwmmrPjCmbQtE8Swt3HGSLocH8qE94qPW6H7
2etXe08wB7AaaM9pBHIYc1m5fYKPUm/J7OAcBErdlwr/rZku8n4emjssRQA0E5m6TK1Jufcqguoc
d6bz5azAT/uTVQpNoQVfmRyV4zXPSgc6M/s4WZJbn4EEoKasvSM4wJMCJEuw9G2qYeGjW5xWTNWE
A9QQzwPZqG6k10Ps7CkIhj8nc+J3Xe56LnZFwikrDW13vLQNXZht7STpzOxmMJ1pVc1sLIrzowUf
WmyLJUENgp5bNhvwwvL/gFoscMLC3pNFpCghJiDfPVLWhywLOa34mrpXz3po4Pj0XTX7nw/QiEMP
/bouLN1T6VDyPaIc4+UcN8vxQZEhl6r/weWaptgej8hZtz+UVW5o6lGz2EiDjX3eACjco6vupCCs
ew5+KXDRfk4HHZ2sEJXgyBh9Tjv+wNoUd+4iB5lu6aaVVF26LBcF7C7j+pDvX6/WZhSW+sNVRsNF
LQ4AY6KZzFZNucibNFsvO+VCdU1qgu7z6R1tfeGbpujHv3zR77vmbGbBq34b/jPbti15fluf47bv
Um6rwLimVoiI+ni1XlwUaCy0kBhbnG9I1IPiREN9RLi0uhY1lq1SY7UMiTtBFE6EXPnR77Mow8ie
Z2GU4sjKnYynR5G0TOTC5DoAXkRC/qvKq+E5CuDLtWLYC3EziE3q3N+Pep6IgPXciL8hXCPOhbsI
omraIZZkMiLkhj/YLU8yo+1YPf78RCuAIgQtgCSxzi5FIN9pAcuKI5xO4mJmY86f/kppVMdPSfLx
CXYP1bMRsp9+52A9dd4nI2zfE2NT5kpU7B9tc+RmDWSi9S8mEQm3WPbJOxFfVCkkhg8QK2hitBTg
ENdEpTgzieQh3zxUoDGRf7GPm//IKcoo74Zr5qGi78OI2f1FRwHuBTQJEttv1wwtg/CCup6clA3c
xvXYkrvmUrqjq1aQ+xjB2QIhgqr4k2yamqlroDLAFkGfpmkfx3tKyEKV7NumQJo99dQyvHBX6y/n
znIrLKxnOxX93fRryo127fr5E4ASSY70qm1nN/I22X7os9gPYMfe/pmcWT7YY7zjdjxEHBsnEwW5
7xENWDgUTCP5DAjBeBfLcXEL3uukRqnfa3GL415/PG2w51UHL7dEuBaFLSZQuRkv9rFJx9pKjP4d
xLVcMllmn/a6JdPk6qCK/ADdhcH5g3+M0cH5+DvQ+AU1QDUL5y+ku6nYVJ4DBpk8KQYQSnO3orMK
8z9RDzO5CH++tqqN9S9ODkDaG9Ab9z+MTf5CHRnJq5VhRI8VVtGCU7pi3fZ6KaaDBbsmky2KxFT+
yjeDc2Q6AMpDduEsxsoOx4jhODMa082OjQHgUe0PuNSIpIUN+nr7EiJcwip9Bpj32ZYVt/J5Gg5i
vr4ExN88EsCKVeXbylStp2Mx2kx68X8o8e0KSM2xiR1bbC0fCyZZ4Gue82c6NKLLt93ax2yspgjP
mT2EsD7xxgUDPmNpYQoROlidF8VlDmYnF1Zou2AWyePwePFj1Fm0+KozWGsfYjgr6M5lc7WgwX2f
up4gPBhyGWFW/wrb56ln1UlY9bl+E58zzEArHwadImq6x04pjbEjdP+RLE0BhgxUYkmNx6Ffb9TN
xWxE+jZRki5kqKzckowrKeTl42FvzDwjC0QqTREqHwXjWYD2UKaF0B47fH4Ik3O6ZzO3sDNYBfO5
eZJwWFXsVgFyAqdaa3+rYTvLLDQ4PehwsRaMTQhV7kkkI3AxAbdCFSyQ7pmbt0DjVQtmg4mrWzQY
ccdE5eYIzCKo+tEr/Aa0NnWNYh2IYflACyS9hlW8zqWz9ffni2F0WdLeNy6Xqsff8schXrJgviLL
85LavKISQZbsSk7O8mJMjb4N7/XhNBcGcBiVN1CyZJDRr5Qn6QWGYLva4t2abDtE6XRuHCzaoB0O
1CGo4L8PeD6P722LStkoCWSon1nTgsjzOpQEkkyb9GGsrY1ldW4cDc9UqP2Vxe8xIuuDKSv1UKtM
tPesMXm/kORj5+I1bymtWxFjWHkfbEjl+PPEdJxSY8tK2Vz+6gohh3qL8bvmYdFNgfaumSt3p+jr
/AC90xPyq3qnIadJ33x4+w/GvM4IkOOavZ7I5QcuwTBRG81ee9VIxFU4b96TIZyEcdEVUgSKZauW
zAaDfZ/0xAl7ZrlQHvCqqzhD+ZIrv5Qe6Dg/xR/TA7WFU/DI8BPuq0wTmlLzY7KWfvTogfI5K/aV
wwjz76H0tQoV60hHrVsNo8vwA/OXTn/ULuZaUiBQZHHJH/gUdF45j/KWTt25891e4vg+Em+rLKIV
C1zOdFPVTf0e+Ux/T8PPNfHs8FzT2mG6/5j53zfzkqzT56eYLPejfjugJD1Zgm5q2CierDyJp4Vy
/HCmkF+86zldwiHCTriQxyRdEn1jrWM3EHir4VqUSU/hAJX1DD6Udh/3ksrw344NFxU05BoWwXUv
/fk3GB6hm2sGZFMfIW7oQuDqp9Kd1QvUjbqekBBT2vlDCrCyTqQKaATqzwHEJ9TsLbI1nunJG6Mz
ehvlMzR9iYLkGU1emiDD490AeCam4GbGk5j7AEWxhc77XNKMN8ZGY4RR3VRaXk5G/JMePvVUc7LV
IVX58onK7S/eVmMQ6ooz+JG6ckJPLqr3GTwmyk/ixjgbABGeAHQTkyxQAJFDmNRjub+zyYVnm71A
nwZ5/gSx6wXw7x9NoraXfqlNINuqk49MadKofbq5MvJYs2h4FNdrtd0hI7UC8DQG5AKGqgWn7iKC
gA/kakmO2K8tPGvtqWU8bHTTeBVhWu4rLLdTrgRogNeUEDno1uVWcaIOE4ofENckEobD0FKoIbxz
AHOoJQFoA1RUpuHQFQjyOLDrSnryfjrT3Vio0bi7oHCUeY2XP/XbPjlrTced0KFbNYB4MjBukxPY
QQlyOdSyA7wCJ+v/ARaDwrI+ocJsky82WJ+q8J49R2AzFvJokiRWZeD8U0fk/mUNtGMdpbLv8hFG
jEBzSFrV5bym0aT1X59teJfUqis5OhFzhwME4neiWBAGgCGaLsG1Ip1raj3BpY95iRy96MJf3YSr
OGR7tWVunXSzicL5EMewlhVzgevWt5DkYiK7vWCqbJTct34ROmVr1jBbehFCMdYtC1Y15aV/NbGn
FiZeUa2lKE7zlXu+q0yY8vuNOANKmLn6Vt9C9QePC5FV5zCu1idxNlspGGbFVKavR/SqlyGP97vX
iCTudv7weyBilo3zOEHbknuJ4StpYVXNPXP+Ad9fTV4og/IIfD83K674sjEUqSOMMQ/BrFeaxGgl
gVCCMMTUTTzZdkncopQlNK7Y6YJdWhuer9qV7RZCfv+/JQmR/cEBoG6oVHzyTNnxZ3dJVKGXJlOn
vFYordbh4mGp5ve4uKnyeh2+3QoOVQiIdvfxg7+Jl3joFLNZ9p5eZi3220PH8AfjmunRUNPcpk5D
D9qu6DgSVh9mw70thX178U5lHJ2NYsM3JfGc95Bs94ddyScB+hB+JU6EwTG6pYroEnRJ/trCsBps
xzKMJpkC5wge8Hwp3z18QC4WFgWD1yW4jVnbt7LxM0iQ7+aCykGEiIvoUVn2E/Q1kQXUL2Uvtm5w
vZFKuPaK69tRNm1gENx63KA29z8PIuFQ8yfKAYIZ0+mJCAg9O2sDgmQ1mMz9wXv9YBVEopUi6jiu
qPBQmQLhFzTeLhyvNbJiLNnUC4hGrQX6ErzQkKoadsGCTZnnQnO8WlEk+ooCXDdHBFoTUgdd4+pp
pHC4bH1LeotKDWtGHGNMO95A0wo63i94m4Qle2zn05RaiBNhbFx42afEwH5BMPsDQNEZpeLc6SVy
bZmlWG8CYkigc3Z9tu7bGaB3dTs3WXgWQ2irHy9mnQom4FFeEcO4MiLZ3gAsICl2xqgDi7jcY08r
fAQDGFP2q8JE6ZXfNkesd7WMwRSwnqnEqknnVWww2XodqNuvqU1Zx3OnG4VkabQ9QGc2HZM7J7cx
8x4AqwWR4/f8te4MNW3pw2IEWcMsrQCOpf1e9G4Kohs6P1YsWHuulfLNLtC0l8nwTviiMwBNEDkG
b3IJeBA4YINRrS+nWixNpzvYaXZRE3eFt54hsesICUIOoq+ZXwgTT25c/aFxCbS1F1mypQioUJuf
Lmcha16MN8cLKjW3lL9lWTu7R7lTCSqVbFPFucL0ZCHDpHK3V3/mUxj1Jh6xzvs6gw+LapArwxsf
d5zRNuJbkpakFr3UWackSmCAGveE0lo8dLYMEMRSux6Lpyy0863MW9vDW7Sh0j0uFhT6FvveneGj
JnwzxrwYgzxC/5/CqARch9ZfUaV7GLL7bHCkfHn/C28hn7Jbeg0jETAwHumADE9aS+FJSG9JKzcX
Cdns8+Z+eurNeEmKCkpQaRjcb5YhfI47xzOuk4xFQCfcsOf4HwtKCqa9RRhQXy/J3elmgW9xRvwg
kL77NyRAjcgIdAdT6JG8sur2GG8V0cNEJDviVNXCidImgI58ubjs0rQsXKvlpL1+xn2qVJK36tGd
4dk7iZz03kftO6fJdGkCbu3BmU/fAeF7F4xwaUOxBA+ohcwBdPK8LCnDKMuUTdX1yNuJVFwg4yPH
sLd3pvYy1lOIUqrhLQ8DCOP2W3SG57kkkqFa5+bTN4Bfey3fAjbDgotIZAvXwX16jpXnuPI75sx3
AzQYusdtrh4tHrY1crvgdYErpyFheE5ZUTutZiqfzyhZZ6ONxFpZKYMqvEpUJq8Z8vfUT961oy4w
K9+XgRe3lsg+6XDVUmFUs5dLkiQj72bvTgiXfO+e6oRWaXd9jCXH5TQNgZmqqWaGse811xITrW4O
8m85cS/2RO4yV3FCjkUMPcn29+ClOZ3N90wWOVCCtVxwhKuLB7NMmz0g1d8vy6pDF5C6EyIH4GUu
Fngpco4g4RR+AEHD9guih6LCvSlmieQZ9Ugw3UbVPvE/QhjoEU9mWZDtKzR7ps5MlNW0o/gKww3N
1yKRcbAHuhE9Lnc5+JIdwi+sK7gA2mLvCbedWWtclFE4NFu4TlDzQiMLSuhN+kAXvwlCeYFVY8G6
/tXrQiaS4/4UpEdz7S6H7cmNwmSM/Mhe9U2DD4AKGSCZN/jxNqBMi40+VO5CFv9CEmC27nQFprhJ
pJRNxv11Ws9qTwG1kOKbBx49DJ1iwHlDM8hTzcWEvRgTiivPMC279dE2icEq1L70INax6Wbet9N4
QRjGQmWJDtUyCJa0nMtcqSMTl0/jcE9EemSNA3ybzAAbAwh7tCtgiiBdGuyswKb5kUZgJ343aOaA
3V+Du6wOFgmlZ4daQEb8Gi2JcdfqUNFR1IDFrHG4gurDbl4r1KdMeehCgFNnGR/CKz0L8wCsMS8Q
NQPUSyinDszMMjXgQz6g8zf65Nk738a6epcMGQLA0iLU1ObB3yrt0EOnTYpcMdtqHm9XVwDxHvrs
ypFmZdTSy1FS/ox0+IqifhThOhb19TTyc971noPWF9+GlY75wGGZoyO9sZXEKNUkHIUDB14fQ/V6
g9GaO/4S98roVLdRi3++rLJwRyzo4oaTVoN9eFTDBk57MHYsrVZrjEiOAz2NnHm4wo1VHw54phkI
Kyp7j+cAHt+n2SCOn+a8QBxf7EdwFN8W9YZBOCj4Ps595QHHQOExhvusy+Mtn67DFrxgz1zAHifr
fCHJpW+yTiPn6aq5GZBY+tQpd0OOxbaJ1fb+zyRuCNzz0fv+2Wh8TkOs8n5ZuzWC46lo4C8Rx+gJ
8Na6kcs9nOBZlANtq2381oseKqbrK2DfZJIm6zkZjuT+rFVO2iY84XH4LBqyEttQ6xxNE/g/1s4o
EsGg6/a7kgNmnz9Ik4TNyXlPI2xAJ8Pn3gCQcLQI6x7X81k7MwP84RChXJKuy1wkgUuSWJ+8/Pk/
Phgsh+JfnMJWGCsNSbDIrRb6Rz25TWK76OB97ccTbqwVoSYyz26BqfVyorSKZ2plRLKzRSf3NnAi
qR6l7zQJ/rD07DLgtTKhPCt5eP/VaTafBIkZjbE61eDkUJ9Z+KpMn9/bRnOHnCH8Aqjygne0ejzM
axtT/QQcqlLIqnUmnW14gcnBSxGchj6dq8dqzc0cTlMfK2Q2jfu3JjKeGpxz/crV1Q9mjoug39Nf
yZkTYOIsLOqTTqv/Fb7rqbTZ2cQXrM0kTaBkYE1079THjxMssxJBBWAGey41tP1WLPD5U+yrs1nO
4ur8PeZ7z4SWUPmncCJNXZgBUzf4PAwt+F9W1FVGl/xiiKSNv8nrj8ZWuIuJtt9kKTSP+ayx4wLl
syz5rlbJx8SOgbOL+9i/1SrC03K/ttwPGgPFqGnqp3eYoyjxnKJEXoKZr6O4iOg3n+YRxQE/HOr5
Seu6VNzP3/sLPQgI01sHSofagX8VRSxzNSQdoi6MLdhyKkAWNRWnpKaGwQyoLpwDK5MStQ+FeEOQ
+dKmBUNCsufR1v67cU+T8/hymoPMbVhEST9fhId+l4hCoAT7FnloVPx39akKkYekwOrjL3O2p2Ih
vd22A4O7tsXloIlTusENMgKcvTE2I9GVj3ioY0vwgfXiproTQ5hJQwP6hzYxqi6Ht4E0xtgvvb/r
bzvXMoehIKgmLNZOFxtV/JM1hVSIMj2zoAsCkHj+Ea6Ky9wGb/Ud0y7zgMa5UNSXHYzhe4VwS2am
GrV5NL3dp6dylHyC6IfAAYVM1gZyaR+CmnELTPE2MO83e519Xhdwd8EDvL0dXAvmsBv4y66ATbQP
0ACVVbSjtSdfjPzfDGJdHA/6IfsoihdV1AV2Qo+CpFSFYANxdXqpY1loT+EMz/bp54K3AuhtvIt0
8JuFex6C6Fy+dl0/xiA6FQCtKAzBdOq91HVbz0FYNsRK6XKimh3TgqoDxHt5RoQKHodjSomeZi+u
2rNks2po3pKJ7S8kTmGHx4MSxMK1axP++E5kNgp7gOJ+xJFX1qWNyTtykI29MyHy0e0uuq6ZGD3R
hHN2IrLJJwnuC7YLg56NT2Pe74W0ULtO7rWZ//M22hREew24jy5rY4HcOmsUkZME6hu0m3K0Zm3b
qpSUD9y+je+DKTiICV6wmOw3W3OjPYS8qCkUyxN2QjL5B3Ey6Ds3Ban9rjaxN9u4t/mnVvUc/yur
V1dVXBSxNbK8bsPTNvdDfjrqnwmeh30P31CniR9jF7Jhnr0B7z79RcAoPgMrMfWD69D17+Y4Z5D9
Yv7UZK/xM6EqBFRKkvuix+sp90jP6nzCRtCT8B3LB5oBu0VQkB5sya9B4c8pL6mhecL6j50TjKL2
QpoI+18c1AQuFpP8MIxDoyv/SiSpSx3wZeARkol30PNaEO0bHqTV7OY6ntJSKEn2RY9J0SVhXOHJ
FZwzm8fcKlxpoOs7mzgOlHbattvfYVZbWJTZwN3obvDGC0/K/nC6A5J3LjljigQvGSOjZTZOudbi
4Wsqcl4nW2YMitRSMYhlU2/DTboyfhPjZeR0/5soKKYD3/1HYJLaINXiuf39gBfiGQPGhnfHCsFa
cJpSofubFXwEE33DKDeiMM6xh9aB+FSiednUYjcnY843NbslFa8FCR7/sbM38EWOBcVTfDbik9W7
QDOjuc0Iuf1hj8r3NZQ8t4Krvz2Jg/eSHZenD4zudjazV+Z6dgVuBmg6SuiHAm//PwgJANBY48J0
9rVAjZlO0DrfTVc35Qm8Z76JEaF3PPonAsPN66/Kb5SQQ2zBdIxVOokAMhBjn5DtYrasuzb/X/+c
skK7drQVJ6S4GWUv2E+8nGMxtCVBXeSprtYfSltcm05gmJfDeEPssuG6ixJV2Q8of1VmE2Fsgq04
nHAFCjcW4alsuv3niyaMB69Ai8numAhPTeMiRvr0NFfzaPwp75z5w3UK7dp+kalzKAyPGVB/MHae
lZ79FDF44YgAkiItzceAPoGzMqpEz97jBrij204YG/PMIIheFmYEdxPNQ14slkQprVpnnX+1S9rA
FTZUxjUMf9ERuTnvS2jb7Tvx41c4UOtkEiqDuDTtottYzsWqXQUYMPgeScDMHcVFLUny4j1XN4JF
CK78iVAlqNvSbQIwwRpWrk1JZfDcvrVSnH/NVgwWxMwvwRkQ2LGlZSsFjNuvGJI01508kvy9mtSW
nVqYWt9ciOY8efAsUKSXR5iovcavvTMdT1PJoJenrpD6lUhJeQbdBE3xVUDVFR/lmgg1wzFnFaS9
6zXIEI/JiBUfEZKoSS3rbdtwG69R3gDsOWgx5NUZMupMYd2wRFjmyrv7NV22oFtedmYzSnZ6yPQ0
067/oKhsQTuLox6Oiw4pYqmj6nn8ZARM+Ax2Ihe3Sa/Nicx6jG3wUFRf3Ve0n74unC/xhcHByFp9
bTFn07uzuy7LoC7lNW//GmNaBWW4SWY6Osj6o72DfCByZTlubs8412bWsouwWGw3vY8yCPHcXuY+
IR/6dgSJY0f1hVDk3wzgQCsj9JYG8JWCC77h8CHsjOUM2EQXgEK/3XATj736IdP6QjIprd7GQ0N5
6IuDeNr8Y20f7YdpXnVwGifuuOpaP0bWuj7/jqTvHGgA2dWebGKT//dgLnTmUsdmjg1pZOtjtSCo
W9kY/R9eOwQRxlII2qkYnIOQzYrKdprRGUBs9qrc8IXTEPqDeqcK1yxS9Rr6pJmZIVSOOt7Zakan
f6mXj/InMVr0rU++tuYua8UfNw52uDVaDdxTq5LEX9d2Z+JC7tq+27qijEedv+O7Wwv1KGHblo17
7i3Jihr+ZHN52ib97JmoeT2e5FgYGFASXJFSLqgUTRK2dknywS6MDwxiO8cBjVNishho6gyfFmcG
SKBr/hGif6y6KfnO7PawzKLthWQjy28aKy7O7nzrCSLidMmH4YYgWgcDW9Vqh7SnyY6THvurQ0H5
3qmJIL6ZrSW6LpYXIRLF5ozhr+Ikm6NgdMcQ9KqJ4s0AYtQf9Wh3cCiMI0nvaEKlXjA/F2J521KA
b3l5Ysi1viZC/Ml/hMYPuTMX75voY0QWeruUJF5zSm3GiE5XOrjqOWgNShaZwIJJ+w9oGL5PGAyr
rjzK8kxGDJpEATI8/hs5mQqqJgb9Te5isVKrdfibQhYZzB8bBwQBKXqrae7V97NJ+otm5ZS8i5By
E4al6YQMHK+HYTdhYqxzK5427X1jaKh8/vFXnBCt5RXhRfjEee9fc1VgqfaykZBTMCrwCoG3Rogr
8Whc/2XWtFikgjLgFY8dqw5HfkN+SEaCpXPHqgo92Zs2TWP11+OQB3AoKqdi9ZcgD+k1Y6k83obk
ENcpPhzztMydhZIPgFPgYh1inLu4xaOqBgRjxQvh0rAujNaiX/rl3f1n47Rkv2+b2RO/0UjfexC2
SHF3cXnqA6IgSaqnBMgSDv2ZMq0w1b8Nox4OWBG9GfrZsBCjmqS/0+UwFzmcYNovYx95Nl6NWNPy
IExC9/mP7UHa0Gq7vt4ftSyxrQaEOrWu67SBqxBgxGh/gxX+KOCTSAxpUzxfEiExd7oV9OJQQG1u
8offdwwTO7Vfi3OoYK8Rx8wC87uwC419ugTp/lQp/Bao+U+KkV38gidOJp/2f2At1IFrcSpAL46e
j04Ryo/bYva6qENh34AtleOdi/ybZzumb2fSEO9cfUzjPfoy8hHIHgN6o3W67IKoMBlI5GF+h+su
iUTKrzNG0vNjJolVDiG+5ieXYhWHaprQKhU4SMKYN6hZZcRDU2nkdyArM/TYONWhY2Q+EFcrfjN5
7EeI9cA/MCh8tG73+XXHhvbLv/KeiG/OoEh0vMy70jBJVRnEj3/i9R6G1rYhiq9jYTowzbaTHCVy
UOCFwZL2lE1VyZSkAh1Q800vRTbKY3v9uOFP1hd5mtLYoeDGiGZYOA89c3/CbWzPNWj5q5Y7PXsH
US2OSDZRw6aUxblyuWD7quL6q2uvyd27pSplKb5Jye92JB2KKjlTYoBhB3fOd7eN6UcsQAFDyMbg
aO5W+CMYNd6b5DdEY73JAhcCRIW6EUYaB6D0flTECGqG1Ss/eSgFr4OmTvFqq/AvpLApWmbMz5cp
9ooIbD9Thhx1qFZs72vrFlhoVNTrF+48Ky6kFURV0GzQIkRQ2ulit5pH7AaM9Ql7jilOdB1cnkd8
7MK16LMLzBlrOcxtzBkCZnvwR6WDhVYfGdzoTiGlooER2C6s3BJdF9664ys7r2/HqVIVK/umhy4j
FHRc9F60wOp4atf0DtFWCZkYB1PCHeIuFJnhWMY2fxDxTijPhzwlr/CYp1nDJZ0kna5yWsRsP0CX
UV5bJZr6m0uM6DReBG80KDEZu0sjSkzV7BIyBwFWkwGa8Pd5zVbMUqqbGAvkPUm4Gs1unGJzKOIM
WIo08+Bv1tpTDn2gvMlbljdEdrkwFbKzPlpw+DpFxIk7aPwD4j5F0C2uSHKuPcfu1hByOMkqGEjc
Zs4BVT+KuLQi6AH5JK11fTfwY0rg1NPb8W1R0Q+mASe014e2HikJb41lH0407cNnDW4PflkwQ/w6
dORugmiokNKDNUv4jScb+l42OHy+ryhSNXvOAlP9AxcmiXeZHzM+869K0foPS0Lz+vkJiWAJFLVQ
er1240yyqSFs6xBwtj+t7yvyp8SeFyffX0r+NQVi4/Er30rmdbxocTqwLfGi2ah7N0whbaDA2LSB
qFRLs3cTkmJ/x4+KC+yT9Wgvq7vETKPqs64VnrwNA4C38I4gYVnePxjmV8Nafgw0Jasa4jark6kp
P13Q6rjtnYpN4hgDDzQgK2+gE4Q3zMUcMx1UVOL8QVZNR3S7A9RaNxWgfq7cOjAnuA2dZD/z6e4i
NBxWZzeI9W8vkKSLygXdMoaiDnnRH7GXiX15ZJ7XFCXMgHKTLy8oRohEselgU9epbLHxzkZLfkAO
VKIuWbFl8TGJKWzyJ+nldu/RIovn8QR7OgIKw2au6J4UMLkjjjZUC4pgrnkYrvO2B5cx9hr66dyC
hJMeSTvV+7Y6Knh0EdEcfDvT/WiX3eLlLycWTI3zRdYBq+Z047a5/9rGRv5Z6OXSUTBFOY4UYZG/
dTRh8RqNkafV2u53soeIaJVONiAtFE0iFZKM9zQSg2HXGWxswskvhjkAri1CS6zhoiXr53deVO4M
/YoOStKI6HSy01r0SCraNtdSI0yhwBe+3hpAvgCBcgxVbib0q334qxuYnOtS1ygs5jfENkIHnvQO
xTFhIk1JUXOZ7WJrTuMRVHSZXLSpT0dhiiJRIOOfkF5CJdbJnNfOg/iMBejHZAUQuxOkeKQKwpUW
7qaG4lFbVPMqMCpBzSKln6PQXtBtde4KP9/1HtypCFfGssuPUuFlVn2FwRmk0CrH6nnd24IpvFd9
pGW+P4CI5NZPZcCGdMW1CaKvj21anIIpv5zMfsOBuL6iW2QP1vg2sYZUYReCfXzntnEyYqne7o47
LkNw451hrvGUXPD8TP+g1bmnQqfnH1RJT4CJjsk78RqR9WHFXhgsTeS5lr4kpC+l/ugK7qZ/Uyxn
OUPrpHlbNVdXBDSJTILeM7XZTT3aTg1q5eTS2yPbXVTx+0pG1K8X4tscvij2EbEf6b4qPsIBgdbt
r0wFSIZZJTz+3k6jKFQoNtJdGx+S2R3OX+x8CfaA4vsxE5rCFFjiHkFF+vX6XvHaStgUvC7ZteQ0
G6iifqyD0G4/nUIHRbt8j8QEBD5MTFiRe/g2Vo7D/+N80WqX7F9vq4N6MkgnTuFeD9nZNY6QSshC
tGERbSUiwyBIJdxXAe9hV9HfaMM5q9MXIYBxb51Lb/wRy/KKzFlm4LbtrzFUP+bv1QKhgtAX8qd5
5hdPkLfJ2BpYqh1BmhO26utxgMp55Ute45GvLUq/uUUJmd9fLarm+enB9dExjZetEwD5vBhp5qoD
NtQvRfwSDn5qlxZkVE+gugZQ0wlRRLijhMwInH1KFVK495s+g6yfRACoHHWTN6kfVz01fkpSZL6h
SMQIl68+PfN+bZZeQQpni8srQMddXr6DB5DbIf2UKKtphZInCxHQZH1zV+3E/q9mun/qCrU0zang
Z9ej6vh5xI0y+dm1bqno1zr+JWlJCNW5b8fNvbRef+m7LLmquMrn+foWZiUGtWf3EM5F3v3iVmNW
M6Nxd/VIZzv3n62ARtU/gS7JRQSvz+Ub0xK6IWAmRBzZEyGLljScFfeUSU1Dyi4ighHyaT+ChDnC
+uOnX3gLf1sNrmcGHMqy1Dos1UkBqiFApvlOuEZmgVsLS83iI3+KsI5ZBd4PnlDYaLuc0ZaWUy+H
gVnIuzSuR5BL7FxxtVwRHZtjhvTCsJCE5vpd4xyoxbnEQc02nj6pJV0z2VJy+StWfKal5ErdqPXK
9wipMUdYeZ9k7983FtWOIMcPOlJ4+gGsNipRc2kX1NFw1DvNOC590FmQlCClXul12lUnS7WG2PP1
BJk5wl6omDyGONIaWf3Zut9NYS9KfxQjXCXs/0Vs4cv9g0jeKr23Nv/zU2FZ3bgu5QhcD80vbvDq
4U6UDljXBO5v8/eN3IqKK2S2/fVFT8roII/EiTvQk0pjUv0KWo4WT/s3wLVHz44lJoOWV3njuzqE
aZWgW4uV5fbsX53eMv78BJyKfSJank9+qx7wteirafevyLqhJXXE0RvDNCiDNycLIn6GaN2c2PWY
vNzl8PIP740fGpkokjNKqUDvJ2TDwUaIKbkaq9goKM7oqaIdQnp8LPZED2bWhtyQa6xqoshl5zyp
1QSTpgACdpTRXcYR9tN3tWpdeN3DChchBFPHvdTjmbL9gt5Qu4lKoIfh/F8sSTo6fKssTHrhKL6J
x+3WO+c5/kgz2xVglZ1RXEP3pb2yY3mhkGYZIQKeZ+qCSfUS/+0QfYl0yzchLikCnWI9p8ojnZkn
jkQcUVAmImhLvszCDekLF9/ap2GUIyeCFpOw/R6nrd2UWRVcBIceF1n1gylvXyDuwKRFMUS5bYSa
RWdBioNwdiJkd3Y653cs3CO/NJOfP1vfGkJUpDYRKMoshs0WmYrq0jVaSD4P3LCgd2yxvtlzI154
7/wkydg+MKQ36YQZisSEYNgyxFRvrXImx1ivTxi3uz9QGUsifOplicz3g+WjzAMjeuFF9SMPoCXq
hTeNn0FEE1lqPUnFj1+P2zp1XWNN3rwlbAZmMjULWzoUtvT3FxEpOn+NxbuxpNyhXv5EQzPNx0vc
XhdRLA3Mg3sRtB1jKdlNnuSxIJuWOka/CdxLlkCvj5xrd1tA2wVSehBDrKq8rsLIeeJsdqeko2qw
lonUlu7bKgKPXg9qt4C1SJrEgmomPrzD8U0qg7BFZuI8WE1kvBF8oYdVpJtZ9nHeh/ccFtqEb71Q
2k8xbTf5hm61OnEPCL1+JNHcR6Yif//XrHTmSJMBI9P76M12VFak8UureTUek8Iz3XDmF92oLoeo
7Bt76bT0qsncdlX0iUcOaMhoXAngXZ/xrQvO1/bsY5k5Rt8zU1WFsITgqtx6469qo9kfVXXbtRF6
y2VBFZ7mjBp0rQZ8NVrxlYHoG0vXZCw6O2ymnW4JaKcJnbJ3GNA7oVQVSzMJ+8T/Sz6ou2o9tnjO
SB5UNjkamxBk/S2feudx5WZoguy5PBrM0frV+5z4dkXPp4intN+NX7MUAVBanyEEjhw0SzPOXZPM
0T79V0E+I5u0KIqpSi/ZGT0vmeiQebStqH8Px3tP0qvFfNDwmbf53Ril9RrhCSkmvk7MA57MEJp/
Y9hXLl0QO9ksi3A6/2x7rstQJI/b/H0x4zCg3YPqqBSGvSzOx0mbOxIngIrM+86ToekUlLCuyXtY
rv38KcU/hUIfByQ57t9UkX/rSOrQJJh51f6U3f2llVvo89xCnCB3asrJKTOyO7kE3fJYCN/PKlDp
PkWwkLtuCGysJPrsUrBFEPxygNp21WaSJeziWDaOhEPr1wQoKtNRMuL9ufsHS3DpKg+ta095VEgp
aSqqGjGr4bzW2Qffm32UrtktALofzcrkW5d+pb8cte8PuGjswrlfU7R2hFMQ2q2x3F/yyDzer8RF
ZbNv5TIJdfladIpnkeCbXiFp60jT5F/UjTTQpMFTbNRJ/UP3G2a0A/s7n08hZ5z2Y2Z5i1D6RGmW
W2PvdTvAhEIywPs1U5hLtBA45E0sYPMqDZpX1BjvSsZ0mbv5C4/ErfobG/FYVUX3sZf5GCptqpQL
q1/SbaRFUrexE3nuwqxt41385vYOCt0q/8cutE5joWpQuuMwZ9HDgldR/O3YNYSnWohoEP81gO6t
UtF9gEyqngy6Xp1AN1v6TclslyIO9pawhzjRT6zUSywwYDWccM2qpdYVO/yLLo4vMSGo/3FJ2Ze9
bHcKYL7vLgjxJHF6fstgZCQk51iDDnvx3q+fpqCTlvQSGEScUCpW69HQBMTUHFgcoJsxLLHrkuKB
LGdA5G6/hQZU22hOcnhe1MX1ZlB2SrA1SRo0fjBol5byhvpiGvrjUdo3WTIUAo5B921JU7yZNweW
zCQ4CcNzO8vWjF2qHZ1/v7VzquXgh6Gi96kVq2v/9bxjYh7Gbgf/fZV3+SBs0IJEk+XKNF2XDMP5
0XPSvQ+17pv+OLf0Cqy82dDTGNC6+g+x8JDYXkX2Wr6I7Tr6vF8Ao/PVkY3eNY7TAm86+SyqNcva
E5qnGVXKtovPUXsSCEjAzCHn973G0O1VwjYI4wFQe86AhD1EdIXThWvkavXpLMQ+kRo3z22VRNLL
fxWHxKWWARFjD2IrXJAvH4SDp7hJ+h92UvGxKDAuAyehjDUuNrj/MlHjq9qqnZMeX81plujmcxD3
tzzB78xVJTMt3y81c/o4/a4N7XlhWwPDpDtiJFNJlw/JwQSglXiI6My4AWTzF+pglVq7eTGKIguw
GL+v21ImKxfF1gUTw07j/eq15n9rE9/Fq910DLqzQXkoL3ilIfZuIAbhUtpYZLZu/QK1aMEIgj0o
y4X8MSDYJ6XBGRzL+ZwyK4EzDn4QT+Ftu5jKWfiTgSys2r4mvLup+So61etIoogGV1BxCBLO81Ux
D5Z9In6VAV02f2rlpxFGXct671u3te4ZgxWZ4U5jzI1zMq3vZ5VlzFeKvLUibhaoBQl2dFWmTJXd
pVYAOoHC7bQjqweG++GVYcWxFLNNfON69M+2E7SOwTEejG3oO+yvaYZU8xbJT63W+7aX24FaCG7v
wwjxzuH3wOGN2YrgH3HzFHkDe/BGn4Y9bKNjMbeP6PX7PD5QU/pWxFv7UcdpRRmUBs9pXzXXqUVO
l1HkhZS9/aXQWFe7ZbdaiEyiEtp6CVkKQBldl+U5g0XPHu3zPwT9pDGA8EVNnxQrBsM06RUJYM86
hy/d3mI7C7TELWQl1O2k5qZa5efMT7DLOIC4KuqPiPXs4muKCHmZq6J5J6KGcd0uilPeeX4KWpGB
ZQBrnBTcMpPl9NppN0I6vq2JLVdJO2i8MnL34P/5xNVHJwi+GzoIZ953El77OwEd72JWisR9OUju
tj2lcWFOXqeV3OTZecIMoSqi30UM4asZKWyOE0jm+2MQ2DoMNk3JWlXiGX6nbNYm0/XCLpii/x6U
wAAWvFkCMhOn6rD/+fS2ATJHDPaum70wBEf9uVL4c7XGUr2S9ekz0cn7EQZe6DmzuKAq+ak7Lvht
IIVvQGGaKpJxFipc0y3/iqW4w0l2tMDAdTEi3aj+wxsTPVAoOgf/TC6/9EcQVcOSouBjk3NAl1el
qPRnxz+NBYtuLh+oOmibICIrhgnYCUI9RksmdzIaI0O6z4aO6We2AwRigb5oBCQ//mmcmldTpZHU
c+BEJcMn4MbgpB9fHCrqeHK4nF4Yz9IgHUmjgKofN0urAzJGSP7apWTkHnzgojYX0fJBngTRpXTP
tLDT8V2hzS0AkLOvigM1ta4JHaYItaJ46ae5sT6j7CgSAZVkcn9Whp+DkkMwv+Vqm0Zzak3TvE/c
jo1tPRYPDl/qLvwWFmzqFA2x91YADmCVyiq7fXYdNWyuuES63jjHkSvs+BTZ34dhqO5+LHsS5mVx
dexZoCPjS3tcezg5y22E8oSp4qYJj7me/foIk25SJVQdcJEIciOGG3XjyN9sdAhDEV5E6lLA5aG8
3xBOPvscdkLOLfSzyla+egqry2bdMsmk/VWFIwAp+uBv7DwiEPmgeTdfm3dY+z3NXr6LwXoQqrXM
7lM4PiAij6122aLGy05TOS6TaBUWncZopPt/S76BVXTO3BBH0LItGtytcV0VVY2dmgXcyx7Ymioa
IrK8OoC23scmjsnxYjE/aY7bMbMkVJTb/c+XT6e183VDk3q2jzz1umTw8F7UzbEHKADlom+jIHep
IixUUnT4/adnup4fSnMuH0GUUA3A411wOK3fhfpy/7vA1lfCfIvEM57SlKbqgquZrltRRDJzCK3o
64e7jnabf1HzRPE/t2EuVxDFezue/wPOi8/fZcUN3KI4KI/3oLYnirscVRGcyUWcFXVmkxQbFej9
Tvlk4Hc2mOtJGadqIrpeu1aGIMQkEJ/tq5xXnmv27oYHapWhsARndRyiuqP3A9yhPCIphskcE6iW
XKijHUBFTqPs0H6isekstFCEIKkYGeNXTxGwlIvUfkmClxYJTbbIhSYrD3zJrr5YNNNZkW4fdemE
Is1tPX7da0e9z4tE3Wwqn8vkB8xjDVg4PCKgVPsLvSDvebKULKflH49jXiTZyd1AafypjG/Sp/YS
oK0FAcNmOfH7BZVwIgsVNfTtpJvozh6W3d6t6bJLE6BKJOGUAIsGD09qjSYGOhvxjKEjyVfc+zxb
b4iwBI9rL0542n+ZNmDJvvfRfKokjIo34/nDKZJxI591AtHNydZBgXSWAeUoTbAMH/LDQX6JZ9pm
nDYtY7qY9XAmKRTCeAehJaon0F7c3IzW1Qpvex1Y7N/+/ljsAufJkmH2NnfY7XzbX+eSYp+dbBgn
MtDK6o9JzRSxLoxKDd7Nxs+ERTirCeR4LxojdMawmjAP1bHYBD0XGy/aU5kl/rfBC8S5yTihRd/9
OpsjYrWFf0CGujadFaY2b3ccdFinshJqrS3gkzFOFmax/BGJuWGkGwl/D5jzYk+mlCBSBEYXDnK7
PdPNyRLIY6pVo9T2rK6lEhzKgtAMnS2engX6bYl1ma/PDSNSMA7QKuwK8k88rV48NB37DOSeDler
rpy8nOxwQUuhLDQmiblRX0QefrDL7ximEDEexoChL14CUd0bar4n5DFZzQAhOND8b/qTaZTFpx2W
Qy0dubKCbQo/EYhMOvsX8JY1Wxh/RTQshxmkdKY6eJgTlPsoUkThyQhHR9+JsdiZQ+bM4jxRUUyv
609qwYyWiXMvjWt1pHc5UyPuCyc56722h17Tk29iIsWmQJn6z9PmKSr6tXHXoNwctRF8sgfSnFoF
wNt7KBF7+YmLPyDHujyfDGpJDI5IQbBqPJDx4HsMrXac4pBnqltI7joM8VKy7AKBwQziE8WEHFp3
VMUAra9lXDA3jyrBnaADgkHkfRw175qZIcZa+pz/BjqQC8QqAOy357rHcGdDw7EJBsnBq8RI9s4G
3V6s8nT7D9qu5+4ZB05uUk5SghKgS4f8Pjtpf2Y/hU8ZpkDzmBj2v8WmHNzaIoAXXwo8v5EpyLaF
ujknsCLdgWtraKxgp9+Xb4HKPD76K03nYUJlv0pi38bEEgBaLa4RNAl5pGICk5YreCe1naFftpl5
dwFa0U8kYYVaLQAOfZ7BD6jis+lmv3Rm/rzevZ698ISC6RaNzjRap8uTMAf6ZPuRe2A7/1Q+RSu/
Mem02oAFR8JLhiW479wr+nTlbe6yPAHwnTEbRynmWLNm7Eq4/htUfqLaNJJ5073rZfAlGy8b+Qf0
qyAES+z1OFSM/XW8yIc5wtTs9C+o43Str/VWyH4K0vMtWF7mK6vYHa3RC5QfdiBQCmu9J+UTadmb
845WhXS2m/5olpulczglW5xxAbjZafEJIz+0ygAb19suMr4fT3slLA8PSp0FEMuRPkgnGXCdlmLl
U+dz9MhCvo3dxer9Ft/MSiMWyfA600oDlGXo+A7qnZNrg6nTNmvC0N+Wrc/JDVBm/Teh7jgcIDwM
qY7ihOV09jdRCkguhNzJPRsGbZTRcvN1QYuDmjbfc/9tOzsuCI3VFEaypJCZge9nlLPgL4q9rxLS
Wy1PC5TK1vSOl1JDjONW0qZrMozoF+in1yyKH6mqQ+Lq2AU3mbuUXHKDrBJbbX/HWQ82TapIa9xV
38J5+luXHS1wrpyZKzJ8+Fp/e8CKi1oVTAmZxzGaAsMEhPLeweX/15dg24ngYLS7ZbrpBEs62/5F
gZ96xzklM3+GgknecsjMB8UyK5i3d92ZISTzktyVlVauLeFj55hEZsk3M0ZcO3AazA/gLJGxbBcV
QAqNOLp+DYdNKZuOgEyBrtjkDvHRigyGAwH8z0yN6DnVE4SiPKttvPc6ZQ1cTz5ba3cQ0eeU0D75
sft7uIDDw1DNFDEjT94ZyE4I0CsOF49IcgyOCO32Mr5smVN3yiSIQYnw6nuxC7fUu8LRQT7zzVpK
TbIcO7NJxLBq+irhJz9ewexptq5B0BPxHd2zMyvZ8QdoqKPne8Svh89oEtDBE6zMw9gGnrzA4fX8
iCQTCsDoUtCp0qpUIP6Awxa2oNvQyLjzFXKOhK4mT3QKtAmRI3OG9xJiLrRRtsX4Cj7nmB6idt0w
NjXaKMAAHAx2Lu40N22+FoEsSA2Fj1NSHweRF9zXwj4FhdqjCfNkzTtyOkl1d2Rv9kTMiIMiOgPQ
rDrb/lZcG3QAHI4kPgykhNbCdqrWOaJ+BDuP6K6yhsxhulBdlLHvM+21NYXYPvQYMk2QZCR4zuxI
Pgf5I/0oR1u1y8EHRGNRI9vkyhGJ69a+JVszKqDfgL6kNfgmC/tCcasTRYP8dUi8Mp3JQUMeozBt
fasI8b+r6AH8B9Y3Y404IlsOq2dICyFg5T5VCgYAosA9xk8sGnbq5eb6w0EH4jZTdS16Rx5+Z0Yv
xmHiEWc82RIGJYisOh4Vo+fArP8Cu9ako+9PRxIKzP9mvO2BrLML8CxUnJVB/5tDOI/Pa3pnK3zk
32s7u/udCfhoUwntU3Xbfrw7H+0+292JGtWXZQKz1p05QWE3jdUUYi7kdopsrrmaFrpayXe4UXx3
zmdzyEEBk4pZ38r0XzIAh+IqACv2rzbSyxS4Y6u2fCDzb0gOT7rpyp2HeXLqR6jpsVHu1f46Ukpr
TIX1k8AmzVk7ghRQI+gY1utus9QHsc3TBzoO9k/T/bz2bsxVYmiuYP/LkAqljIcwtLAL1VVwaY5X
gfOvrKZvMKMS6ESTJ/cUzGJa1uJS9uvzttpnK/So8xnm0o77HLLZzSVEy0KvOv07qFssfLSHOyYG
OZ5Pbm1aesmHJzjsNAxh9Pccoi4p1lBy8vScC6UScU+grTVW4OECiYVym9K45V1ngCz4eAowp50h
/8r30HSvb7KGXa6FHlU9qR/gKQjjKz09+3WljydvQX9hEoX7uIoLJQ6y6RbrBOiDcvjn8lygqKeF
kMDn7OHTa98a+hHA5t6AAhaEKsoTxu3YGSWBzLgHXfO3oXGykiODvRsSGLdufHRo3Uk7JjXhRRtl
yqLTlGUYC9ycs90Zsy35VPlqzmkzf9XI+B3sHznqT2jJkXZbc5VruT95eygXR+S1BKYwD43WrkF7
fYLTULlYHPvHKxFnPgmSTVpr0WOs8h1YFW9/BtDGUF5IlzVko7BP1oExCiHPPTDFyVSvmsCxgkeD
RP7EcqQWcnwcebLDV3dY8VxJcNz9UlFLLQMrZzNlx8LoeZN3aZtWVLdKk02+nXi2anhZGhJJ95K1
t0mCxEvlTVBJX9EAVM7wvakEFtRFtb6vAf63FCvb195J5LU7jbLx48hAQpNGObzMszGzrfuRceqJ
22GP42kD6o4rpCg6J8+mnfAZGOZfPFMrnueC31jzw5xPVaySHAMp9tkkYopGKiABFkFP8cZZKg1u
ppPD3C3q/h0bUU8/cOZaRT7V94+TMAeSq4kxfaHquxMng9oo23/IzgNavlwxtI/qD8Nloc5mizd/
VPIE0Pe9o5ZcrSHoYgpE9YsZeZN+pf7sZmJ1iB6JSn/Dk5VhXwoIcpNBnT8I92mUqfUOPcKVio4R
8xCYPoQES8iY57Gam63jbNVn9M48LuO0CZF96a9WpHAKPkqJsb5wEVClZ/CiJnVrRyC0YqfSi+nZ
cXILe88a7K/uqnHEE+hk/ALBw4sS2eUPsCRvtEWEd7htYBXBdmXUh9HFlKf5zjuK1DDtnl9klml7
+4+D3Xy9qxTn1OG7jhybZvvNBTYjgLY2VkPejAlp1qHKUF1fP+yrEBcQqmc6i4KCOvrbs8axHhkZ
BN1YmoY0Tp+9hNYiALGTbzi49AyOpUpljCj+qMpSOqYKixAL/0pRFfp2egcO8NGvcBDDlfZbo/wD
yhjVyKES2wvgwgjnwKq9gAt9mV1s2f6Z7jSLhU22JOnFh/v5AEP4OeX7HXRrNfU6wRb3hME4I5eS
zgcT6GzbtvHwayFAN7Fx2B5eGf+v/nnzZcMtDO6GxSk58sjj1uO66KdxSXN+DaZYW2pDnLr71n4s
HUM31cSSZC7ltNxoQj96BIQPe9r8UkbF6I+l7BIZtsvhSwiP8ivN1NUori22pqPE2xlC7M9d8hCK
+ZAPaJn7y/pSCD105AiAikH0kNBA4ZldhjlZnhHpDoAPIa7/BG4D8Px5wb+B15pRkwOOJayebJCX
QbtukkdT9Wx2e8vgb1wOe1C6hahECbP2NUesULggY+60lUFVJkyDj3elCCjzvx8Rw78dggJlcKUK
E19vmrT0aSe3Bxs42yZdjLUO+Urf26ISG1lcLf1CADkIggpedQVt/byhAeIvq0VxLq8ErSP/naKX
pI9PYOrTb46ckjeJ7XBz3kAWUVTAVeH1ECUtm0/PnyIEb0zPeviJ6yct0H9rqh0SBVGcbrz7Le6O
Q43MRGd1Fqxbe6QHBegcLfnf663YPr3Skb41Ox7ePZZFFD2AGVuIV7st9U1JExTbw+C2yg/PlmGe
RnsFT4hM94ph2V2885W8eCcVb3CKzTH66W2l53RJrirC7o2Pji08LEbbk2qSZF7ZY8fhdnV+hCBs
2Y0krzoGIuB4jheRSemrajuASbH0lYq7MNBz5Hlj9YKN/28XF2k8gDE4IKUTS3Y0gQT2EbGjWtJ1
qZBxftSeC1z7TL5I06VGzVanGMxXBFn7ebBLgYss9BQHspzWnIEkV2gN/vTy/U/bHff25TNhdR9Y
TIbQs2ZmRfBvKliFcQct7v55CIsbbsBn/TL58iZ5OXGJssXQzC3v/UAGEVUaZ8321fJkyUD+Ty/Y
jeYccIUUz29rrzB5P99rJp78cO2MnWGZ1d/Rwq8SgpiDhUvy8teTFguB3wK2iVsd7fhwGLvt0D86
fl81BSg+KebQScnbBFCfN4pTSyyDfHQ6gZ8sGTFd5ZhOk3JtDYff/hYZo2AZ9i+GJqj273cGvNwJ
4wrgP6/DX0B6TRItxVncJQB9y5NPSDtx4FAiab5TtPfp0jCqr689mZll+LJYwiqTT+EIEFH6g+vN
oqLvtI6FAl+41hTKx+otktgo03SDglmU7MUvcyMOORKmcihCELBcFdW82B0YLvT/OGP/cDtCYICF
WlJW9o6idZd2v+NV8RYVtJOo8s/Z6MU10P/6hPkhBXLFxIsbESp4gThVe2lgLaM5hWIudVBXclu8
l5jForOIeGsgaOwpLOa4Z+l5i04IBopz35ka30VrErny8+IWSI8qKeBFb7ZOSWH+nLulMhKLs4vK
J49edPn24xAEvRnDDhK2Gui4Cnv0MLYQ/H9lyf4qiKy1KFXUjzutsuIDen1CdQooFIgLAfuL/lGg
Ab3DKMpE8I6312JwoqhjJVV4XA4pHPBR6d1dllz4odRqHuja34ixNq0DlnlTqmoZ8QFR0+pohtkN
r0L4Yk3RVEvCt2e21hlpThqVA/sclZJxvFYI9LKuPlm2ZwDcGKOLKhzTK8lyKJVesA/ODMKaFFDI
4FQ703kKCybgzyQ1MZd9oQZgVr2e+9oyxdNeGFNjIv+h0efVM6vOj9niYzBiEbI+ldO3qEmCozZA
3bE+ELYnHPFK/0kx1381rb106Plt1p7HupLX8kQWiapHLJhef4JNE1c76JgUPTVER+Uc/U/sTSH3
CJQHvoQsFW/NSuBvrO9WINvNl6yTjS6EngsW9khRAaiP+hoejoGkf3cJqnZwTLNdWWpFQ7u439Ae
T31NG1srN9jiuBUOoo/g/E1srDA+nkaQcr01Z29uphbnC5ISVH5zTg1rf8Yc/5bMN+bxFExVh6W2
aCM3HbqIMEWh1eeegY2sSBanbPvFvWFBHpen/CCs4uGaJdUZwFGBkMtlx1pzWPdp2hNmgALseeEI
IfZaTBnmJbRLRme97DCHceOa/E0AiQhC7kG5HUYKIEN3MoZVf+0ENC1jBVVu/ofkVnJ3eMO0/AhV
FULtZYwLogtnHEkaTFY3Hz61+2Cm/SPiIA7uM0YZPpnqYwvmv5pEB7BuMYTFCGVMmglxY+EbqaF9
ygqVk5g3lMI7YJ4wS7GZg982xOPWvqCEhRN0DBScuT/qE+df3URb2lv3T7L4r9qdkYNdCmDFzUo7
FA7Eq5p5HgooZhZ0hc6P8VKOTimzAAzhlw1bTvc7p89R2OetLGZHAgXSkM2KDztOV0NESyRqk88L
L6P+Ki3e1fsRjoKXwNTcii9mtEJCqw2/H89JVYDypr6Rpiw3hofHFtwUfNSVY6Zva4+cqbCD/cpB
1YMubg4XRSNXoLi71BJV5nf0kElC5H+I1Qb741jfc6Xfa/rcR+9GjzRKbPLCKadMSY4lWNJs7Fd8
B0nVPCAtctaqFJ9E+8ZF7LDXOj4N6myA7+IIbb4W044O4cuvfl+aD4AokskrhWAZcYOPe6NW4g7M
UXlmNIhOC4vn6aopby3VVlO56xh+X9ARkQBh9fKpX4snMs48+fBN3fOAPU9CO8UAqd+t/dInv+dv
2v9id5STCPruBEtjfKrPvWbvOyyy1XISpk6Tk6FCZf3y04D9JumjO8aJ/+KX++CaodnqOrT6NhuR
jOdHz1S/PAYGRDGOgbWapTiIvqwHIQ8oeMpEyQIyVLDevCwrGOwy8jSZPaqibCOwqxIDg4/kLhCQ
iNnEW2EKUVkqmJEnzrguesEIs03p7uVs+GtoMKLNWNgA6NQMBWmkCe6xPvRe04nhuYYOhY8pNaal
FRfaA0rh3E9RnEZPXfWuvaiPYcHHGhXa8cWny1liOUTBrIbKfOOpTFVBuyHUKDm3rLSkQGQh5Pqn
mkvkA1XY31UZzb3jk7uZEusxzi6Gk4ChyyNAFmJAJoh2fe5W8H1o+YthPyqYb4zuslpqJ7epYP8x
oLb+DM8oX+lZ4UksrTwfrwsHzM7Ntc6vaELfiOgRyUr7CVEJmdPkubmwm5//bbwLcuxeFLx8SuXd
/ER5GxM6sBCUYNtIWGxQa/CvoyeUa1icwDTakvNdo02+k851phuUCXKq1wYF0JvcNSOvcnuSvG4y
3khVv0xyZAPZ+5TYP3H67L24ody0pLa5TxjeYk801xvc58CVOlf9KfdLm5CWskd1eSfm4jZh+Xp4
NZN3OWbGj1sbkgyyCVCp98bvDYOnhTjtFJcJkbN6mOtwhkrln+jXCbI9ymWTSSaXO12DW+0r3EUC
mf5LVToLycDuX/qtbc+CZpY/oU1HZYGTXS3sIMAaooEO6O/gMAJCmgOlDYsVcpt6kLumyDKtIpEO
Sz9mZJiOmcW+pZmm6SBowbjaOILGy8OXwHb/rhnb4k4TiQl8YhG6wcP6Zf5jZ1dgJsnhwl6abnYE
ApA64aQqOGLdwy2RgDBSgYO1JbVtEC8kuvwx4C87Dupev33bPPG2UY/cvT0rlZbuUB9vmgTcMkms
uNM+inrNzf9A1c3T7bCQQhsxZoNJPWxhtG8NEt6FoesL0EXJ0NfaVxJmz5hw4Drjp8aMoJ6NG2ic
CsjfQEFvGnrnXsD6n6WKYWUCBchgm6tNnCECjdhu0p1/WW1uOB7MhVpsqmgn+hrgigb92wg9rO4o
inBQ/7fnRoxDxG+F2S5M5qwyN/aRCCzXQzLw1q24V9Fx0VYHywBNzMs4ehRZkDwgkJPSymQu2NQc
M6y5gDBEFAB1spenNucx7cd6JKWGZjGsJlPGjahALEcg0TfN1rSjngtNL6NgLymstVFqsTDpHfqk
KHZa9dM7YMsUBb/Znu0rORqRMQxIEjzh52J8hAK189prJ+Hn+2rd7ho6LeygGBBxJbTysSAbKoMF
OH5lOFJFUHB7RjFxPfCBvHjWqPUgvlpeYxTNTr0/dkiwDhMS2f5GjmgdN0TIaXUWScOJ+7AIxJY+
+YhBOnsAobQ7DAl6oYY1owd4VtIIKmstuc9n5o4vHJOsHcLhQ/w6qhuvybX+CNUrMKTy1jn+hbKJ
oG33MTyWC46iM8gYJkLMPwWD6qUDTHp0v7QScjBDwliTVST5ZvQLzlfTOtWJ4f4Drngf6Qt2P1Kq
QODhAwqRKQf3FOcY7f8DA0vHw9XN70UXr3mG6MNuVcmqnvdAj/ti2eeHv58xjH/d7A6CBBmdj3u9
ZFoWQcMc/fmr5Zlv2twlBR7cJ9vgUFLYcvwHRyi2aeTuCBvTbVwpLJUpcvdKrUOK1BH+d1ThjXOH
nLpLgErlAHJFV2GuLSCzPbYekqvllD6zufa5zQHVJJ8V5u2lCuLQVFqa41eP8kz6cQ04rObLuOy8
06KIVko+RMR3fY0UEOQdeJAfOB/j/8JHTPlChxmDvt7zJh6HHqzKymNgnKAQ7HuTbk8hphjFEckv
oCJr3L1fVVzYGvqsOeNc5MZy0q5VOc99FcvL/WQJPSSKHCSDXLVFauM8kLYtKDQkKR9E/7LbUUbS
BIeO2pKQfvquirZZYyXXhxUvvBxnXgj9sYQ97yAhtKGFhHMjJaOliiwUVPWJScBK0ihh5E2brbuG
haQDk373ODJ/6CBMTWQ2VpA6KhmgtYMZmjTBqkIMQ+SFFmVIhxqa3bxBST00kuwhwz/GDRZ+PpIK
DHDpon0lLTDvLY7LdDaFQdfPC8bw/0baZ+GTjd5bozL4s6N1xvhwN2BlMK/amt7Z+fhTnjglRYNx
ziGYDMbjBCVEUsCwtbijT1qMHO26PWQt9Lez3xv1qOtFu4RSNxOYDQ37UfE2YeNTTHghUDMo4oAy
e2Jh/s+UuaJygnS5fKLAqHYH2j+nXf2aTg3lnpMqolqMpN4vmG/+/TGg3IJTscYyDpIDYToqyx3Y
6SSXK2Sr9vdc4v/E8NxswzmGilhZRTWaupx+x/+Xn5KM+FAZNgouYxfrtGMyzvEPW/0ymb06bdjQ
eUHK/X2Yq/dMMc6DG/Ur1mTsdr7I96lpef+xX0FX63VXZ8Ctx9FhmyT0Q6qMvE4ssg+kxI3QkzLY
BuIBvTWug5TYF3h7darHSUoMcSjNaTOOwTZ+Wlhxgf6+kCVQgfZnJSPbMI++GnsYwqtOy5Dg6+zV
XT20OFzdhySli26Wbcc5zoBSIrlaiEzOl3jsQyMcY+G5GGoSrHo+6yoT6+svvUng7f/NLQUUp30G
B1Z4B23TP/vwjq/ZQ7WDYIGTNAWzsrpA+0R0Yh4Ggi5pVRkW5NU3q6iUW5Th5FUZQ+QXPPiBSecl
RlSvud69/PYcxpXsyPpq3fGl/ZlDn6WCzWmNTlNJLxKZpTTeRxH/uv4SRy5udZ5wzfGyy205gt74
Sim3MgbtUx+ZBvdWGGMH/pRBtZh7qIT2J40R3PW8HkdymUcOQeYhNtpkiRZc2J3ry2HU3pWGHAgj
T5KRB860jpJ8Ypii9qcoUzde11gFGhX8WktTfZg4J3rR+rltHQ8H2qZHBvVDKvnQJ6n3+72WiHVG
ZBrWzclqz/wTOZJNn+tczTPORdVX3RyGwY84+VDwK4AEg+bcGT/QM65WFHFvhQx4UEaWRJfgJrDH
otSLpdLQ+rDK63xpeoTP4pmRBANP4+H3CNRFm8E7xmwr0CSSIt67X2sD7l3a+0vMPLSFsUmjKijl
4WclzZNJ1dh2sJfZCqNC1o40YMzMVBpHP5E9jLblJkC9yV/oXz5QLMCzOj2o+5s/vq6f5+UatAjL
Te77jtBX+AMapp4WrjAagRql6lrzSsF4W9gRIi/dl8p2R13r0RIcX9LuyrNNb5E+IKQbhCZTqFfX
DPOyZcaLtJq2IKWe62XH26XkY0M32PGXyoM6ECk8JbKYSWAVVo5I8zvlcsV7VVlgFKHUL1JPtJOG
PWRzXh/ZyOi0HQt+qwSy3X9BLj2/m/hSwvRvVZGKI25p/PoZl8ISnucIHP5N0c5bcFlVMb2mPzZP
XmbPgmOwUzp5vWumz/auyYwCjDoIOS6cctxGNJx3Z2wEowHWzvkSC+ZJ5qWOnRKkXr/GGYw1uHcw
I2Y2qeYMPXnJD1fbVXD7IlakXIFLgDK0Y0u6tKf+bAf4pi+C1qFs6bNjXSirj7JD4Ds0Dz2AUpxZ
2mgIj+oKueHV2po2+o/L8dDJihEV4OeDb4qgBJZepDnHTMIeSyyYbhrYBtSk1lqz/rSu6zPOvf6s
3OKE3rj7r3pi1u7VhjxNd+EyEvZH+kHVFMcgXYQxZtsfLVUHYbtqlwI45nbPLPcAvaoQJStisfGN
z4SR8n6jt8PXPYXOHcWQ2FzhXofKcVrrzpT76Fejv6kazJfJ8OP1fLNfITzA2N9RWPL1MrhFu5iy
nWtCshb8blDWYfppG7sJb99x7i39yG8SwX7+TqsszdIow5tYB9d/yrwRyjGpaVe3ro8B7KWTRD/e
OM5a7yVq0prymW4iXScBhqg0iVe/Y4SjRIBioOA99WvgrrsrFOtYEKZhlkrzcPfuMtEAMK80gidp
UwVc4nkpelDHnH9BFYa2WvXhMDyfNlYGabAwzu7t80zyCF1a/gFe1soDCXW2DP0ZERSW9fcTmaXf
SeftVxig4OfIGn3IYlBB7pCEnv5XBaKNVUTD1klFwif5lsoJ1gDeOYeSmXhHcREHu15ggk90//A9
57+mDmmoEevPrDzJpVf5iHZJq+RmedVAaGoZphCSFcEaxyRScAoaI0VE5k2yNjsb7JHP7gBOn48J
nA7/IkplARSzOC4xxs0k+LtLwLNwmepFCHJDqkGZsfntIotvXlMuG8gpQoiPnVqaoihKDoRWeVGt
fUGKiE+nDVUS/j5YPByuivnjN3FWcP6I4N27e0bnQit17rBzvc7LO/4Y1oLX4XV2Aq9ku6E+QOhD
VoMVv+cRwZMNyyd75y+20oJZEu4MLTwQB9F4ZTGRzS5WsEtJ4Rl4L0OiPhuzmwwOg+g1dOimC2jO
GapWbpl4MWYsbGHCfNxNh0FQ6Hv0E61wTHo7+nRBkbuslKJzcffBrnAhYArxMYJnWei3Mp59nPrR
cNlP5I7g10cl9lQCiT1tQVB+PHZ3Epv3pY6yyMpiVrhO4LaTsXOGKZMM3KKe3IrGHQXyX/yNUslG
fF8Id18cVg6aXnYwaJL6bPK+XZxXRngqFadOen4tTIWG2pI0VYAlMNAv7tG/oFhR03oJwIKyF2bR
IVi0HUQh+ifKEneuuZ9/1st8VQLgTVrXUbybywrTYU/64NM7eWzg7cuG162GHfDf3g9HHDnV4KDn
K1XGWbXtFmn8LKp8BhA1v1q+rj7PtmLqhsw+G85QnAuI7Swmo0oi/FFTOlxWfLb3GKbb2zc90nZz
tR+DTyFaHTLUwkd3vPChJgfF4CEuDbAnHJRaAKT0PbOUmUyCqe2QJnQI9eRKarc1rG18PpSsIb2+
QMWk/RYnJtR78fTBaLf/TiNPlQg56OVSoO488rBzBJgQ+fs5qjFTBjoCqmnhZAkJqB3ftsI0vK/l
vXS2VNkO01A48H1fix8pnItz9bmv8gtNUPO/juws9nPOFj3ELbnp3di6m1csQo70eJLwfR4SCi+m
uQkPni/9erQYEIYyKt750vOareZfZyLFQM6RhIqdl4oOdBaugerfYVPe89xOIgzxPDeNAirrtPXk
mMBhmBgse5lHkxiDOQwpoTrpCgZlg4gOmhuHufA8c/9Tz8G8ngMaGTwnUfko3Ymu6FByTIIr0uHD
b8VWOu14bvc5kVR2rNJftG76B7hvziwlusgQFyC//46nKLcQbyaFo74LkYM8kOl9Brel6EYi9RKz
hzSGjixbplp+CgOHac7PMsYAAUGhWfia1SHb9p1HAnYdq0y8KoiU1DyClQnYvROCypIty6eRBfnv
/XkFXGPA7pShaOO+Drdvi3x+0tikANg4gkjt/B3ZjlwNJRqIP/NK619wuJoe9D6vR7/WGaiUYu8v
GgM0N/Sq3H7qKVxBLzlJFVx+O1Kp+0f8Jx2W/4cBcAEtg2AX9HV9lJz8i5ybVGe2m+S1YkS1pSuU
v6SUiE2sC8vrFxA8qPh0SDidhGpED9fTFTr/TCT+TBTYPDv9WqF+mhGYc6LG1L81xJ4tX9od+8Kk
7+Vl3Ycw7FKjn0P79xeGvitNztq5NP8i4Add27vkR4RT45jaSu3k+Uyc5lLJtBCVeUdz2le8oA83
2cVrTntsgwyahR09Y0V6Cx7Qdfn7LvAqRZGSLMLAKz74ymta8i3Ve6iJnjtuOPggWa/vakQbWf2y
MjBb/44muT5pxT6yaN6yTavZVRmZLBLjzz6RlLAzoqr2EOOHcCnKLlwZtiz+cBJq4LpjJayf4MUF
VLEUD7wAfg7eE+w+aPshxsnsobIepGrNZ4/iRz/dJfvEMnfKyAJimbzl3UZoraAbf3FvCNxzoR6L
A0gO1rDABmui7YIGGZTyaNcO1wbf3Bm/pc52BdJSTPdrtedXxohMtWDD2FrpIdWag8Bpprg0xv6t
dVw/MGwkoXYpteEgHenZC2dKcWAU/KAqTmwxEqqP6ZM3DzIbGUlOXNzd3Ih+RU+c0XmwrVAK3RMO
izVXOt/PCeaWOPWZeYZdv5OTFbPYTFXJszC+b/pCLcnylf7oimZYloKDsJL6sD1QzKecx/CW8f1i
sZnRNw4NZiL2UujpSUOJkdwYRE3jtx4C+MdSgR34OJIubdFWmJ6QUHB4VL8DXM24Duvwf/Xp7kOE
W5jbpb4bkaMTMawiw9SHGx7LEnO9gxWgWsWEE9AWphph6dkiBrDGd0lG5fY8Ya5WOz/UanNoigpC
VacL+uRXFZWQp3Jy1sH4xcHcwUfnRANq6QhRni3QiVkzKOPpKaFm6c2QRgLC6QszHb1CIZlTGiGm
0KbzkWtSYmq5p5GMv+xbkQCiGXjTnjojQzuYqVRXYmYB/D4r9x6g60sx5FMRe2WJwzsIJP1dGVQG
kTL0Savc2WlerLTmN9ny2L02C4zSk0kcjx29HNW+4lsb3A6zwPXshWg7RK9/TZXn1IaAj7rUE3AB
uu2zDSWRb0Lud6t552vz8U0zsSVkGLrjSYOIFUCvLGqYx1UVYruLL1YWMGFinNAI/McI1Z8xh6BD
tD8teOkCkepvFi+cU91NdWD/GUJcLhgGCdZgg2TCYZErBgqBQUF41QInmHcVR5s07mmXDwD5qp2Z
UOG0w/MWQ0w29k3nCT4W3OntAaqk2twlU0ZvFej7CgoGAwHI4vHMQBlaPMxQ6lj8bteVbXQnUtBn
EbTtHZQr4J66BIqghURU8hzs/22d9yk1jANuCNluB7L4XInbJAXWXSl6N3YjUziopSLTMRGM8mnF
Uf8C6u33LBzC817ETnPpmn+aDWbAYmh6951kjx8ctEtgK0B/N6uQqTTlTzlds2K1hBVuzJIj/qMu
L7w6r3AHOq4RyrpxJSWBIq/R5/dHcuOy23GvY6cBu/hC7mXSrca51E/OJ5DI3mhHhYcY0FbXNYks
2TPewRHzdu3zZHkWCYfmKE+K7JKngKJfZN9AAciVKTzPu+61CPukOFJpuyfWtRxia9hE/Q33UgLN
GCM2c/Q1+W5UD4AmqZD29mnM56svwVyZjaBPFpMc6H0TGlWlEXOP/mrBx/42GLzByO/y2O9OXbG2
wQhwUCAmsmoJvLesdkEbFGqaBJKeARLwuDC1RavXEgv4tCuZzVni2Zv3xcSaqoXyqDlC3SBGpkHH
4gMw6m0VmPb78q0SLIBJ1O8mWVKHkGLj9PyZvG9T/4UlmHZeHBiuI1WRFnh+cOmVpq4SV8L/DMVO
WXBD5o7NVE2IaaUHpQ0FU3ZSVEzrVRATx2qvtZZbmJsanednEywC92IgKTs/gjhIbu4y5O4mvN14
r5efpULZmqsT1p132YxN2a7HT+6ERUp1xp8AFLcyCgQIAnCEWKivbDjECoyneJzWZ9Jh7+zCer2v
MfGHhmNFTlyesrFX66feLf8pU0QoNEpsLd2xDP32BZ1SI3xfq2hXvREWnmx+S4LqhzFAX4nvap2L
sjeN4lOIxbPCZJ5BlGqSVSPmq2wgmsafryz7Q+UYOgjfdGo1yQ9B/YE/TkWUaphIwmWy7DYW0vky
3tomE00dB+iNdviIqttXMngjEH2aTZ+vJXU8vvkHT4PBFJCCrbZ1VXW+jVFmB2u9Qn+NWxgZcn4p
l+kXeU4KoXPht5FS81orqy9rEvu/evS2/Bt5DZpaMk0R3OzdO+VeImQmSamr1ST9WKP8639qatHg
GgOYdYGN/LJv72FVbBOltyYk5nZWYsoN2pyOgi9k7gViz9ZyT5ppF8y3n1prwBm7fdWpUwuPhUbb
F0TP6EcWayYywzmHic8P4+AJH+6zbr0lOVSQhG6+4hrajfY26hAU8tLKY0iLOZhLFZ3xLXFaV/nQ
RvGLLfV1qX+fyT8fyIW095UdGh0e3A30P0J/8c89PGTKvktYQGVT8z4QH4gmOKGXsdguzSj5KseS
MJInX1n7CDul5ebPjIFWZWHf6Y7vRaGFIbb1Sc+dbN3TXrx5QUAk7Xc9h+jukqSu+/HI2AzpsQ3U
H1QlHH7V8sL/ty2E2XP0V6WSIrR2v3w+bBiqFaKxOVFXJz6OFW5xH00MvhqjXi2Kcc5ssW4lDd2x
q1b76fNtRDAB7LakS/WviY7euCdfUsTIXUD6l2eRbbR7lhhQchGDlZiVhMmY2cmcG+FwVdfKXEhN
pxJxzsG40KQHncrp++K+yQdf1GzfIXFv45VhVXehEHMysw+chQLGHrOntDi+8cACoLxP4YR1iV1A
sXARIn1pEpKltF1PMr390+Xt0x7XzdhXP/ri4nrnjtbMud4jFvHYJILeefWxhgLcnhozJJusQxgC
nWjUqvA4hFkK3cDz9P1b4XkdGhgJC7ctpg6VLFGGs0+iTW08km88YM7M8gBNuQ97tMPHUHS/g106
PoyDhPgZFgZqKbBcvI3TZllRo08+R2QFC05VV8ynIRe7DeZGFyM5ppSGfLetPjNOfWARESEivUHF
W7is3j07Kq29LH80CIIKKpeQjuwsai1urhMah5uOa6gEm0iO+rdhlerGX8fECT/aYZWO5c0z2JMd
Qbehm1vSns5WBMtGl0eKjuijBecwBX0HBdxBzwVruFN148CQnY+sEwrYZh6+zafRX9MCMD0O4FfG
zvgAlPieLDImvQURK5srrg8V9AxhpRoAcg5G4ig/yjQJnIX7NmCWHGry5mQRlLp93H1PHfnCZstM
S/Gp2hHI3S3Vosj03zVv4lm0De2OPt2heQpH3h7+eQihLxtJHYlLpi6dEHLmj0CPZ0kuKvXuY4Vw
zpUe5y0BUNZy7c0OrhVYMz5HCRJGGtZjoyTZxJH46Er/U5MWV9fTfNsfBSZtZ5N/TkSVv2T7+53s
CoNXVZTa2S1swrN+DQszbQ8K8ZLRpwLzVUVH2kHjur1o5FOi/YFUvRX5qk7Xnr2Xj8zcRZgv90oU
Q7qBvPpjilrpYoUmo6awld3D3HAz2EGi4fLDmHGNdHgPOuu++BN8NjGhObM5HTkSrE2F9IXx1+Sp
nxHEhDTg4IbxdtjOTjn4phDZyisHTL+ApyfR4kfoWm4Jaq/YL6n0pnaNNi9OtazrjpQdYAZt1vdo
cO4T6RvJLbZvfPz3oNQgMa4xXmHDZB5f4xI8qi3sEEZgZaBDDo2r7P5gqW0C+2jdEaH4EHb4xA7J
Mvf9REdAowNxaAW1i7/lBhSBVftm1Lv2Ij19cEiAw1qPW/Zb/CSEWLs4VBv3JG6zJgt15d+Zw31O
FSM0yb/boLvJRJk7ZNcRoCeuNHjgSrlxUB6rjgZeVyJOmuhdU4ZaK9x9D+4lzbfxZCeuOCBdhR80
7AevzkUjPGQ9puB6u2J8+0FgCR1Y1ESc02ZhNOiThEJ0rm5awOUjGtvjy3ACspfCCqGcYrIyIYZ4
mUjFJlWOMPEZrjf/aTnzTB9mtzIHa4MZEnmpYAdzcmGtuhipMsA8EFozvCusZPPlvDO7/9g/tyHG
+UC0EcOapy9sskS+/gVG98J1/87biMGeX7tanyAR04rTjKmT6z54Q4haV5C7sawXmaFPpm6kdkp7
eWdFvIfy+gt4h2SNJ0gFw5chAvbMVDw6luj5ymg2WjcxXupQnklI+NA78HTH2heWnsZ5Tixg6tLv
OGViZSlizoHg6xo0p4HY+UJ7p+kt/7GkUEIB3B2JSRr+2kE8grCLaoCN3CMCQVPb2U0E7te0+Z8V
uJCniObXZWqut/k4v2cOevT2BiweoL55jUrqtF/fe1Uf6LjDA7EcZA1U0YzBjPv0qI/L/ppzNmfN
NtfevuPhhjCyWqsqV/y/ibqw6UnxKMi3Y1vjqNJb8W/hiAZ0iZZl+MvEEJqC3DKIn/mEAxkQ6En0
7oZAvGJb7PewitL3kEJstm+NuuIz8Mv58HbC+CEyXBDKQAy7Tc3NTIMZCuoSGO0NHDYCdQhV/iIS
9ql9Su5Bjk+M9vLbJcWxP8wuHDHb1MeS0P42vEzEBrl6Qgdx5v9OnjvgGVo/4m4ZCJHx8epBM2IJ
b24I6f3+5Un9Z7lAKWZYbgJwslrrShWf0opRx3WhnReGsmw+a5G9sI8NCuDlPsGmvHtoFsXZxVRm
7Pl7yVdYjTjTOtpjYlQyhVLewnS+Ozd8SaDIHblWbrXo8r0zplyiph8f6wwZKSl6FVJsJ0Vr4pZI
a//U/wzJV1//dtpD2RuR1lSxgJG1Ode9okJirB20pVGoxXvOluJ43A7c0MTxQDVjHT6Tai6MW8HJ
X00WstAO01WaguYuoJGxrU7rM794v7lrWdcLBYV/ijRrPoow6Sb2NKsZZErGaEVVdaQbDdhuxILA
3WPqZ96YNFW+B6BCyDQsbA++Dh7K58qnB3FoBgIENIfUGZGIZNm+YbeFT4BrDHOVR/bs0C0q/WSw
NTsgK0zf4nMp4HgAVuKkZiPiiqRql/jJvmiurDcGKIpP9GZgUmw9iRxe7lvYhD6/wWv6Ydpn0v3J
g9/gym5C57VDo3hjsN9gdbh9X3Sz+vdXniEpLSeLFPHIVf76A9qGQ2U5nnmVTj6CgB90GxUawXbv
1QfhnXNZiCLF6WvWQdMyDqG8t0lapBuqYPDXOiMvjel8p7g6tAKo5CpyU6GyXRzU2EFgyVxGiPik
NYgBz3QH+huol3R+hD/zDxN9vF/jTVfmqihsmXAjORqDuSWCe4XoldJH5RlEMPObMeg7I8QV2cS7
auXHjktpl2iMXLOiKzLATP8JKioQ5fQwHLLLneT6P22MDniGYrzU6N1KxiXv8+UGpB0pVfeIMi6S
jqKRjILArtJznLlXtCMd0oktKIpgfIhpmWC/+nefgKcUxwMH5KAmPjrnDxhw+eCCsrIrI4fWKbqh
HhtIxN3Zx//Wiaaosfvh/zKy8+3sjPqKjwGnmgi7FpQ3e450cBxlnW4Ic8hf6d+6rJ5jTzgHIitt
WtSt0X/5HGDB1WV3vqcgoFPXmUM1vPGSx9Q4nbTFq5RvlkDUCvX5NYYfXWoiTJY/3Dv8vuS+rrKV
wAvt4seWyU/0ykMGY71SAK8EZe2gT/Vr+VRyOcGnWqtVfRGHbhZOMOFcFX2ZUE5ua95/7pqRzZcf
hJm4BKaDnJ8sWgVP/Zbczyw331NprbYllc9g8K5w2y9otT6lQLE0QRmZXTlI5Eeyh7xAMWrlnIzJ
RbnV3LcdoS5tT7wfsQNzpSytAXkHaHVyPO2wqNuB7fZ05J5qTi7/GUUAhdAPOmX3TfUNjKmbKbC4
xijdlMc0ih0SoiXeTNuVF+xn4gn2dng2RJ69U5IBHRAOKFDAPysWD70euvuaDP1f4TSrefVo9zDN
sWGoUKK1FXhA/lKDjlvjSh16UYWqkKi069j0cNx4ejeRv34u06HuH3RXm/TVTV5nRrFPAjY0sonJ
VCeNRPOvHvTwcCMYMZ4Rg4pAvUFJ9ObzyyLMJjRup4F2ITTHmn0cu5EMc5NAbE2EKb4enn7EkCvD
C6eNaVa6cFXMjbMvbW/snsNH91bCPZMcpbuhmOoiVVxSRCSbeebJf8S5UHqg/v8/xq77m4lDsmVt
OWWdo0Tok55Mbxi8kgdoiLT7v4vTnLe/B7roJZxl6r/8uo5OjQ2JBljDgtYdWKiCDtiXCDgKQjgV
xOQhsP56bnhwlz+NWNZcZb3JH6/JhR96ACVZ0IaWvKkL3M+t8u7pAsH7tqwiOLFE22OpPfNzm4sW
mS+oyGypTheeYrRcQwxFnAS2r8XG++AjNtLS/d2AbaOeNloiTXugcH79skIGrSjHakZ5Wr9Cc8ER
fVdajV1yAATEgA4FXmkquuF6qBzXSOxwwjATiqE9oop4Fl2GFBpNfbBxsFn1qW4OZSVglDp0kaOx
MOCOHXPWWcznsEcDAaQilaCTQxllJ6E3PS/0Bgb08S0f2aQ3GjNGOcPtvi99yfH7ikqZPHskHPJR
7chw/2eaQJydAlW9QZI8YEh4zwxM6SbS6fJveyQIrnGz6ancCm4a+GEjQel6u9XQCCAIfinVTKr8
TCkvGmQXkOVF7vChOKiqmlKqsBFHIc7JfheG2P3ev32Vj45YR4WLO94VPpzayoFu1gB7swjxkdCQ
Mdzqe4Jzsn7UgExngrw+Ae09fsYlHZmvR1Z+aZBPRSibCrvAk3OL2okpV1XUJ1qkmzfAcdxq4BaM
ozjAugZfY2zqiEE2EXHpenz0tMwV6GfEzienAb9xjlKPw9iQT/kWkzB5drmnaru1gOMCksJsNZDJ
ZggwU4mfkUd7r64Qbo1V+2YoYAaj2BiH4zC6V/+89GyBmHp5fuX/1jO0i6iyc0DRGnL0/frNdM1e
Jm2rdoN3QUAVrjQbhWholBowUUH1RHBEfSU19RHO/if8atcW+5tLdz5GbYHAHgwsGQ76H2ZvJS/f
RJs/xpJNJlPwxEv1nv83oSP4liJYQ5fIbOMeF3rWmKwLXEH2vYKc3XWxu0fYuU81Is8aEorQ8UNk
3KPX2k8FFQRwHR6hwLP2Tbcux71a538in1ZbpzKJIO3Z+HMbZgZZFG48pIBaaTQEhu18WsGjFeX0
bdhhkbonuJPkouak7ERC99NboMtpYCNtcpaOlYVcMb4tA875rRwJZ1quwNaZGYUN+5jum8n8l/kd
FZwb1yCRBR6rfBq99OPOhnxyMv5xWeDCyS2yjOG7iUXMC0OCA13ELtSNI5xGIFGW7fV0jw1orAtW
4hk2Vk6XnkYXtyyxNvb07+f0GNUoBHADHMtmVQKdIQCa4SFNYICV+EuSSiXITKybGZaWLPVZTtO9
wcKx9StnNCopFxRk7VT2hkds0Q38YBOgS7L9BHbdi2DwA1cmmlzjSQV+6OwyvQAi/oQ4JNtO1miK
fnumwVyxBAGNEW255oUbwGMi1X8efTugl6rk5/cWofEhizyTnKnRsQxxKVNxDk9hhYSredWW9RA1
GBYz6FxJUQ8xFNmy1AGzFIHrFW5D6FTyfVThYwW0xpQRZSg60GZuH5ywIeg8AxFT7ZuHxY5jyJ1r
7GgR+q4WlcTHE3w4Zboj+aShqTOoK2Vp/lB39JK+ybsldatG+G/3Cgte5MlIHkmeY6DG4+2rIme2
cV1vwD1L6/6W73lqntxl7EhVjXSxpatNPklKHVnpltIhNDkNgX1TuVcpSIvsYQc8PcMubHe+O6iR
LaYxUIDAR0MOlUYeX5t8OUFu+8S6OyjP9Ip0lVxHehGao14WosqJD29NFgDtV3erY//6Vvc+Ee3R
zxza14/B0mStcQOJo7WOCHrYePizJb2MsS/+YoyKwaLYls9N8+W3oEUG9DhSmiSdrB5i05pNKKL2
qJ64HlxpcZMiIgZTqLNMQsv9dahMUY6fU2WbhRroixexdig04iyK6sUfwaEpyjNXE5EplQcozLU1
mqsYEAU/rlutnnOy31vaWM/v9UKD+Y7EMjYfz2NXgpAgEybknmWvE7rBBZJIWle8hsgz/xDiFbFw
IdeoKlkUrurk0oCfZMgm6RE754XeH+2yKA3hSoo9Ir6mJQ4FfyvMkWXAFgQpEYI1gZLR71TtQ0ED
P4i1e8wpuQW7HiRX5YFeAbcCD4HN6qUaSnhW5i7D6BXO90iSgR2NywIBL65d3kmBGCFdZZFF3/KH
01UgJmdPz7pgc3C19n8i19vTDMsMqc5C/Os1reuGJucJBIhWN1xOJQZCdd1wGvKF0uShUXQYoRbp
TGNHdRPMMEGhw3WfMQ/efoGck72Y2dluGlWI7XVVKFyh2nhfBZce9RdIV+sLbVgb/RhZa3rq8wlV
7rElBFn9UshVVs8o1RWy9+isG3Cm+k3TaABg8+rZ7FR1vbzhIu3yWAUbnsgGRoqbdnE2Q7dv3c+f
Tnyf41pKt1myDzYvRjJCJYUTtlDaay+nmoFskQFyeI+vYCr7GPL6aPRpufVS1lYWODT5q9YB2CES
17ul3Luo2KOxMzw5B/9PdNdPHiM7rEtjaAU+yxTmssJ+OCyoqpc0u4zYnqLCno8JL7V2KZfkT+vL
7YQ19GMzQ7o/XStEqUr5N6ESg2I0LNDaEAXrorgZ2jNqdrdkVDV0KSPsqQNYigNRWJ21dRhfKIF2
tgBVIVnGraXhTtiPcer7i+nEvmgFA51EJDTcRchmsn6VzRBJI2GmFmtnx2FF2GM1682gBJ7eSmjs
war+BLMdCh/nu45bpF1ITjeRLbRmC5JBvafYkjh2yIKs8iq/ZTj6ocGRq36xb1DFpU3R4qPIEn1D
KDrp49vykioUgX5tg/YHYGMI7L0oeotPojUsOauOI1XcTGcWxx6LSaGj0gtA2/r2CDQJI2HBjZnV
E10qQ3N2bAKRC/a01hvxzwsGG1HKFkJNaHnIcITP557WybZpy0oCx6XMfi5nOlWXfKNbPDa0hNDa
i1kiLaUtx8nu6N8mADxEfauJ8Z8CvrY0GM+aWLPKKsYzGR6bgeDP28us4iXhZrbpzS0s95wwHinr
0ZKa2sREjLDTymcQ84KXnTqMBNzhZZ+B4Gz6I92roAytOjABS5aud46Hka5wQWn+SOdQWP9LZLDk
lsFBoj6zJdZMxHQEpX7+g2zc/ZjO7v+dNsOm76LA0oovEaZb1+9Oo/Tjeud49Q6yteUQ6frKVdIG
tAqDKj6+aDqFJLJ4dKUTmPAPkQEWsg/KBTmpLpRYvof/Dof197sD7wiaDj++xLp8fr8RcaJV7AyA
Mp5yJyARJfZIgKfEpm8eNBMFA1A26PVNIIGS+bKzWEggfYNHvAXkaBhKnoWEQGWNhu6/Dr07yCXq
0Nzfi4hmaizYumz8Ly5U9twUx7WV8qwPbuZFk+h7BxOplBIBA1EjCs5/ASe/WgkKZAer6+BS2N5P
xvCTlu7/YEPOdGEk7+PY8bVv8ZfVIvYZIiKq3otWqxG4edTz7/3X9DFb/NPyWIkwe4q+sPyFu+GT
4HqQE9o6JR1rM4sUDZQAg4TGKqBNtQkYoAZQW/FFXF0vK6btomZFEwIf/eXH5PocsLTxsWjGlS9H
r/biHxWhbWCpg/5l6U0CrKiGfLpKXnD9+2hQL8L+tv0t4wxw+ZKZesEh1E9jCvPgDzF+3Mp/SX3s
6Knzp41HbQCBNFCsjpIWKJCRpUz5Ox+X2MQKhr5XM/ltT3lbpkOhaY2dgB2Y93MRdFS9I4Yf1Q2X
3kwA2YOv53N2u8P5K84FN91B7dF92Ktn45amsiPyzBvSi+wR5N5VErVpfS1gIkChKNuTey0u2t38
0kUlhrTMQ2Y/iW4bKjyZnugTM8oZUZPowtah37x5Gvn39+9qUPv2HTYhOBOBDYqoo/MeQbmpIQtk
BPyDQvY74+vk2mvfl3yioCxKsZgyg4bCTzZRDAvSXwu6RaF78rqMDfcYS9r2YslouXi0RxLqzz3I
jT2hZMEOXc/lccecI3jGTbGDGr9Ax3bOWDDhQRonhiLzAhth0fcyNzGoSg4Tdr4TOQjaEFolzN7w
md2uHWhxl9SSbjcjHA2m8fnI0s0wUHUEkhozj+FizhyaGTaHl0qgL/4vlh51QoKrla2QoN5+MpyP
3nO1JX/9xsEOXJSbbhRIaNt3UItawHBSZy6MFl5zTaOl/AwrVRg7ZEXPoI/W3Z/AaqapKBOmZJQ4
bH0IJ1lU5ThMiKHWbUtdL+ClrZF+d9jZ3BIEpVaEBph2FmG735kAT6RfZWIK+FcDXyuBCHIgVrCN
enbbVaJKJbsCw5LYF45jDH5opTcYQNUSA/sttYY9rf33C6/8Jq+MvyWeB8Z6Zt67UuS3p+2pT2dy
iNemoojYFRhVJOlTPak8MKP4zG5zEPp2OVKo98e4TQxEuLydGSD0Z0Y7lqFXA7nfHL0TViCL9w65
TfoPSU7kpDR+pj5zMP4u1dGV7xBHL+vhtQqk7P/ZmjnnD3fuQ02vDc1izwk4iKFKeSijRbT4Nus9
mZ/RWzAT2pmGoiGR/DwKUepRJAFpSpIolgBCc9IxN5jS2WFol6kKLA1sxcBvcY2X+6GfPskTbxY5
P02DY+ShEdQJ9itZd+KKbHhc3LDlFiWW+E0yf0AqKV29lnCqepz1YedpUdD1Q2KdahZyMIWqlPPR
cH8MMuNAixbzFyYltS6LYjCxpqmfnk/SVYGq3rqLtGpj8ltJE4PrzuZJkLY3+QHumEhoIeGazyqF
b33l+HfrETKmgeesXdHoT+oD/kfISYr1yLP3o1N0ghlulmXZzAwHvRWueHrQN2vzKmUl5MdfK5Gy
YCrcUHzXcDdcuz2ifdqjfptlAW68szoGyor6d050/SIkhsV7eCnJ/0cFK+cpe2dz5XaOtUxCE+yQ
xhvriN0Qrq+ta1io9M0z+CodB/P9YRZhcDr2+/ByQ7kDOJ83kuk7dOP7lIzBB3pwIMjvp0jIE512
HnMwt4IsxNWJwWvWBUS+iB5ja08N6rViO7vr9SCSZn4aD6+Fd1pD+JoDqOvZQOr36itfuaCy+Y4u
Y0+WfxGrL4hHwjgGx+Oo4NMMjBf9CGEfGCedtHLicr8k2/jl05CU5uX9s7AwPiD/RxQ4CbITMF4Y
9N84xsv8cClyExyAMWrPOEmSs/Cl5n33dTt3pC6YDQ0pXcsCgyYhaj3EMirVS+6EK9HtvV2ocVt0
5Mcjtd23kiiE39+bvPNv3hYlNarSJrNUwjeo4GoMpsJ2y5iFiaglydM+JmWg378onSMXPxFc//ZD
OxkMD1x/cFhd9tcgbEyhjn5bFHPuk3M7plMJ5SULEiUN23BOTCBQd9TcIc/p2l5kB1/zHVHedCNq
Prr1t1wSKQBEGDCzRUyxu2o44XMi/azVCkv22YcKA510CKJEbgkd0p0NQMyr/CEs1TlFMUqTt6x0
3Hg+Sa8BtbfSZr7JVy9QgPP+5i12H3KA2Md41KU3hTh2WClT7GncbNRhr1sSkF3ZEa2SxcAc+xJf
D1xxKiF4eEOCRlL0WX1THk32GGW8r+WfZfOW17mCpuGOZiZQBXG/wMOEFl4y4KqD0SbUILcqAJGJ
9lFWp5iNNSkyS6/MjXUQh+KLoRgBxoBiukNXWPq416tbqemn2w3W9eoJIGP5WesDu2phqTgw8RXc
eWvFSPMe/GxfBmVZuHXfKUipDPzCG+jrWJlsCjCtpccxLM0jGy4dOF7aJX1rpq7Lh3WzJg5PfAua
TFlS+f6uNG1avOfw5uJVBQy+e5VOO0szWOmMBQzIyvYGEdI0eJBRcFAmPeBeglibr5opNZV6QjFt
NqdazxyAQMMJMzSroZFhgXmwNVUqng5ywq4j3Ast5aFN4YvsdQaraGjEwN12/LA3h9iVg9muuREu
vo1GvsF5RJsfdgpK7SC5TPD79tCrp50lHW6Walx5i7h8w/DAN4l1sXgqXXHJnmbKAzdFYvOCyOKV
ME6LNU4MxIpT7WwdQZsfWNeMjMK/al4zvwNMQGQnQ/4VZLJ9P0vwYky/LEV7LfF3hJ7DMMxHaYOa
P0Ddsrto9aw4Fnscrth6I6CHjvpBkcOmM7gd39DM3iiLsFv1ws8nmUK0KqVVjNdY7m6z8J5QpUr5
kV52CwJ516iWpYkurPdwNn83aL1aUXGyxir3IStKoFrYusSsGQEkVi+CQmi9kF+ncPwI8l5pgprt
TtnpD3HGudPJl41SrvGWXo3Zxm0HpcwJVLc94mI4MCCWD2e7Zgp3fdTtWLnzawz1N3PfElYtgUDe
II75JLc46wjIb0bnqcj3dP4X3QYI1XZuQVinwreIcIpjDEUMnMv96BX1PiVT4qmotTWPTCDsh7YM
r0CvDVrjrsose8EY/63KopWyF+AAmyfe/6D54p2JRcAxX56MRLLxInP8dBSCxBO3iSSEwDmqOiW1
4tfjJUxNvd1OL2m3jLDrYG0M8SZOPWED9tEx+8G+0zL+qOO02RonMlA9lTO/ONZFZj4iFnUikSFY
jlW/K+JWbmZbtXcSO2ZxaQfi+gVcSrrfs/DKr/OPCWJYiMfeF9vPTOTBPz8N131PMAd+1MQ5ayh/
mIIan7ZHRDAhW4YMJY3q1han1fIRjeOSPL2/lISlsZEQUMEJVHiXQbNNp6Ek3H6RmiYHFkweZCs0
MdIDuYbMz9EoiumSo/eRc5JASzWl9Do+SEYx6B5Srrnm36A3HIWmEA95A3H/bsUMa8VXLwHhfCxN
jU9WrxzKeoWm4yc6bnXsS/W2X53elz64tP3wjtb9zggEkU8RKBEvWSVl9KpZxUu3iO0fluTqrNdM
pYBiKVaueXpQehDaqXwh3ZOLrANYDe9oed3wBhzvqqryNP/qgAZUt+y1vo6QzLt95RSRZxLKJt92
B6iTRzhGudAesNtbSlyPt7UKGm0sN4pLfQrXZx8Byi00tIScU8T7crw323MK02fpMT3BnZ/kk9ro
lByTZo81cTUXvc8gCt0Tg76PFkZGKIjUIahBIKHPujFDHIMhC6ApkbK19ucVAO9ZpvRU/Om1BOes
nDcQonlVt8v3mX19ZDXfnKsLctyPeilPud8h61fAwa/AYBSR4DfsDnXRd2ngRIQDfTvH9+8ebP3T
ZDsqKkKdCgTCjU62laVyqoeXfkx5m69688YKDbS1k9A8+RwcvMNzMRv+rBv3ypTuK5M3LaFix9ru
L0b12CyxwuSIDjZGlBvL9+Ms6SEsPWYZF/c3nMy7ddJ5aK4/X9JjbwnSoDnkIz06zl0oIqsPCA9v
kZat52iHNOOVXKKvEVpey6XK1dIYvX2uCSuakCm+jefQje8tfxJ4J1dxeyojtWDRm8gbQtKM0GEY
ZGcIYSCfrL4oc122CJTeKkWR5yWrQTabzazP2uIgVEZg669hKj6njG2C02j+AVII1sP5za6CVt15
IyK0oDBOOj2c7JPjBHRFV4vu8jGdLPNC8om9OKbqi71E3XyeIrqSCbkwh6cv4rU7F0A9GYkiHaNY
sqZtPU/rUVEaKWn39ZMR3t5zTH0b/2if+GUARTJcgTjg6gVhUSzkGRlZEnMbrbe/l3At2SH3Bodo
flkGqeCp1zBJhddTRwcv5KTUly52/tbVT136E7gkT+zN5Coi5pFLaWsiBosOIdc1zQdHzs4FTv/J
fw/O65k94zwb5yZU5uInUwiumZrNaFmkoYCTNJWBANUFSII4ETRHPNGXY64Ze+9ZBcyGy5uBqTP+
1LgmgOpnqVSFyRQRlGvfSG7phMl5rIVISUnnqbvoIqOK1pv4VBEyolOycwEI4KIBk/+eogvOzomj
h0hq7F0eKjhpOiVM0UeEpYDABE27gXtlHVMEj0y/HNV2f4Xedk0oG0Aj4EYsudW2UpbYJZCYyIcD
nh5mWT3fu6YCwdNYxcmm1hzqwnYueUobzObjP80ai40uaKjWBjYQt9ndRvOogVF/q0KkjjYGrbu0
fW5sCz3anALB5LyCup1I69s5uGDd0Osk8kvSOVZmfCLJRjHHlXmgufW421Er/yDxpojgMnoXKtY2
IUxbA49/JeWHCAyw5AD26G3hDl9wz34MbkwpMUAqcC0GSqi+dg8sE7dcFZyIOWrR5Mgk0o3F2h8i
wFy09UOOVT2wVisNxU3jcS1IY6N2k96yMiLulU1VnZWpbzvu4xzrl7UkALe/781CXD2OSo02z3ct
P5RNnTpA2ZG39DZjxJ+JnZeoYW+gLviPHI59tc8GdwApLZafJe7pSz5sQTYmuInnTLguWRZ7K9m1
P4e74F0dSOeiAGC8mMtejqoyxiad/23iNpD+ID7VuQJb3OpCiJzFsjMi9n9oAq2wvnUNcDa2SWrv
78eo1HT+eBhvnu2jh4b+f3Ly+hoiH5FeogCvtknkT/ckuXiBsce30auCmRF/gh+34Bhi8E6sGn2D
Qhbviq3BuQYWjCLpa5zJW4Gd3VuLBfazn88sOBqPvzdjIXqwgY/Hl51ULgfdgC1LEuftNhNqUZyZ
pNCUFJKCVRBtxSpqqkBOwpdpr3Tm10qggKGIFvKlfa0PtaE8C0pX4ZmBggb+tsk59xFel+3j8ZmH
TOhQ3ZxzEOSg7oM3AJ7RBQRfrij5KVWiT8sIWXdUZYHV2KRRUzzTGihvzbphcfaC0KCYV4ZXNEy6
wA1kq0VxcvGYR/SNTkpEUjTd85X3kirGOS6iF1bdFnELjMM/O5vu2XG52I2xyVXS28dwdKKvWces
NaP6H/97iZLoyyzqnpeV/197G2/TooTwTtA17TRQOh0YK7yWkYzq/hKWFKD6OvsjzDLylRAY12dC
CG7MiG+MTkGLN0/uCsE3y8z9wGz4eQc+CJKrr3+iFA5KM0+mAd1v5Mm/QMkxkyn8h7C8dfBCoq2a
yogof0K+g1uRoDBtAXM5yrJySpF3wzKMYOocZ2mOp11qpoZ262+QBsFlpY2UlsOrpPWqpBVfI1VN
umStH1saLJgaa8zx//OZ4+HiZXRihD8X2m5YgDeHCVWBSZ4iNVLyAHJ5tIobLfyu4gQIpTl4qijR
rJaGiNw5UYgWmKZT41gF+CFzeiykI97Kv9ccCRUFSNTofDgwZQwURuY5XjvDH475QVi4y3FzVn1r
5elkeoV/EJTFy7/PGs6POFbwZNGtSuazgn9ALqHVeLk20BP7miJtRBkg1d3UIIbDeGOlV+mBJ6ew
3AuiCgW7JVJm5ZdX1sfMAzjHxXDEp/zPj/ynXwV/q0a7kZyk5j6no1u7SFgbZn64qG8NS1V39LZy
ENY22QFtfEr9ctvj+KBm80+iAZ2Oi+C3S0Y3sHMR4aWu2zp9v1vzcBxdoXa7hgIqNgVihEtmF8ct
h0RkEIm/hxStrSabFIedHwB3zzV5g+avxgt6QEF3KA5+ORRVVvEhmo4zYGTje4nHQj419J4vwRFU
RbYurBVr8tP8QEZoYbJMM+FqeYbtjMS96P9Rnr9CqZ+nCp9HNMVVnPwXeY6zQgI9lH49yJuhkgaP
erHflTwR3k38ahoCEAXSrzLMbYJf5f6fV/IDwiohktDxa2AO2IZvqE8h2j0PZmvSvJE57atvQ0Ug
fsGIE51KE+rO5UDJvABCt4IpuNjdcgxhJtfof0HuLjhDqdTInanV/pLz8qm9pdrRO7PkFWi6QA3g
H5Ur78z9w6KrSU2gAn/E2+Twx9Q5sCHJx2jqkIfZyuk8X0jfS6+eioYys/oinO49v/7UpRk1dxzr
PDxjUY4aLFC4co3kdn3PnqlqEwGtwit9wPtnbFDk6/UvAP6Hu3xn1988jJH8OiYerIBLFO+yzlpd
BpQrugEZBV6uMZbRzXVhyExsc0qTEzkvlipCK6pfu29yJokPp2GF6c02sUhe1rAgXzrsatjlvwIU
mXMksVWxWp3OP8kIkXRRMR7cVe0OxsTdZYDz3R+HdRp0pmebDXd1cpvw8PRJEOr+YNZuYotxWIMO
MAw3KaRAWh2LdKUBm5JFpy8NYJxp98Z84A2kGdTSdTCwhuZQQ3GVKx5iBIq7dfW6RA3OOGZzMrrW
+Etf04/YZK4j5c4QbgGqgf+m9zEwPCtznAyKkYFzxLmLgb2NAlmtwq3GkfOEwmdS1YXmQUwVT85X
u5z7/2wNDOV0nuPD4TmoMrNS4oBFnylJfzYo+v9QvkwsBurmSfFZw+TKFJvtI4nYp+tqy3BJilAH
H4hWtOjMhpWZqGMjkzDD7CANJhUkQbvPG2wC2WPPbf/ScTBfLadf9YqT16PtyzhwYLRGuq7jb6DE
hty+ouP+OI5cKGW7RXT9+oNkD9wirutocq6RK8r4YR8f4Rfofbs6lZqZ9XxQeY8DeO/DX6lPmxR7
qIPcj0Sw32aa9ADOY1pCxWS6b0rzutgMeEsTO+knhmxXGYMQ9b+621e1HCMqU5fgXDpgYJ5d6D51
Aloy+oIwzdHaQ1eBCXirdpZBr+Wv8TUfsvM2t2MXxy+zkWmKtf2YCVNbXUiijQxfWYf6G722jxYS
s5MpgCk1MFJ6eoqNZyd5tKo2oCsPRQKHa4rhRYKRKkhsVsj53t55qMigTGDJ665EtlVtz7ujCmce
3XPHjDnLmSScea0vpZi7+GHBi0Sa//Fmrp1odv0GRCnQ0vLfl9WSVEjgt7Upx6UI5JAo4LRNVPTw
U0CvQI4ZVzzY+QyY+GOrgkoicTsFnSxpG9UyjHjiu0jfjelkgUY39znup0Cw1KbHd4XgzTdBrBgw
q91Ww5tY4StwGMJ8ts/O6xGzn0pWWZBFvKFMTxN7upqhDPKkGFLvhqYgtCONousVYr7ExZ0Oux+Q
2Ysv/3T/uY1axGY/lmdBDOM1oWMfxrmcnsvthTG4b+lSU+WoUeWgWGcD+wKm4ZzheQn+abuGhrpI
uSg6K/GCno+BV2PugEtxNn8jvNKf2rgIt3518VbDnBhNZgT2/tYJlHGqsjP5beMWTBzflqqlHfPq
7qK8kIs4c2jN34ZmJXUCc+Cdg9ybSqkJmqUMar+iSX35JosXp1uG8YVHdkA2M7Vn9Ex3YJY5lBbG
yNejhDe9VqsF2M5ErKb7HuaSdUaPn7HMq3gxLwzAyot7H8kBTG0H9SLiD51h/uCiAuZ4bDDhAmhC
yltVgNgpu8uO5zTZobQbLzp64wccNcLg75DQFnyLeK0AsQmD8/hDksvkwvXwyR0Svc8gGyrBIUHk
s/TS9U90ZN77RLdVaoVIXj6xmRBtAtaREA2uhRuAQdLFeJlFLdfGbHsj/apEAsMQWEtwTDcSXoR1
QQp2DImIDOXhB5gubA4UA4eOm4jWO6cAceah1D7jtntrJj2SBYwAHnUrSJ43szW7MFIR/wLCy0wu
nRyqQ/1Ad3ekrQMlnVxx2ej+YgHeevYS1AQ52lHfQiZmMqyE3xozghPiKFxKfBlun/bxjo2Om4lI
A5Nadcf9g+k8mUCcxbWuhlN/9eJRZTD0A/Dd5VPowmd90cgSWxP8meFjLKGEspAzIaWlJYVrvqzr
BazMi/mm5jbXQoNYw2GtLXGGKwg66NUJrAoc84+n13FSK2Td6yEalZQEWEbOSGrv+ASN/LXgCwE6
UyBOA4xqQ81qxCsHLHw0MIvs79fOl5p5NCqbyFJzHhbaUi+lrs7fDT7c79eca28Xn+UeQBxwPDl0
llAw2QW3lZLiwe6kPc0CVtOrgAumqw4VQdkgsKIENxC4n0XiA2hVYKXAwMivatwDJP8Ul5EL3eId
u8WC315FR+5JmREO8bwgjKeDBGYhk521fmt3p505KHTdejwH61Cz619J41IAvjvduFKCX7S6RxP9
UhwgwQB/8q36jv0Ofd82w6L+BVnrPgLbr0IkgTkEBLQQtYr7r+W4URXraaRPgGDIA5pTuGc5yyLl
/oVDcx04NDzoOlDGcicc4JPtXmqHiaNp/VErq1YTP+KfwkqjkoRYTBrzWtRQBVTOasuJlQwCmtoR
p+jmM81oEImWKDup96Du4JNOyHKXd5CNVT0390oo6HsqTlUkMi8jt6tg00RYKqJVs+C0rDkLrrAq
5joUUFLIfGw8oNppYIgELAJLh1Voz1cZXAJ9md4ZII859m9M/SUf9+2sTdV7jKiwqeJlSbVFOCih
y5kWlVU8m3jdajeXAzNriSGABAc7+FFkfAHxLdIs6krW06Y7PmMu2FcZxI748hDWXNVEkJ7/oW64
0659cDRZ653E3CRGBuqUEocvWUIc5LemcoK76lei+X+j0mEhjrNg8YpG3In0hCE2BGkRIn46Dnxt
tO7y7Itvk06vvaowY3sb8UIKErbsZ+4THS09zhFTTEyzoMffRIRmWEGgkwsDwVtbF6KLvzh6T/nu
AXmHIwzEGvc4JUG42duOUWF+28dkyFRRZTBaSo59MVUGjB0ipR7Y63LjT0/KYTbkJWQOuksB3bsF
PrqXA2A0BDb3QNnKlK8oWV37/KNO05qekSL29Zi3Rj2E1jGASYwWBiNVvnre/Y0vbYzmUtaD4vjo
8WwmbqnwR6vpJ3ivAiihf31jB21JjLV5u7qjEu8IcOeON2lSC+6kiOV4U++kHIJxQB1MbWEK4Yh4
55cmeEKNJJjuzQ/JThrt7TSSS/0pdWPJLSzmKGroVWPbQg+t8rImNClA06oxn7J0iF07wTzxEnuu
fTofKmaopwBqHqjuxPyvpTx/5dprdTRyBSidkK5A5UTsDH4M1tOxzbPd5MC2Va/SqjipGotqp8Rt
zhdsJ+J2lx2VXPPDsv981D1LOoiBNAy3A1DW7IsLbzDFCEjR0quCtH/CuUByYrM4hkQw0GmiloFF
+p6p+pknmtVy3H2I7Zb+KmMtt3Sp3MBXbiWXaFOCNZHuO9wsXYjlZeuV4+byEbTMXRnUfVl2fcSY
HUJl+Jfq+J8G5aRknygIuh5dxv7bLjG/DPboRBNS3G49KtxDe2akjAqZducf0CWcm2p7joETl9D1
Ca+00ieXDVXaAITaUzHqKBuMi9njF/Fn1GVSWzbykpfNBoiyGmMqRVy+XMqyDF1GBAbex1cuZc51
plZSLcJL1kTsXhv4Q9wAEZZqvgIKBzS2Yt2ouqEiJIFyzbmw5s0H33bGj+gPLtEtLup3FaGQEfS5
sCcg+cdJFISbWMuezdzRZz1epbkb5cvaUPebAeMOsuKPBLGqhllLxtOapulrqsSWC1dLp/5vkmMw
x8LLf53feDDagq9u04mkKwvdHDN1nnBz2sprq1Zdg8fRk3GFA3SpP/7oxxS36sMtlyaxKcvjr6aO
56NSPTrJHf7v6jg79+JsOggDcJFKPowSl16/yXVO6edXAt/bDf1mk4pFIX9wAHfaHuSOVJFx4/I/
MRHOE1ubPrOzcRJqOzo4igTqP5yFFjfBFUuyJ4OwAscSzAhR7joAn+dfR2vHHhzRwQU4NksJmeF3
yiZ289bLOK7XhUhYZCngdcMWuec2Y7ZRbvAsCcurzRjk0RipX3+eCJW6oTgywQTMQE9jbiOy41r5
XZv1Owy7f2KuV/tzrtAn/ty23vW3F8akWfELzAfQ2l1LRDVUw7Age900U+1Nm/awkCyly+GCDBxA
UrJ6dH7hFopJAC8k+sIpM3iy/RaJbt8RsHlYoiJuHG2aFO0L0ryb/HG0Qef0KIPrvMGDdir+SbsJ
TpfLaV04HhxOxs94RPrRipoBU5iERoOO4zW7vEt2cjKkRnbj91VIiYrciZrNN9W7yIdNzyGVCCaQ
+X/a/CGQKfBkLzjkcujQHMyT/qY0vD9vwTrAkqOR7IcL63pcYzM12CFXGZ6PBYGhFeZLwIeT7nlz
4/fupqxCTP3OXvGIp9vovfa19LUVBQyv2omY/oUNTLqxiA/DWcKyIo5h1BxXdHo7Qtzyt+Jau7fd
AQnI4yHilyC/7q70mERw9KeJHIPsIlBX2ShbZ1JMu8CCKI4yLDp65mkVjzlGTgmzP8FhiOP1fKQm
1huR7BVxqLAwrN6XUQcUMhB7Ih16Sx1zXxLGIB2UW4MVyxBJmxhYoTmJ1Az91VruzJikHs9EUQlP
o0bRR9AuVLJVXCJI9c+bFQqH5kQtvq7dD/nom51b56oKc9KGohXVOCAgwC81fdecJg+rbDuRII/7
ANbbKinamvZhV19Xk84ewn6kB7m87wliqVmYToKua32eoeRP5jkQw1ExkO4QpylOpTVlHMRa/njX
yz2rUX3kOd97TNy9j5DVtsLQwkKLl4UIjQj315VJMSDujebfHl5a2jP7XeeF4BllXRhbnhBBQ5Na
z2HBAu9RYOKOCoQJW4rVPtd3FFVD1DmgaNBr6u9vbaMZbaxwWocstXJRewYzzDiYUZqXZqge7LdY
1FKMBAWk/eRSXdd4jkNSYDvoJ1i4Mft49q9lcrbF1soya/khVcsxdRPIqKmjJMkRLut44w4ul8O2
m034ibPQ+Fk+oKNVIaxp5RH1RWfqf7PQz1AN22kvXe30edIf0MD3WEDdOLC4X7WCntEV/UNDtZGl
Nb8lqU3AYrIT51iIRLkaObJU7M5ASFwDMTGIGZt6y7BdpbrKLW1movYO4cM8tv2AoX/btseaDJFS
ieseKMywavco8bhFI00xm4y2OVDvjprNFzr0BCz8eZUZc3Mn+4QN98D1jpaMHBBAeIRsvloxPQtC
c5+V06xmLBCsgKPS4NPYtkI3QXUJNkIDMQTPZ4q22B24uW61p5FNOEARN9cB/Gnh630cR8S1Tp4g
yfZwZ++cHVx4EK2++3O0EX8Y223rX37edr6aGDHnETCKwsfXECMW0ELQiOVQqsDRoocDFkWgP5S2
fZTAVF51Pc5zp7VaQJafGAVSee3+ajTmodGW8zMZgwAawJm9UgK3TxApYuZLYg8q64azjYySMCGZ
uAkN5ptLIWUckv9RXB21CkBQsyGTV0IjNEQ+Vzro7JO679K+ShwRUyKyZ4X8I8Tr6JKiTqm/oyw5
3BzWyUpm5XGiDRc32pss7FGnPslOScmV6IvjlqY8hVMYFDUEMv0tUMZdDq00lPDh6sj6tmJRkpqC
8+FCjeCQtMafbD8ImQHKbdJ64VYPFz5b3mKDDhLDpPne3rESoY5aG/lzr7NHgObicZHDYF6yYwBU
BayrJmnAT9APPo2ZNroRC7vDqf6Vtiz2tcteAChsbPVqyMkKggT1JZ8jMnzhn7Uiru+15IQ48JNP
4YxQgS8ufLe+F3I145K7XXhSYBH9lFbDvIViAFYoZaSJP0QsC7LDjTQlJmgnN//2FpZBo2Rbyr9Z
LEhwsaynks/qUn7N0rlgzEu9NNyceeDBIuU1Nh8VK629G7bSLVJwBpmjGXWoyyTy0Pb+VyA/GEeF
pHPHmM1DU5jdhk3ltlJ4/V5qk/+TtBz7MGAFKuYm6xPuuAqxg3HNMzagGYge4vY0a+TPuRv4OQ5B
tyWt8aeqWatAgbEvhD7xItftX6CvsNRRKafdMF7VWABBrrtmWs6INuqCb+d/ZtOUE6gNYN1RzrWf
vzQ2kpesbVxwfCjly7qQg/khMnXmMK/3AUSbjy5UGgI3N8GvserwFecL7Dde8Dhwr7gvWxp/nATd
x7DV1M17xvxuXpK91eiIQfVxbjtIclTIHKYtyyu98qB+rINdLxDdaZLm8hw3+QGglgu9XjSCULHN
469HplDfv1Zl4NPYlF3WGPU+J/3AHEpKdX1iJtrviUe84/PxQFe7qA1C9dgVyCfl65whOT0cT4+5
KN4TdT1FLnPSlzDURXYt9q47IpuVW/s8chGQBqLMa45hOFIlkg0tZyRO1uRZEv4K1I3C0C5ODSLk
a8Wj2sZzBOkU/Z35zQwZk/EXznf+8zG/crHBmMcuf75jENFGP/KX52DoPuYyWtMRhTorN4seYQo7
3ZHs6CmARSBLQ3tfDlFUw9oQ8PRTC+GctgvYII2cc3ZgaEFscjwMGXY6BUraXeWVEZHcF6Tf/CxP
3VlXfM9S1ZEWnu9lBuwuoIxOPSDGtjDvvlmJwOurl+xdtt+jhK77EEldFhO8Hy+mYi1h6eH9Wx0X
8+DKqlBYSjyBztRMF4EHyC+4PSG/4obT517zLJB4hSf7hp3KjsktciHf/QGQE1G9NHOPtAl81fgo
gfw30DzAszvPkYghKGqxyXA07kwmii/J9GVQlAuoaTyYwEIrpJIsdUDa7R02+ySSotIwFFF2VNpt
z1awcL9zG2JxU3/Cu/aGyNx0reYZc50VAUdm7f9w+u9pZOKLO1BCkSUBsoOrgWijTCvwdXfGZkOx
p4iDi2CvEduI4V9pEJq7nJtQE1gUSwel1rk3zMsing+zU8MEYc5MMVpb3F/wmOmg37ag/1tnLvEQ
192x+V6B4fPqoDXTFao24a5zr12AH+9PeyJmZpEHHObDdntnyZAbOhdYoC14bEzmuAYyZDUoYOfE
pJxQ1HDnYRETSzaPSpnX8DLxjrMH6rPFKrV7QnuMs9CkaFaSVshxrVXIUuh96y4iGoV+uXMYYR8j
sp+Oqlz12IuGnp3BHZ86UvjbS/RYlblbjtChRJtm+rBMRbjPBs/U2Sc7O7grXBte7ABGqLQdPbLi
9dZ3uoFj2uHaYgCDjOL6InIo8B/cSYaW8gte4MhelA5bBactZO0ij8oDc6vL2onv6XLoHKqUmZ9x
7LqBoz7AOMU9A6x+L1vhmLMcg2blqXteJ4Y+rXo+kkmysK0A2m2oS/oY68cMPeHRoge75r0K9pp1
rRxWZOnBtBp7Ad3w3xCYH0zq3/oP3RalgAS2yaQ17nLbQlp+MJ/WJaK1bhxQXJtIyalU8Y8NSThi
F2bOJzaI9knXAXEcHe8GiDQsI0Wm3R+kgH3PVJMISE8wn3sE8Ql/k4uPZuEWOcv+FDWGqNiJSKhK
GpiJq12+049IvD1ZGq9xPCBPHuO3hSKEkHIUb5VxHvQJ4WzUViyLsQvy0AgFm2wdqBKKyEC4q5Uq
cvXAhmcusZcTd6In/6mntWRDA/dAjjuYQWSBGPdWEnZGIZ5++IBdFl3IVzYKfcSvPaIyr10/TnCV
OiC+Uioop48iEwzHrRMp2cM/O1JDPZJhpipO0cKh04DI1/R3WlFiDyJPLGxSYBGSJt3kDEZDsO8i
5DWqIwpZvd5C5+l5j8Q0mCK+eP8phBkbcic9otMXvxieDxhZ2lb+XfCbAZ7q1T1WzeA375BYNTIo
SplUF6BSiKnslSWCUdji98oKGnAQAtgvb6rLY27/UZhpdr2Y5mtRULZt3JnZTScyKLx3mRLigjJC
L/VydZf/z4O+lIYv3kwgFUHPi428nhfHrGgmnITZRC+uaxCyJX9uKXQMnlSGV0ypBJWSdjYhobUU
oGwaJFOO09B89ebONUlFHCZMuYGO7yC6AHZAjM7jXHzB5Ot8wReP/YSbxyWmJhSwSZPMNm6i0guu
C79ytmDhEL8LmDp3w87WhX+LWFM46pmw5ezDEJzjFofmyJz6YmZhLILEncY2v12TbviCgLjQqIIO
lXB5KK9UrPhNpSpoiHCsKaj262uQe7jYz2/J4pRyg21RVDGuB8OmqgVAFvzTay+F5Cm51+8/OsOg
XsMwD+9yjJZz/fOXFBBVS3vZ3RLFNMc9TJiFuUT66SJTebZ8g5byQjdDbDsnz8hiJFRWfENrFi6S
zpqPDIq7xy/q6eitD1WgwtCB9xprCC9B5E2ulgY4ZGtxdsMZzorVNSMJGb+SdXASnFICxbzgBBw9
itL3WhhkIpHhJrNdSTARBFA1Sp8UGsL73xoKrc4mQm7tFwFqBf64slc3x3ymXUK1NJxMNLLkrBJX
QN12ifGVz7syA6KaYt6R6xZrSRhtb/gV53TKeyY9FbglvoA97CibOahuDGirxT3skCY8Xmla7YWv
EzcLqMpOxJed70gGDbBgGTMrMdYJCH8cNlXhA8EIqMWoE469Sx+sE8537F76mJgVl1V72ZkURADd
Ig1KyNghJu3CMpsITXwoZ0k+nTyYCmX0yLb2MEm3U6FrNEANjTbdwtzAwf8aiaprk69mrQHY1+7R
Gcu2VIRZ/uxQGThBvjbg7L8dRMehdaRDGF308Iwsy8pwssFKKXgCttJ59WlOSh3CnX9P9WLhH6Fa
094Z4vCrMV4n+IgKQigY/uxgRz22OoT9h/1O3kkONdwc5yqla5KyociUT1mxyVcvGT8jZ0c8L9gs
RZS4AWH6bxry3cVAVSS8Z01A0sv0aKw0emJ94VGWDBLRxAXZkXkCywbbCdV981PwD/uG/KmzIMbI
XO8ckBK71/TE1meMrhHNJaFk2Eb8w+izcP+7eR/tToENoUELTbgoOc727TgyecJ5JYtGwjj8a1Kr
TcsV5StQvZ2aFiKFn51thbf07IaI2HINGplIauLituSBHtYZLBg9wvp+VBqugrBw7grC3TrtUsS5
V3YZIalqqV1xGufPvzRPCq+Udqb10fQJpnOTbRy2L04VZN7q1KGNyUs8swpIMf59lIjhTcTQHv0c
sUmk+8i3dGPY6nyFMWsKf25q2BGVm1d8evAG+CgFq7xKYfV68zvH2ghSxHkIIJ+WpDMsF/+tZ14g
8QQsV+kyJ4oi5dCccPUJiSUJqPdqoAjzhOgwV8kYsVnqlMrrwmQORFkJmHHjeIO5JCOBbD3noWWo
SAh2j+Q7WyAvfiwbTYIITUqrxFq5y9gWGNw37d3w7ZsHfcbskGzn2mDcDrV2OW4Tn4H/hf+8tap2
Noi1sUMQgBFe726aHKPaOL9Go2O+C+W8KFJkGAqtN6dPVTuTypULxOMZ0NsGVizObZlwqbSghZye
Nq52fSB88b/wvd7rafm4kxIk+/6bCQizkhRMZB0bktT/lYv0fa37P1U+QNJby8fnCdaswfPCJ1qI
527POBI8zOLqQhkLfIUn0W054ZjxpamGQ7uTETyV3Eq7ff/8gKG2bkHqzgLFE3Z5j5yufLA0MC/F
dvcgkzTmuMz13B2JdxvMEmPWX5LHs0HaxmW0UREE5ALrR0zTGKvmt+O+54+XyE4xsM1qlauo1pXD
HjZsMVXsr/+bPBvZgM3cmeqZREMkJ7qMy3zDqRRiE2TpAt0pWMUbrAkumJCXmPhNg/DFtjZUbMkL
rqy/PhKfVIyAlx1HNgDZ7yBzzHpQaEY047CcA8AcRSQ53b6LFqGipbh/0lLFPPPQbOc9bSv/onLg
Eg2YN12AN/cwPBuSBNRcC7cTdVnKll3VgNjQZelWCZwdC72QxtkEE+TXRUsxSMu8dwTnSRoqZpJs
IgZ+2us0vnHx7/vWkwGs5/y/dIXZ3skgxco5LSy0gFL0Dn53BAlvHmp/LNP3X4nH5lkEyi20kdcr
fn+HjH0otEkx9XiDzIm2CduIy2NGTB3AWzT24mv2ezJPvHTCQaQXpVe8GiwQN1rGCususXNJs3cr
k5J1EpmggWdqMFYorUUxuCb8cWfPHh5fKybCl9jA8bxndu2IrUOt4ovd9oCdkPjXjTxYzURfKuPx
3IldQD3trZzEuKlkHYJgUiteFRHax7tpvpjtjD06YKspXgvAbAOVBuNvu8MD9A7tZVbwY36gRwC6
etfGILFVpCMy9rl7m+2SiBlJrOFq5rKJ5dvMyNz1++Fd3m18iN6Ye8pMs/JsOIHxTovJ6w9nUo1X
BPmdQnl68vTMFLff4LhAZjcyBI8YV8HM0xlb4Q6dUXX/kFphMa2eCXf6RBk1PzeVRkEtBruTHsnq
nlMOrOZbv+8UeW9yeoQDHrc/kB3y72Ga5TND9rIFO5L4HA+FuXuO0VWl+z1RDuPkaSYH6tTeaNNR
cwLPGI3/BmM+hw4GVVSdqk2DdFTz5cwV78FE+ReieH2b6auMUPOIR3WY/9xSqWJ5SXXl+XsfELPI
DcvnZh6bOy/oA5lwLU0XpxuhnjQ0QgSE8cJuAmfIlpCv9ugCpr6nnVCWxhiEN4KnuGccHopTso8c
hLCOkHoj81ryRXqpv5nU9s+1m12YoxIn72gDrftDT4x/4xcGJvkHLM670cJ+M2E1ZAljJhm11fgT
QTOdABPOUG3Y3yRpnRdB5Sve3V1OXu4CaIYpyPKep3Jo8ZtHkfn/ylPF6JGl0s2JELuESfCCBABl
S8Z3GXhajtey+2qs/r2wIYJxh90m28CDqpy2g832bi176ouidN906/AHLUm80u3d/zA8kE+fdelk
Lwm2URwpe8GHRLTdhaoo2IN3GbsKzmM6L9EwhhYWc+6sy2rplQaRR3J/CQ8FT8kISq9F0ujt2t1R
Qxi8zW4X3vkjYhieiQ8YIWi5RDjIZ/9uv1UIEsKVBj2iMzfP/HEA1q0/FhTB9G03t+mfsNKrGyED
R147qhnztESQVlbEq7aOWj5OPcM2agxuJsMh8Fu1C8w1o0e/pMj/N3sOh0uwp0+ozMX0HZmxePwC
bNdpglly+HuRv7Odm372Uzk9HX6eUy1lByue6msfqg8n5nhV8t9ZWtXe/2hTFww5D1F9UBnaZP8K
052cYyAWhoLgf9p00PMCuuqG8yzML1KE2DwmDz5dam+a5CWmnWHEWx/ysMOSmUAmB/NVF+xj6Q6x
049X+cVAK34ifXQ2ImD8fHjLMLEsJPZlh7CUf/4m7fogPpK+FMn9dwxXbREJWiBpONheXqMOGwtA
8ueGZ61jvIF71KGCJxIlbrEiiPoqyGs2tj8bZq2de3d6IMUZkqxkwO6yPAGMbaoTMcjoCPkisfzW
kwCF7UwrGU6lgDvjxvPuzyY1np0HTtq1zduc7CUdgNEsd2hEnOPsl8K3BVvkquTzAeARylxWCZKg
zI5yUyMq5NhbalJbHNSrh5kvtZoxXGZ8GxsKi3Yb/jR9+H/qcGALPUMX/v3Xf+XG2QlL7VRFpVll
Djz734s6LocdIh6VOpgvgh/e7u+4dhiTebGg8nZuXriqCUUmjSzVDwNFS62zODw8LDM7CZyUjtSq
A3M6wV8H9rkyLzLgRh4Q23DsyW4RfZNd1kUMfKs7NlZhTqtqkZdC5/irHz5HegMn1T0YF0miRn0C
xsA2oxVt3WwYaVHzQw8UzTvk6EBinOpgBeal1kc7g8f9iTj6ctDATIBJQfkwdugl0yuSJhj+3Cxj
WEq74GcPlNxdfkZoe5l70G0xrSUP01k0JpDXjANWInibKcHet8aex/56k+Jiug+9A0PCrTNG9JLY
bjroSAilsY7zDApFDo6xzq3Mz4nUbApUVHP6CLiOeD3WA0M3nB3npUinItt5KmLlrNGOpPBxcT6q
ubHWBJu38pYRRvdyG5nY3R4to/t2URi7kqVoO3BhGH7B4Pb0yf5luZVyp8O4RfoQ04mvwC96auM/
TIarjeObs0bR/FJRvVhadYZkbG16ffQA/OToh1jGr0MyfHpdmKuasbkHYrVYlmDUTjm8ybYSdEww
Yx5f6d3pSjzts1IY4Vx7vZSIrKyjP8bya00Og8UgFpO5vf8d+MEpOOuNXXy+Ws49bE/fES9STY2h
nXUENDqPYFmpoFkVtavqgSnDLjd5M1FMjD1tp70fWIEvCZxG8xzRBmdxWuvhQW7owAnAqgefPQ9F
2MuNpokSBCp3QjOBnCKKl+iMqhKgSFBTxPybojvVc9HtK1Nnwq+uDABEAyDJtr2UcBzgoG6a71ku
Fji8b5f17hj4VLtnjyzsyhCh8xRv0BcaJ32CEgIr6PzET3kjdulDtfkrg6UJs7yAGK2BjQSeTKgb
LtbiGSuBhsqeXLIejh3qfIMl/zCOU6CncZN+Qwcy0q0ru1fIIM8TbEi2Q/tWGKlzl58tsWttdx6Y
//8IAiTCSuJ87380v6O3m/VxZesKywIjYawtYVtfCpdzjrFlwacuNensQrFRbJ6pJSC3YRv+iiBN
Sj/og0jS2faOgdnjDT8WF8LBOpHczoaSoRMFfwCYO0a4LzXOwPhTcLKqOoaHlOsWUT23GQlbPTL2
O+ATzLkSsuOYhxYDxwiqfPFdcUdZgG8J34anEwc+pE3B/2oKqL9WYFB7DeDszvNLYcqRzcaMmMu5
RrLJwCXMdDOqEgPQz8YHkOaVQzVYmjLLpyKOpAnJZYKYBnPfTp9T0psZKbFhYZsSReCIofWizQ1z
mMVvkh9NNWAEDxWIMXzEeHXLS2GtTfN1cPYs+c949TkOMowAgopEkW02Kgw98lC8P2X2han+42kv
oF+mzwBR13YopLy2A7s2DzByWvZ3y2ViURsGafyTC4uEweoR256vNCEq7y3tcRsY4Gpofvjw0AsR
WXy5Q9Kc+ouRC4w06RZJ1qShUOgiy7vv9gTGR6gVzki46FNC9rGM/6gE/zLBgGRLzl8SGQ5svXkv
FMbvOtNjbm1ggYrbWHX6JUWJ4DaMRlFDP1qfpWHF+jcaxE/9H1z2nCVwB56NDOfZGhk2o+IZSSbk
ObpEiA9k5Uzt/5rS0A4Le8Sg2ycqJmQs4B8o0b4KtEoWSduKxE8Q7g4zF91yn2TGdJjKb2nkkizk
srcx6ewjEcE9n/RyGlRMMzyy47WQlKq1MLi6r6JXDYT0QSYiY5J4LS0F+UzAUYD/XrlW3XQRls4O
buLfTjZIdtJQSGGKVtF82dXpwH6d9ahpoux3R50eO+E2w9QS4UIvJblyc8eDDpMEBBi0DzWAkI4Z
TsXFmYxY5wcXZ5m+dX6ii6hxFbm5aHPyWneP5MRk/fVJ+gd7IpNGG6sts+ifoU6sF+EhqOz4rRXO
OH6NgpHrs0TNM+9HP0qc440/6gujz70u50t4VBTJHRbjkokZbUi2rrzfMRtBZGnzicVvBXGm1tVs
xLj5Za197KTMIeH9QHTo1Fm5X3E7Pw/XZpeuLpNGCLnxBVVZh/myjkGiRZGxJkgHi7dXyiMoHgbl
euhO8HqB5jA5U7yP9Fbcg/h+MbjDP8F52o7VEkvaABI4nj0345Oc1Kl5Cx9/WGQ6rj2dXGEaDrJ0
EG98S9YPWU29uSY13I76wfaypL4B2YdooeqQJSB9zHk8XPTYwkVblCKbBzKnTPMb3dY3sdreOTRh
dgvfxb8HtsRUB7rIzUmGcR4p7p5wpd54BgtauBl2eBwqUkP2srN8xYexpOZDsmxfktBIT2ViYKs1
UuGf+8Bhr7zdMfStn//F/MfYOeoHm01s47FaG75EeEeVZy3ZHIHEOvx/PTv170n1lKtMEWHFFrJY
7R0XS3vNW5RRUhY1XnRqH/csZnIdcpbzCd63uKmj6rVlq4z4CEq2Uw/hxbNTTdEjP64Xihh5ovPx
GnZOUQ+wc3zQBVVkLGSzwT7jPDrAFcPgdAG/1wFfGGARmPBAdIgkd34N0rHRG/Pvg6iDOGTPWyWw
N5IZWr/bvwN4XwtbmOlpidoor2+X/ExRiIumhLnF/xCL8LV29s75fbYR+8epZ//3U/CxepK8bMXm
sixMtsP9fcnDUNwNMTfaaNmi8a7KZRqJHZNu8l3yT8FbO9Gq6iSEZam8rvLBHoy/G8s2v0EAXG+p
0zvgtQCKqfKzjo8oBrwBSs9mmLmyOlQ+ZlKnY0Pdg78NUc1o3Pp+UbXCdhrgPiYqTUoK/SD4OxBh
DuWqJnMBlwmLLT1BcVWqPPW/TARzJAydY60W4vV82pG924A5T97wxuRl+y+mjmwbg4S7ERP7NdCc
+1SYaNg3hTG4SiEAeQOuyLtBQ+bZvYvAShszmFWrtu91uPX0ymwujDR1gatlwnEhPYwe88RdDLbB
7a7scoVuXPTN9xVSMZGmCu750fMdsOP8787j8Xr/qLvyXZT3QJhWqJlvoIDn53sDSOksKbZ7m0Ge
grmTwdx5ijsxP7QPGc5QDRvCgeH1+cF+0SDt7VliYeSzItG5u6HpGpPL3P/K9iZLi0xUZkWJ7d8L
ZMPOAVe+8BFUNV8rdiFM57yiG7rFSzFBQ1x5LK1phN1QpkqhSqmbR1oaChsxRN1UnoMly1yP7x6l
exijFS2Sg06pocjHngOiU1hg8kyKA7LFW6LG6O0vDHw3tePxr5po1fR7nsR3TkSquHlWLjuD75LG
HLCMwjLY9/N/afTko7gzYQ9aOsBfGzREL1Szhluob3aWchUaCaoPsnfykm8bXOVLIBUl0Yd+ja74
wjZIPyRIqSSN7hHfBC3itS52reAfYM/gIY5jq55ax6EbGrNz4/UQc77UOc+YPkv1CbDqsjMtB6V+
lmwKMKsU0TFumVyQJPiw+KySUv6FLCfKIOWwKUiEMCi7Hh293vXoHgxVs4Jdn0WVCum9c4iJ4C7U
K9Tu1kbG9TeF1jsFnUtsfhs3yKKtD/6UWHHFkHDnPI8tt06S3GLVDKcCydxOuGO7siV5vmYmi6NM
Mkbwtj24cNvzl7H/4sV3TMZzmYzvpEUTvDz5CRKCnAvAYfs423Y+1QgucSqliB62MjhtdYDZJK7Y
mSPVLngOV/jA3TBPgQ9P8/wvYbzu/911Ve/FhBpfUwjxzdiRx0W4wHMZnEfLyOgdA6Qlkau/Oews
3xGM20mxSe1DwKPPHYqfzsOsTJXEq2gGDKYGXoHfsD6VCi5r3oONmM0zS5+vfIamRIlx+UAYOkJr
4ShlL98Bg067O63Qkw2xzuNqpQ+6ZrJFOCUsJ8pwCQ0t9k6u6PUA9QbOdTno/RJ5FlXotPhX0YY2
TSHUxKt+xKsjX0kOq+N1AGbkTQnWl8O744jvYwoH1J4hNFy3xm3lqQnYyb9i+g6ua6nhFah8ilBJ
CatqMsf9t6dkW0TFD+yuEBXdg4QfOmdmah5Ph8dLtTxy9hPZdQOQ4bCb88brN6WCkvCkcqaxFdbD
K+b+LmENJqfDopzNTZ14u3+By/0x3G5lAGNxXy/Z6gGcnxggQFaa8aaYMqYAY01AZSQamDIGjSKy
Yie6DS9ckqvz8HPngzG3oiG/4pU7rJVn+ujnEUnsvh7mYE5Qw2TC8+xVOd0KJ0laTPdqRaNZ8GdJ
/W9GMCL1OXtXTw4Qm5csYntZlJUwSSlEAAX8MIhW3KYFXfxKL8iAL/cKr+12I3t/1EMccCZjTbtF
yonahdBBU8OPXNpD2oqwYC6D0lvIO+tUmryU9rZL6zwbJwKb3HxtEg3Aw4tmuTBaND+roAa4tSMZ
C9JOAsuVtv9qc79QPbDyEJnScq5QPlem1y5Gxdc5qEU7iCyRp+fMh9OrYTAaZ0bONlSAhpC1p7OT
CUhEgJdNuH46lC6WtQLcqwPVGAx1AGdX4OmHdmGyuknKFabPcMmHfBtPst0rKozI1lwB6ZTDLVBQ
ivg5Cn4FW5Ck1C2xvMBzCfhXvuJJ1A7oDD+vPWzAC7CICY1wzh5JqPW+dYqjZaFYkWNQ4Qg9eZCA
FHC0deySjzEg16MQ7+O/Xfi+lfQGK9I/sO4ugl7EpG265Y/A8GGciLyrlXuLYocboWCgBXiTgh2w
2reL2IXg86gBZvvdB6t9X2rYt9RSc8u779fDn9Pl/5+TdwKyITfbuWnDDVIh0e9+06G2LWY1JJXm
riOvnlefTcfOffBfTV7NvGnvP93bBd0GfI8xKfK4JtktL8mjj3JbBz/trkEUmOM2qmZqAxRcd6WL
/hpWK7VR0KeYHe+5Ifab+T6E5GZT3eSAcEJIiGQhf6sBPpHJ8lPlXkISxlLYDvc9qzqFcxu6Xnsw
hcGMZqQKWd1eGdhze6nXWZT0YPq/DUYS8Cj3pTv1bderthswONp/lK/NLyQIx70RaPylWdgfcK9M
Z37+ZizZNgTkdBCiX3vQYhhcGogut9gLStkfwbfozx65WZ+16uAJPyYOrO9Usj/k9da/GRkb1H7c
WvmbPmufW0kWtgZRCnhpAhYKIgwfHnWw7djfQWB2B0C2kplF4h86JTyzF9fyUn4fpwJFqQy3T9jS
lv379ZTa6kfvE3mgkvLSfQRIgcxvS+Wj4iN9El4IMhNUzN0qdZQk2Y5WjpVtj9njFrn4GhQipzOp
ES8oQgD+5O7sz+silJJSP7ZQG+0r/CLoos2O2JA/+xI/bqYgNAbQmHbV9MdVSrCeANi2zGBiXxmb
+t4M6r1AnWS+DI2MLG6bGhkPiq7SPzeHHdjHiR8yNyRsQqJCP6fA2+VsTmL5PCguvdtKBH4lhdwf
qgyg/z8FtF+W4MsvQ/VI4xPoQZ3peCCiUpvRhCnuVHzC2dE794PJMkkl8yMP7+vwnYhzno9RvLRI
QCMD+nVqIAIZfUfLtC1tbuoq6wm9P0hT7OhHQDzzyYv8x4D8NYD38e3kNFJYYV9/9ayUO2oX/z/k
LpJMF+fCQYxxBvQKMlXzxy4tsxTyqVOdUy9CyN95DbTtnwth3dHICKuRJXXH5qPpRzI77cLCRthV
nL6jzk9g3EPJErRpNNgsg6fWQ4XV/M4eF4yqgXdzRd2KIBB1Ck40wuopX7vkv8v5ECA3M90qx/44
tg6TWrhcuJkP4Qs/alf6bQn0S+eVMbS7lGuPEXTVPmW0UiY9hH+uVuYJt8n9SOFPJT3Kq5agpdJN
903wMTsSjsIZE4T7ygClvmyv64yvcNOsm7rlwrZdFH0gF5ZG2QRA/iNb6k42vCaw28gnyVSO1p5K
717sTPIMENpvJs0gtJkbiXNgrip0Lgr9r2cDIH7BtTfJ82AqoF0um27Lk2j//G1SaJZ7s3oL5dHr
CgCJZ/rTwcU0H6On94zL8OEDpX61rsyXMdd7VXhOmC8/FHuid1CNfn14KsIna0SqTxwyGBSF8Q6l
N8M2C+K+UQc540fpcKhmlMBbRAPq5cOLS8UBl7lx7j4XnuNEX1Y/bluFq7lJCbVVWii+S9t3KwpY
HrMX48QcIvb/Hp9YBOuXEOo17Ar2SMWkmqR9ZxpFTM59ZMrwUY1ee1/NpWycl7A03KVgaxuAtAj5
9DyWY7aOiOf2gH3Yo7CZiAhJWB8bqXkD3+xu560RBtTXyqRD6OSqN6nv0iE9n3jV5GRtXKOYF1m9
5glxW9XrCEnmSCjnkL6Q7t+cYGmrEcKHJYY0+UQyVKqwSkgk4/qpGoG1tlrwk6Lzrah0mUL1UAy+
k7mGbDlmHxbkgm2M2hxbwZ7WrmoE5nDBGMTOF2LSeT8oj4Qrg0srANJZfkDXc4wvz72csy1IIDEt
yUwKSwfwJALC76YS9L3eqtQxNZqDKJUkdhjU5wEsKrLvFc8C3IrybkBunbZpOARSfnasxlYCjsgn
66UvLnhqQjejlbGTV4GzvSgi6xjt7HlYzH7KhR+tIsIVjA9meYPEKXjL/BrlicW2mDEqRxd8K1Fd
Nw5CGX7OTPFjNKa2itWZbmTfLmMqiTEIuHmxwMau/bHeOVu7qhTsC++CI+1jQ2vWb2dgz9f5lyp8
3bQbzBLjtYGzK0NTDkB1eG6rQ0v2h2egqt/qLjYErhyUYq3BGkbG1eEqtL3u31b5lRnd3r5fz2t0
NrT1HZKgKSD24wtUcvn4ngaWHPF8X+1fePxouy0lzRXLv7qx1/FnjwtER4l0toIf6tIwTchllRqg
FswtoJLV0Ddj/4O3qpabF6pd1oEYdCaJxI8IP+D+jR28V2uVwA7VnH3SM+oFvDQg3TcZPmAdgLme
2x3tvjG4W9vMfRxGuQO3i6AGRHRzsUp6zkC0ZxWOQ6xCwrTFwNJ+mEFf4YF5DAEgOFYxHDEl+05S
IEvO4Dox+t3V60lRc4vc7RjDWw6laS6zG151bKklOPVndNX7HKn6o9IOQkZ0AsRaJfsVR8GMbwH4
KW3kpPv6VTsGCDtAKNJKR4ZsaTgqvNIMfW1jlOuxjTYLidWH3/YZW8TtFJn957pK5SXqBd7I8w0H
KJlO1ahc9jIOlLIgx91uQyDxgFDQ4qUeqhUbgEx/HekkvZtdNJHKdM1a+zwBtNC2zwTrBbWtqQ5B
5Gekn4RXGHcFU9qx+Q8eIpJBNXK+5vAiyWaeHmJZ5xLgK7xiKFGtHrjUcqgwdyYhPpW/mrbt1VP/
Du3sMOCSrnUOTHnVi3Yp3/G8UkJm515s2ITgy0WELVoS47lc46yMWexk1RGnK0c12nQSKTNZmFYt
rlAvUkt4VgwzBFhCPxu5iOvTY6FKYKrzRUUeB70whTRGW50pmiF7DJeeyVjLqFvD3p3yx+V6CyZx
mKrqsu9qcPdgYryCk0D0Vk8yO6eFj2QCvfwAVq62LSIYKrRc1IQMfViKi4wxS+syDJyA1nihmE9U
VWg/Q/iMWX3sytkZ5E5U2WD3ptY7BcbGCna30M4LCLiBLgfp+v49Ekv4no6df6cuXniHr4KbNT3P
Mp2o1nFTHDvOjU/ft1F5xBfNE8FAQtRjcS8MIwEKXPt5jyMgz1JAwbhetdITNWAiOOBX+KZXGsmC
iYlkpGAtMI8yqd1IiB9xhwu6ITs4FR6akMfw627tK/rWopHdCFmTluNPH+/HHByDPK9FG5EoSfQy
7t1oVvLEzGDeniJQd9G/CBA7GJkJJo7rp9WDeo6OZ9Mwz2g381SgDYeDFWxJmZ1W8pOYs1LZ4opf
ou6u0T8bqs4xkmcWQZkAtsXbSxmdiArhtxXETfK6/0/2H9dvcbr9jxoBmZmst+SoStG5rL3No/Op
J0kRvmsN7iKf+PVHZweRbiWZW9B8pFcABYPKDSkDSwlV4MkNCyKNFtgCgLSefjlw0C7cxskPraht
vDe6x5/OUT1nSrrJdUEf7O3XQHFCgW0FU/ubeARhJOaYrGqRl338IX8UppehOGC7eSMYZ6jRVdG7
HzU9B8pIz3iJ+tS2uzzTljUpESP4uQ5dhl4xF3aBH8LCiAI6a37/EHvmQp7Zr0ZAyYlhX16BFk0P
XpnByI/xFmLasRePX3f681tEJvE3ujS4H2O/UcWNBTdkXBclmu7j9AvN4j39L2aXyWzPNchxBwMb
eaw9/zBTh9nP5pWG0QWpsPGBrAv6L4d22YKV2c6pQPNGKZ3tkta5/1IAbAWJSm63vf7NvAtI1VnP
2AZFfp7wPfu2+jaW4OWcKZCO8MHr2pTCLaab5fqspDe5ZPtoR+TctUKsSbJ0PX9kbZ2s+QIOSTw8
raCmpmUMx759UgKR6EXC9JzvdyK7xodIVbGqeCB9PoW+3WF/tbvBt5Y3UlkCkJfL16XJdamI8avh
Dt0XYLSsk67ljc3vc6cT+Ylq95qQD11Bvk52hgZX3ihD58DeEWgds/0Rd+Uz3RAjFdatdPx958vD
xNPV9kC0si792JJ/kv2ACNAx1udLZ1CW628gGswTELRACA4+P3JiM8EO5Czy4II8gtSMDYVj9/fX
pCxP3G8c4OzKMQzrzUGp3PfBLVMQfMT1GFYUWwTPuI2uhRc9cyRMpNA8yvHvFCO75U6w2M5kkccr
P1d5VdjwNwOZ7f6nHT8DzVN3BDnchaLPFeShloxEQOY5+jeTFcrT876AGZwE2caT1ELpaGi7r1mM
VXlZ3vpEJi64dnyAc0SqwZXYkbMs41cwj+fsAgZktS7nEGow3WD3d0NZ3KOuDhmdZzsfDd3XeYo6
q5uwVP8/Xjs+TxksCtIA5aRWfLz8U6XcLcni4NA8bTCgDsuhdeNSziMIsuEW6yWs2lchNU7kjaLp
/h2ybel5pUusj5WAHIqufCMnLkbjHgTzz7l62NkeaqLlDwmUbHPyaLwna6z7V4KotAPnygmE6QRg
e43yOjDdgYezNDgvPivvTO22MFxb4RgrIgHEvCaFOaSn8fC5gunu9/YqN/QJl9wrk9NQkdHG3nks
XORpmbpMtmsnilIiV7c4+eSO62xxKnPnIkmU+VMyXzagGI0Fd2TAtBIVdqEZdgUmMpiIbHyeznMk
lYrWayvndsWchSuTugPxp5qW0hwOvH0gyV+3FIHW6WkNv53Jwc4k+tx5L47yOO9wgg7rpSVf6C9+
cOPxsvS3Ud3UbbO+lCmUuaJtSY4MxJOXA0oAhTFcfJv51vFELUU0uiMzEdCsIZU/n/SmV1pRGMtw
OYRGJGlRIw6geEe0tkNBIO5bW21yJ8CMJHmAGdwbcWcXMZycTloklUj6HNIPxYA8ki1+C78ytuUE
zJ/XslhwLzOUVcu6gmspFkDdQN1smNkzFW8DWW4NOrpwG7g0RuPOXoZczy8P3St7x5YRGyUy/lJX
1GRMjGwgSSOIDe2tQXfcFLq1Hp0WuusdI7MJyW+K0ctXd636ubIiIeUxP9I7x9ezws1K1pQyda2q
XGGmjOFWckT8hDfDR/vJIxk+VM1vxY4O6+8QRxSXcdTD3IhPJgxRaQ2hWpTqkMQDduh8mBtAPEFp
aRSEAOLONWAP9vcOjPAHE7Iq4xmRwGOLFIfcRfrsy7jjCBVGSTMqKKPNAj0QOnbpuBFSu+RFCofc
SU/n6HdLGlSvrVxeA7hzRgnqNQeEDxR+8Er/60Sw4YuF4L7LYJbDm90wXtuywQO3WVtVXgLOhixc
bC/QdhC7i0k79sowNdEZMiDtIi4ja4KlH9AdkUwHWzvq6yZVEXtg+uND/t0qFrBlt5LMqRdrMtVH
6rSrJnRQRTKzjh1R4Wjqsf4wvT/HndZiaxmeQGjhPCQj5c+7KJFSn+Ntpm/YAdZP85aBXOMHhwd3
GoQw7iCLB4q+39LDDmNi711be3aGiLLyGCKXBQG9Zfpq7zKJwI8NKwRrp3tpttzPj/ddmmNeGg8B
q8y6BVyeYCEj8D3dtu1VE0nA9zJPh9HE9yhJ5MGyVWs62Qf2Noe3v7i07evF7MTdAPY2ELA1fORg
2wgD+ax49wxJ1zk8NlawNRuEHOFVGIh0f8y/GUBY24cM3stWiPMm4Hvqv6kKMzVmZL9gLIHr2nM+
wexFNnCJIkHDiOedsuUwe/J7Z5FPY2PT/qGB/Dgoce5Tw1mKsCsH3jJXjWSi/1uCe17mWsRpNCMd
qI/H2eop6VhEQtpqY6J+N8UCLgvP2Rhvgd/mkjDoPUySQszwaHw73zI0CVKwMTBT5vHbscP9oJRi
r4aPGzmiJzGq9RyCUr4w+uM0R6xMHkBdpvbQxfXiRqgFLhLbMcnnM6FAc0uZfyUKrsyVWNGHdkqa
z28oDFlUQ+vvj9SLIP6cyNyRn+pgYFjuNln3Ng7by9DMjySQ1NBAt1bWycyHU/3hm+hDlt4Z1JFD
QzTtXRRiKs9Ss8r7OjAf19UDZ+B1uiJpnM5BvK5HVRTHGRQmtiXXjuUciqwOwbujxUDY+/IIIXc/
q0i+VHO3bi/VTMCKq6F3Dm1H8lMScG+JQpxyT+QUJsQMCWyHCHlek/8qzIkRRiI+DzpI2cO2jUGI
AccXHwVWDGa1eQgERPOtgtRA9S/lJFoJyNyJ3yGPgsqM6v1o+JFlKLX5OfvHPDyr+2L9nJ5oWYVk
unjErpUAVe6590nHIdc00XtIQi4eY3bMuColjIYU0iHqIB4LUiGEQdBF/1aUt+Qxu9tNyhtXpIWC
Omzft1RvfFi6MCzdt0yVlm2KULyXb9TH3+bBtZWqt5X8qEBP6dDrIHnTvQNLUAuooXZ+cdZTdRnS
kShJAyBjuL9NZNglRYVWj2Sb8v44kbcwUHDIKzZE+sj8+jTDoqX/VTDxruNy6SmtPM+Ji/VkS8kd
N39iwqrvo2HZINONG/sCOVTvYYk6QB1BYy1PaoOZEg8pCOssS246JUeU2Fx3PwEUokx8JNg+d/nd
umLGVZcthyRUfmbIEQ7aMR651EDVMe7foXOF3ZgSiFKtvqXKtRmXawhYrvKD6BY2apcCpNrxRJjI
ciDa/bzJ7VtUKBwJox79q7dcT8oYKxvvR+zSB/J/pAL0MwRgGhzfiE16DAia/QJiJFggZ8GNBjy1
zBQpn2tyNqATSIZtQ4paxhunVCWCIOri5DL/arbNgc3dxHrpX706utF88FfChRvJNB6WoSiN5Ijr
rhSFZt2rX9jGsk9uFyjbhAgpVeYD82pkB654SmBPPyCtBNuqWvwx1+Ixt+wUSLX91VJLZ8I3aeJd
wtTO0vBYA3JYP6UK+1wkKmqJgtRLx1rTuCvqT1sew8beXDjzEQ5T/YdyrJUGyUh6WSj7tOI7aNlR
yOCh7QwIOsmeVUcGje26eQJkmTErG3jKQHdVgnzKMTx3RYeZJNabbk6qAQ9/2yuIHWmSKZ8Xc9mK
LyXhXExGtIpdE2awysJRH9+toZbrywLrXz5y/qmzkslTrd6AutAVMRgshCrGjvMn95krMGBDUPJW
q2ED7stWnSZrYbZFsSc3hJteaKrX2yyAVQ4rXT3yPrHmmCit5fto6z7PEixYBCQwSFKJYZBdyH2T
NJi818y6n3gJ+mE+YFGz61GPhIYg/vfb6NTxYIFABU0MWcP+BTO8Mr41ZmWfIGlEEpc7VkDwGN8u
dVrBVN2bJk3FqpTsIEsyvVOmoOnKtSTyZVJSkUIbpOABxbH3te5jqW+T/Lx5WgR4mfLHAHE9BO1r
ZDZzHXLr8wHQI3IQL9Lk5OLaA1xQLkmdkNVclMmoLf327AGgz0vKpe8ZTRJh0uOQYf1O+12dR+yv
2cHBSUbm8wTYYbNv1e5GDRtioqEi7xxVL85QgkhjAfIAayAdzvZlXA4JI2aNEEXwvoH2Uc2T+GY9
jrktyX48q4qTfmpq1L5ltVqQtaxGZCPkxVFSTtoKatfTmhbKPZRQ66ss6QXh7wFW9eK433H203W6
X3NidmQYsLTX81wRkzmeY+NVOOkTz2FzBOSq+TvzFR4bS3RJM8MHOQpxQzjhrHp+tHcYok4Zx5MJ
+4QcRAlr5Mi32Ep7aExMHxn6Bo0XJMkTSIjae7xNFbjGwTEtiXnVZE7YVB7h9uLofEv5sY1euOOW
fJbm5H9ekadzcmBJ0mAFt2i8x1RpC8h9SdzXXZesMZL8Y2jmwf5XeK9eajM1cjOCYx+EqCMXBccw
/FjM6JXwK2mC3oNlWxsBWaV0EkTeLVusmCpF3Qgl2OH5pOY+5+cQPVC/bfN/O9JH9nXwC3VoI0cc
ghfrDaMitXq3Uc2GndD9La2y/vh5Nm3Tyewt9fitq0piymuJin9u3ZR22faoeduSDl4v0lGr9X1q
MlxMsV2JyGUkh1l79+wna4UyDB1beTC0uBbQhOH4aCGD7zDzV53udSoQXMlMH2CTuuCSfzsMU+kY
UmL9NYtDmmAp0aAtkSklTp1XtRmtU8873imsKJSayLO+efB5yQMKawykwOOuP4xRJSM4UJnBTIkV
UYM8JzfM/vDlSh6cuJvqIkwmJLbEpVjUbFurYvDFcnTC6dCu7CSfUQFq9NwjW5oKIuFh/oP6N4j6
BP8Jsnzcia156bDYIADWOoraZtvvxQ4IELwBtEbD40rUcmgIDtblLPC8vocO4+xzkenvZCPHyhHb
vqhUEz9lghcJmyFZV9sPx3U9VIAdJuEYx0i8w4ri75Gqj11o1xozXblHymkK/gIoxuLE1pJ4bdfr
drKctFZhvzk3ugb8jgJBSIo+jqa+d0SaDMmjXI58lI27N5xhs367ANYNNJSs9JVyI6QicNzxoMNJ
4jLpD5Bzax6+sp9hGpUSkJW5dvGdNINzx2gguPd1/JZXOvRHKJgAWsoGfxVpgNlrAG3iJqt5+plT
5QBF7qUeSM702B9CGrgOrmA6CnIYiCS6/LfWwTRulHPujZ4SALOE+L+7XWxU2M3ozD6qMyEG74/K
Eps/C+MThZ8aZWSc3w8NBW7jmz8qybRjI3HJHDc5qp0ppELFAb7P5ah1MPDHh3Gc+o+vpcrMXOln
YrWEzF0Im2zVG3CvEinOd3VCjfE4VdQDJBH/shprEM6X10SmLCZgygxA3/R/gPH8ZIt9bUKFc8Y9
6eX2Y3WMMBdaqfHygrrCk5P9JM8+Sakg6w26EZAAj4Ny7GhgoIf1NRZPGKjfq2UCrmH6YPylZm4P
3Zj+Ha6SySg0zatoRUdfmjP5nkFBSD2YmBKzawgpWizrpE9R7BXMUty2qsAdlIY1ir38+JnIxq7Y
pjq62x1+DqivUb4nAf680xz+NhfXzGiRMEPa4IEqDr7gmk4KWFrm7ERFmG1vdfds2CetET7RYQ8q
VFC78YIOuuONGvabN6G4PW/sY0jx0O8QgN4TB/9GtMqqY62zg/VQYjr5kWBRUAa2lJclIZNIhtPH
GoFRUNk3qEAxEAOvUbzMI+vTPlq5thvMn0/TW9oYIhqo+g9qlwA3tGBfHsg6Z5ByeTcXQyxowHYi
lO/B6CQjlK07pIGTl2to6gHzxGxNYaFG0brkzg55U24PODa5Dn8HSapjFYtdV9Hoc+NU8i1qfg7N
+iUekNnLcuMK6vo0DPkNCwv108nCD7gU5C2E05b66pODHuNqwRXKEmkFJk4TUENNkT8GIg+mWfDf
6eiG+IojI2EUEo6iDISVnQgWgdf+IU51GccJqhNxvxsYbiN1K9VpM33NM4soBFhnXaje0HG0Lbd8
hHX1tIYVYH1qvBAPI0/K+c+Fq5/jR6edr4IxOuRQulQhLgJMUC1SIWvL9jkEVokFWzDRZLNchfEC
UcEyGHzhUk2458gdjxUW3OmwEhuOo6gGIGx/JZhwwLUY4QeukjSzj7f/l3ymad7oyg6qFIJ/KVFG
v+os0URmjmLZ6EA04gNANVmy11FbuhKub9PoryvYsSzXrpaYBPeFlxNRO9XnbWX/h9zLgUkQw7Qm
e1kfDEs4tRTlUzUJ56RyB4qNK3ZYAT65zyNAcOnZkEjYhJEwqTLBfTFJbpVnLc2cQvNol3SU6Br7
8vm/+zi6WlJw692havR5bO718BbrqjJPhsv6qPTHWaF9YlZ2EMneAGZPX9cmvpnIQafr/wA0rrbQ
Gz5EBWBj8tI3ij2uBjFut84HseUAKc56d+rco/m7ncbmGmB7fC2LXIbz5C5fIhCg1jS2kmZ4QtyR
VmIu1clHW2UuimLg5X23iQICWAl2ot36LNHbO3h1OS4ggGq5Awi8YkuQuXG/60JZvio29U6NF304
2YwJ7AW71QTFxCTl3+h0tiCOLlQ7lFgFKboDXZ+GCLY2g6Y58KKF7FoFlS8NpE4uJol+KLOUEGW6
rM8/9bPo1CLt0uDEmGCAcbqM+z1LrzXJWUOVeyotY3MBfPMu5Jn6k9EI5V4G73rfRpi4vLwmnPUC
QXXlcvw/jAfQfhzxZ5m2Sx8OWZPhKRFh3sD2C7kl8IN73b5zc9H5EOKDsXWOZJ5DZx4bmxJsL1Sm
GX7rJMa1WsV3kTI3ux32mkCiEGGVgpigEWud+YVCsRxAkN9H9n98VOkw/4v2BW6TugqKlLeQAKuH
HpT/ps94PQpN0wt3sWjihI9RZe0o2SfU+AjUYhQI5CKYxeQu1aRApAAIgsDhKDp+62qFSXEsj4Kv
o9d7AJZh+HqYKrZpz85Z+6FxhQqf3vjQHkK4ttBNYn51ejh5xzdnN62bo1gJEC09qGEq0GIvqWTR
YRHnKHZ1nCQRSICJCmyGqe0QCPWN+U6goY+WnrxnTLpkaX1MbbFsHT0tUFTtNK7ZmNJh3bj/WPdl
1ETFVQ77hNmudY+yhXSzu1vpT2deNbIvFOob8RlQdP8WwM9l7wEsp/xSK5Jty/N/C3VPvfn4zLsb
rePc4sLAFS0rVW2lVVGhMA/zsBbscs7QpDug4TZT0urqITlAL1hhFRx/9ECQdXYgTEkwYbJJeNV2
Esr2cNs8vefN2YldmOCwTeC2LykgfFCL3WWRBS2vb6MH/8sLI9ATez0Taq9yaL3kEPLwaw81zw8O
FCyDnxhWhoq22eHVgd6c+PAgQ1QrBbCftdQf8sWZ2uDIQsLmJgRBQtCbcakn/vOJLKOGc5Wh9sUC
Gm87KsisE2MkUyrChPXkZ2Rl4OlRDeghNbhXdWwW3nreqwz2QG7IX+ax+EZanjMGIwqFDLHtEV3K
Dlou+BZlh/mZCjHbW1OYuT3eDs+NmnfUXjMkHh3+HUVjA4JkaeI9jpC/Kt2PJJMA+g/TyMJ5DlZf
mvC4TRtljz/xJAs2v3gSHUsd+p+Pq9rn8dbyKxl5e5VqS9NplBr/fhKM/O98ldSp69crE5OWlKU8
9fsi2wPwsduAU282w78TAbNSM96x8P5paEK7WBQhgPHOJ3mYZVhi1bQWhXz1sW4zqxj9HLuLVi21
Hz6zAhBg8dKW4nXSloU7NS/Cp0uG/WSurw5vL96UtIxbF1sbcgSCd5U6EyKtSEY7QwlATGqy8W8h
jnkW1R2Lys+sV4dRZLLVQFvIU8F9x99p344APhwlZlqSR52v3hQ+DLDZ4DfTsrLUsqaCGNqirjTn
koxaeNMm4ngGgYIWamvsu/sfoNGgjCfZsOUqpToYoIJvDIM0EURVsH+3N2wwTlb56y6XLvG5TzRZ
KSK3kfKHAGzDRuaWqfiHiPy432Aeh8lGADNM+cgLgWa9UBko4gCefeTDKNrjTg1ti9PmdB9STeQi
mcGwLZldmLUAzCedmXB20Ghb6eFQk4g6VvH3gDDYS1bQw4+E6nOwebXH1pLMqYQptyMDnVWpSwnt
kUbo9IzqnZP9YRf3pBLpisa7PXX7qBgYRY6GnIybVCr0tGeSwJFQQ2vmjdnnnTS4kydCVUsm433V
NgLN7V8+y7AvXFCHIEIACoc+r5w6n5yrNRJ5iGklp+uuz5dknh3/nEQwEjvdbJ9U0RdsZ9xPxcv5
mLGkDRGvLHjbIODlnkYAeFvU9ObVspXNPupeTRk9hDd65SJJkvPSx9g95mHLsV0DuwF2rTGVsF/h
YPfJOOL0GHtOj3E4kCGTwBH9RklrY7b4iQDpkRr/QmK13nfyEo+aomKagOeaLrErMrEyMMxqsr7x
p1GunQfnbTipNtFl/TSDhPHFqUa4Of/7q96Gp4CPptgT97ixbjcGhEBzBMZMPFKykMJvf9aP+XUz
PzGNtP/6MPbKet11DfqlbWAwNEYLJUh0qbDBWADYNtRAGWbiTxGOp6KeB+sgwGOo/fxNVroxw9yS
g+EBWf+odHByMddO+YLO2/p7Bo0vjctOJh6wJzkdqZZOxClJ05+XO0s44FGVhUQiGySVAf3uUnG9
xKZAFi0HuJlr9Q4R19v0JUv4TNpCnwTsdX7WTL3xset+YXyezwG0U+frta2qAyuV1qMxBhY2FLG6
L7FKmJztarvNNMlcxTynC/7YnGrin4fdvpaxz1b5CTlHTf4UMSoD7SfTH0JFBhZf1cPIkoMuIZSE
4SNCMadIAUkApC8D77J45s21qFH4yIrcmv7pAwJgvBdkHnFYVdevoyXjwY+aS22984WasqA7D8bB
jP4gCC4sDIOkXc3CxQo/Z58CZjSNjc+G9ZDS1bRsgLUMVS4oPt2Lb3FJb27euqrCuszm4NkwG6Vy
OYH2dxdKTcKNSfYrqQdGM5pEe3O/iuwknyIzAiHngAYpd2CC6c0zfUhBQcLhqfjdryGsbZW9agDb
rnm6M1aFxQtSoxieLESym9eHxwEDvgGxfqbmPfgBTvjrNwO2R0Q2iQZel6tBAq2TNLN/ygH6z3EU
HlP8HVgPd3xuClwf9lq+LMCnj9q59u5ha6fVl+ZBLbbl6xnC3AEDrRTxuQq+1QbHYszEu129qpFV
1KDhLtNE2wmylPrRwyvGfIupjJYm9p3hZmUjU1WQ7gV1n6B0ug0JnJ8WvmjwKapV3tuUNRwZhERq
vXCCEB44J6uKof0BrnFPv93jheu2CQfqAaHNzDbi/p/ErWoew+5v+EXH+rjC3yS8C+M0GQ5pCOSq
IwwKXEshT63eelCp3BdULXpWfmgi6h+vf+ddRa1FYOuTNUtz6jWZmiMNPczP2nDdgYN11CUKi0Df
rCmy+DBMeazyPkkB6jfycwpVK+U29dtUkHuMmygn6wHSRI3uMCn+u8pDIYc9+6pevHah2prCiwEl
kJ733wFbO26gorSVRnPM0RsKoBN3m0DSXmujkUujMU27ScXOifGqsc8DKYM97feOjv/rpQ1iaxGJ
xiLv7SVTpNYx4igvi0vyenz01Kf+OZGDLU3kbiE8e5lBrF5lEbS/vdP4cdblTnwf3IA6C0nZSbVy
IV9L/kBzBkPFffnCDGeixZmsUnApUoBpI3rL3xOHVN6nZB/qtfx9Tl/KgQg/lZVUUUVMjoL1NQBB
jZctcBHMU8tmeJBGvHfyuLVzu/7dqo/HxghYMGZ9RkiL4VcVMCq0A9A0UQjmEpdTDdsB7KTeLeLx
x0QKz/cbHaExWZdcATaUXT+lRoDk5aqJZqlXr3GMTuVuogmEbNEr6/iunZA5yscACZNRjanjEAvy
VLgQRJsRqvSfutght9MI4RHLAz7l/UN9xo+sWw27VfTClY5KdpI4aqd2AAV/MomX+NgBg3HwMrpq
e4/ymQcTbcnzRVROf9+UQ4TfOIHxJIMb5GDoRBFUNBN66kHqh6Cl6oZUpKOdsnEVfitYw8bSRdtg
BS2XpJi54cV+X1sMkcc/BGc0cUpKkX2OSwccQLRxH151c7KFtZwGE44PUzdeJG6GchgYPetNvx74
safZS1YQci49pS99Z37bM4iSuuh5muJqAZj7xoH96XIkhQo7uqjzU4Y+zi3KzqY7EDE0/Zunvuel
Tx+TxlEeRBz9TjXhnB7dR2IHx2gKAk6nV4eUjYEBIM0xyIb4PUSWiIe5WddttaQDFmRuHR1aF57S
rA9HO2eveLjpZBj+wMiI1lb/XJl/a4g7GqnmShWpnoxhnMw98Wu7P3e/rl5HAb+l3PMdkWGSPbXL
SQw+Yy3xltnDCJXEP7jSWKCsIc2iJBQm2rQeZfNUYzz/P2ZNMMVHiQHQw/TTY+VSAhAbE/mvg0I3
k51EWrY2jBifiWFMWhE51sjj2yeYl5wAIU8lmZaPBCls6TCKDabf1yC8537uhh3Qu/wqSzUQ6aqq
Rr7TQlyX2jg0zY0K6np/YD5ELAVdV2/COSUVgr1wX3hNOH72Lt6LxhS6V73JcpxcU9IfCDY8OrjR
992kO/AxUDaZ5lHEaJaK/pfLOOF6Uwq6/4/oejbapKUxZHPeNE0tk5UGDdQNc9nqV3r6yUVBB6fl
dzj3r71TEM2G+Ys0/rmzI+OlraG/9YPzKwavJPljMYEt5AIoi0AKaP6rYNDPOrRA1ICytyDMeRyG
zdHaXDGX90roJ9la7wXDlOPXCQ53LuzZND3b/W0EhyiOW9to4ncoxihohm81PLOdPvtTFpB46sAi
XklqsVoV5Yq0gpsjYglmARYtEnuX51lD/gd43CZNgGySyyrvgnHntVPBHF79hxW4b4LbuAqQBEYW
xHM7eJ7U9IIu/WlvN2QWBD9dUstegwN2aqtzmw5rKsIDnmv2m/wI+f8bG1K7WghjDgiflQEnvm9t
9/bpYccbr5V2jPar9RUHTz/Y2XHd5mubjpOQC3XRl8vzN8M1l7HVC/a4NoIzY9P9voby5axmNhVD
PvTqVE+nChcjoELUSG6V6pRKmVuoBa6l2E9xv/6SFowTuQWYeB5Zq8pbpjU3AJ7J0xh0I2Ztp+SO
DVWv2BQlVVasOrtPgXdvXgeUZJZuu2kt0r8pG1BMC0uvWON8PASbzj91Kvomd2vscbZb0kd1HtLe
YjC7x4yan5U/3YG+qP+bpyWP7Dungru12BQIoyly9V4+D1K9Du6IxcN0Ecr7NN8gLIAj9RY7v0Na
VD1kmYEoHsOPVOWYhbWtd0NiO29n6pWsaFQSmFgefYe0pEhkQlPbhIaL5axflYoXaW4FCtreEUdi
h9iXhk5gnJQ8X3zZ3kQkWL64ywh5EiI079QiDII6gTOwAV0jaHnY6efxNscyLgraroJcxukB7O67
Ql9UmZs2azKYgPjhuzxhdLV0iHI9fVN1/fsM8kxCNc/aIoaSjG1z0soPZiIm5xi1r+JTb9fpguEm
bhiatFifXt6BbhfXj2wW5GhnArpd3PZLKU4Z1hHfvw/4bXwrG1mCfIpyKB35GYh/U+glbWMAX2S9
qRLCDg/h90jr2oGkOocAeNVc8dcmEDOJqqyuPmtNwxfrsOePLf68mF13BABVJNh2Rnek/8D3Pxy8
G8jhq0WgsjfWffrJ8EVv3hqGWm1LY4LkCkfdAbpMMbzfsopLW4S58GH7z/cIUyxeqvCr9TG0TYkR
9W1MK5RTLa3PXM5+HfILa34PXf7Tg3rSrI+q0HGJYnqqGAnHDovhrA4hPFl/FPnw1nwao1LJhtFa
BWCYcD41PERkyIMHILOx3vGemn9sTDX1trfvTsAyQi6Kam/32N2BwZigxYUQ15RcrgfjrEenHELm
lR9d5415llvAEu0bKonSdw/h+IIDPVV/QGUdHJ962Xk2dm4tQaZOV9HxssjPHGfZzI2mH0xmuhoI
uBlr00jh7PrTx8ZqKOCOOZguyDI15Y9A1acjHQjBuHQRUny+DOTPpuyvWu21hLZGtpgl5ZyRty7W
9+tHHSGkdW0dRndFNxBROeKy8NCH9QCh4Hh9nbG9YItt4IRplOhDprdCTWMd2r10pjgfdBbXj98y
gEpDU7hW23ofDVjoWEyhc+DAFzciUg+EiUAQTO7Tj1qdP9WKFxJ0cxlWJqvPBCuvTKsGCVkpp63W
J8r/xuXhed1mXCU925nHgSVVnSAmJri94wdRGIdzj4O0zXjVfx5gbWfsSiz6NnGR1zBoVzO34gxD
Y0kLdh0Qfw5mI6foF3uoUEigqU7KRhR+Y5RUdjvMVLz6vq17vMh2g7eoB1hNaXGgkBjuEJZj1BD8
6mONUG6UiG2vLclI934Fb1d4f5iveAxe8M8g/M5CgJrNlrqmt/UdqYXvc0Ttkz2p/IoB5nVEjLxt
1WbsI4a/jIncAoQwypj/R+gEv6JiT83F4YjTALMan7bvGhn0baNLVTgevqlFqia2fJUHSztUA/mR
+4KuV8Vs065QUCR1WiCziuiGuXZ6wOMsr9Li/KEExcdxMncCUzn7tHUrCF2z/wQCSaCQY+JtyOEp
pBVJjcF1f+Tr0FnpOSm/V8fQa2JaZxzy3Gwgx4ZvoPBgmLVfiTq/UjADJXhoPNZgLHAho5Pu6/nS
sHRmVzQkLxHIdo596gX2fw5XJOoJT9ftpSVyqAAntMyOI1Gf7RBzKkUBa94dYitlL19isuuHBW+g
fgsm5VVxj4O2E3TM3nxC8pRcbfMiWYbT72nE6osY9437HXbWdrIoyd/ON5XypAvpEAa9OtuCkwNU
zekhK629nBdMSde6+MeRHqpM1I6yPCf/ZOOjfHzMb4p4IOESnsNMClRzRbRzoXEYRMIUr4EyohCs
Dy+iK9v/xWc2i5kNLl3oNVMUr4S736ScQOq9NEwyhOcXygeV0PQjXfNPPhJpSClpjOKt2B8kz5RZ
S2YtDsI5tTvl7ca/K4UEEKROT3PwFwWV/yIFlN0fy+2EQzA2uLYvWauCm2/nuJjsnPyMBulCVtxW
UpAE/2AcRndro4tXY1kLrVdr8damW13RSW2KH5HBNp5bzfEhBX3VwlbZo+rg2ksvxzHmE4Peqs9d
8tJLnA60oYvhIpLcp5sFwW+HixX+aAq0P3CMf0czWQVJY/R5Ts1ZZCyYSsvghxYC/2TxOONM8tMe
fEtnaa3XHtugNJTJZuSX7uJbMD/BJsVx9ubp48/BdWMD+ibeygyupsvgd5QWghGrJ+inBins13fe
MNkpPad2b8hS4oxVB7OQbd9vpNHk4LRV9RSHYBsMnk8urL5ZvDsWuUiloTyG8RWZ2k/G6YBIukJF
NQxGME276CDgYJwZwVINOvZsKwatCviOtaZaZiZsgUPLOQoT1T6M5uHdbKd4XU7KqOlxhrCdDTOk
VM41sMiqNWkV0lOkPF+hG/Xjxkh7VwirVJ33XpIMZLayiMxf1Jrkq0Q8k7sIzieZAJb2HeEL6eq4
jRy8SZWRoVfBOnGzFXa6uq7htKKXYYC9uniJlhiy9HG0tq9ySQ/U6Z2Dnn8TB4B7D/xwLgayldrx
4xGVrQ7jenKzrgOtO7fxM2z5MeXZ0ME/7l7Gzhtrjdy0vS7uqRGky0OodzYMRzKGFHxzJUFprG3D
8beJuTcd8OXcbbvekMl0t2/PUwuKGMOeWGSkwZWPkt6Y5D19uTq1ctikRLDKZvF1c3Loo/MwxSCg
mlTZthesZelcw32Dxuf/IJF6a7Ls4rgA5rNkTEabKNs5MHILbqCzVoNuPkZYjCxSkW91X8uG7AKh
mt2x8OMnrjKmMhE1NgDXB3UFtXRGVPQmaZFHyht7jUeTjjkGTUTmxCcKWBAThFTEU5ErAOEqEy24
SRfZBrwjXbJomd2EwGwz9hwSL02SPiqi3ZwzA0OWToeZHnbHPI7xvz3gBwHzI9D8IgVWwhYcaUi0
nyflhz0KEW08AxF+pPzYsB13+VNc0o6lQ8lcOc6Z4XHh/oDa8lAgVO1O45o+j817RRhIC7Gw9fu9
YUWj9WNuQNAaZkDkYtRAZ3lxJjNJmYJKfe2fcJE8EjxI4VZrpSmXnsHgP24N1vx7OAcG0WmSH/eU
syie77CSmMY5KcuehDC3CKyX2t529NSn/pB0CLzc2Q/IoRpLduNQOWVEMr//mUVnufGezVXhPlss
y4U98W8s0B+xlB/PSKGYfx91geXy2K8XZiBeYMOqFD2jZ9M1aoSjwHRbVpss2yB/Y+L9nbYhqnPz
XZrBgU60rKwWZAReA1SKBH4quqni5a1EPD9i9oSx5p1m/pmZ7BzyJwTtVT8OhiCp4xKZmYJXXW0g
/CYayoOssmUcpQZQ3NClaFlk6IbXjWNHj8+siL9mMG0FrH4kP62054gSZHzcvaTiHDo89fQuXFXJ
QvCw1KjYyr4aCa3SogsdJ7nzNBR1PmgkErPhALj2zxrGDPeEaffHdRRyauCk8QPKvSFEutVMNWlu
OPiDo/F/w8y6RhPfzH/Gh+DhztE9QBXf93KsVv3vSxe+aJtGrv0QOT2q8QdS3ZmqtBG+aaYwTM8T
wp28xxOWsKLQZmWeM8VvQ644ApkUyhSogX5sb4f1pWJ7etHWC5LipzNz0G7Rlx8zLlQuWOusZTD5
J9B/AnN+B+Bg0NlVxqRwYs1qwr4vmbwm6EjLJw+D+cQ89/8zafJeHDp71gdKPBw1HU/uS/KJweXO
utEfEu81dYxaGqq0dq7PL96Io4xKKRMtHwmJVKVjWOSpSRaQFu7O1oB7EPdYvc3y1imsBp+nV5lY
WOELFdE7x5HIfu83XCDQJr5xYwOnvmFxPKohoRARQwKuc3enoOcVgcFt3q5wDINn3UWZ8VoNZF0M
RuR2JZStE+igbKm/j7+YTlCZbflDUsLBg0Z3ErU2E9khwAc1XZ0IBm6ALH56FYL84rYCZ03nxIxt
dgCCbex7ZWOgm8hCZVFoQtAcDt76Kly5pO6TwHGiBqR0xZUVXUlPgokFij0j4A/a6IvKwgNUoOj4
8XwBa/FSbKiUncYS2ItMjq42ciGf5fTTUrUlcqAiTIzya6wI4IJKd3TsiP+tFhqQOXdSsj1m79Uv
pITy3425/dsYO17DI1DKZ2z3T0VYykq/zC5LQOjwdBFNr4igIfjeGQ82M5lAPEDn3SVKJL2Nro76
O6zc0X9QUyxHVe7JwEhisTAoU3mQ2vxOsxfFCgZ9SCx2AMKSNkNmRV9H2wMA2qn/Y+zuRzmSfuao
NW4IXWBd7fm5VXlG2IW0jlCTT5ZogJpAMdiLAi7Frb5rF99ko4tsSZVRxJ9B/9OoLL15UTx99egA
a4gzu4cwKT93zLbHA8O5t/+vnHgOZAkaEn/6uxFJJd8yaUPj24rUfk/VYUXxOssRYzEwcoBmiw6D
st8hsZBZL+1GNqCx9FBDcZLsYgONgU8Wgz8EWZZeZqkLFjm87B7za5IGZCt7VYS50NmyuhhqpSSS
lvhPkG16z0JCuNkC+PCANSxqrwbrb5+33fUN7wR8fo7rkaQMg+9UfKQiVe+Lk4pfsBpP3oqHQiH3
lX/weXKMyKsxpNUXTtlKgn5DkHg7BGca8VqarfT0wtSlm/nm1BcUdi/oyQNrHW6QgLjSirRMKCiT
9ysZBEpcgPhq1aen6ZJiSnCGBC/6A9RIcY/xxpapU92lhpHiUeds6eCLLP9XbNOLwgdFDqdOiErL
19rWfOfDnPkuEivnQymNtmBhq5eyExgYRNBS9D1R2shNDYcg4g6ke7L5oqZf4dJ1EfLmTbtcQN0y
gHHbBTZRT+gC+HIYE5Dd9dusZcEdXf8qdNYVhUD1WrnA9pIh77SXUsvalgvuaPH02YPHQa5PSJLk
yxevyV9Yp4e8LZp0gsYHaa55j3vvajCQITCUAI1O4RMRWvB1jsuYNgM0XhhCLJRGQQgf0AjkM75B
Zp8IeQk8Vr95VyEcEqqbCIl4sVn6wh2tDdMTScAyWXBtArd1dQGTxxVm8rq00sHoAApJJQe1WR7M
cC4YO4mqLV9nVFOSg316FklzHbplpLT/gzVBqnoibbGOTRQXOhhjDw8AmFAw5Pa4d5cVh2BDnEsc
rbdGuHVY4wk4UVdt52eduBKRLNpe9+uyeiepBvCeJAnw3zMXWIgipPahKYQy+7FV1OWI5wc6V92c
tBgLRo5WDVF3NMJwpAtLdEzN83lVKWTf1+JAP2/pVM9i8Ylcys+nK4n9O8T8/J9DFe+W8tPzaOr9
CEu3JYOJHlZe5sXP/B8eOVZej4EtXzITyjVjkZBEu6VvV/AA1J85z0Mjnvneg8a3YmlvMEjbp79W
I3dBjhWgLd55ZGmZo1RgRKNjqWr/ym20iHVMevrQOCOKfi3HvApdpFJRm5ye2kmh/xMVJLjbVxjm
H6PdYL3UGgZn8k2pH4v8CvQK9bhSUodlP8km0jWn24AU2XLJmSX5RGh9dYJXxlHZvu9VLG+jhhwp
mUUNK0pncykKkOdRAlwO/rXNhz0LcRyViFeBrLYfV73GuKjQoz/xJ1Sq20NDV3Qq3v2fi60yaQoa
7AKxjWYvec8IEN6WdJJ8ZvIX3tS+nRWAu5nhy7TN6fTuGHpoZ56bZt96OjNUe5asdcGa0tEwgBzf
g3mWLl7I9iVcqPo94BCptzEomO2sghODK/qBOEN3qPfUAGxs3c0YtlFVVoYqM/0YIvVaWIKQwZQR
oM+SHrucSYk+Kpq0PJ5ts7WeQhxGmnwQZ44Zen00uh/4PNxv5YivTU7ubltS/omwHleW43mtvmpH
ftsT33iEURWxnoelYh3EIFbn8yyVobH+3rkBKlnZJ6hqry47fQ7JMTa2+OSgzfVY7A+zaB/dCL+3
fFjhGkNPIjqRJ9bhzozgLV9tGoL0lFaNj063Q65AvSqnk245Wdli6THcvj6PN8qLaAkfdbKK4vER
Wez2TxNvVRLhF4zWZrr2SuyQt/2OTNnQ4eeltDMbp+dnu6rQjhWk23+lViszo1B2Dt444oCuZ+7s
CVCBXM20rH0URX9MStXwiwjw5md5m2+zpAnp0tig6qEXBVcouJwGqMm+X0UALEfxQJDnBXARYD/f
HKHoXD9WW3xZS2O7v/2TwfjP0c+k7F8Zrx59j0y+tqc6ziCLALUmbS7rJ6Ieemp7KL+qBuMbHJ65
0lnYrc+LvWl4ZxS1djwhFrHD4+g5HtaZh5zrQVMmPvN5M4BQRsbPseZ7Ldr8Mc+yEdGa5wGMnLMY
rGXx8VJg545Uk+Oly5/gDafnmwijfPqLwI0r6ycuYu75eY37FUBmxnIS6Tq9ROU1JhWUir2YDQGS
gICQyxH9GsTEjCy6+pIyK8muSrfjVlg1mWNkfkgjKivS7rH2mc6dEhtlH3NEBIBmCkR3OHaAQwZS
Q3kzcrA7qFdovpJEpyZdtNoclrioq56PDq1/KrRH4eJmfstYQozERMWoqkQ5qpnsw+UR6+NUzA3o
vPHDthwzKkWtUzr2xsSSvXui/kqbZD/1p649MUK1t7d17Mhnw8hgZEVLvm6YXr1gtPRW/bQ90NNw
VeFQK3tG+8fFf4qbYCL6jmTN8H9HI41KlQJhjbYdSA3gzfampYG7kADE7vgUQ1LQ923zPO2zs/8e
/XXqyKLXxxvjzrF5Csy7jRI01Wc1XP9ajQdWmFua54DJDmGQS44lwaBjiZ6V/V15KDPyb8e6YrV8
8cQCIntVG+1ETnDnsUZsFO23nu+s62XWS5BRSs1kShRJ+5vufpauqIkRWjuwnuia8jrrFSvj3EDX
nTn8sAMqb3vjNxi6eqEA2D0UjjdQNAclPQo6Inz5gqcvORie00j3pgyiW5CwrsQmO+k5nQ3ZOrdL
vRbQ6O20T1GMu5bJgsVMAJPlhtNRUIW0qeyq6shw9rU0L5ErdqmloOR5ClRQo8raLpp3ocQly6QK
5Ri5xYfXfhgq0K6EvRnWqODmyvM1G3NETcxIPb0dqXY/xPCI0y2ttDhqBM59SW46TxvI7anKOG+W
Xd8owL0xFT/hI8rKg3+eXKaGgC6c07RkF5/AxqUOZ3Yy6SyBQcH6b0ZZcdRF8hzrcX1qy36CHnl5
tFJ1K1PTED4vGGeJ6u9HxYVg7cQyXzBe9Egxi5HYWnTef0yUmPansysahmD9g9wQmMZ/zI0o+5C4
Nk/qAXDqqWq/Q3lK+Ufeb9TyyTRzG/Wsc3venpIgtZWpZUKOHVjFprdtCVoXqZKR2aPMFYxp7TkL
BMPzjNISXkZ/S+h3PJ7S/PIwA05NTSeVNsFxA6X7rjdw19PLoQDMiAVIQfdYEmviEQevj9RgkzWU
XSbHJdKAiCskCypd/He+DxUKl/aobBrT1b+00N/90P6GVCBDk3oQOg76Jg6JpZrgH1546v+G794u
qZJ0t/L6+YUQoCJwBoi5TlCGW8FYoUw9EdlWqKMmJVhM1hVNsKAuCNF2ue6+MCpZ1mIB+Az9YM4R
8fZmMUmB+oo3qKjdTT5xDexxo2xINtUnaimI5iQv1UD98qGwMDYV4nN+T4xnbTlTmnhxqn/GczpP
96o1S7YwEallVXHNVSx+HED2W9bYFVjW/9TibldGjtlIMuF05QYbgadPPV+Xy3cydP1ET6haqwJ5
eF91mlhA5abS0/KLRTIagjGzLi7dBdnViqhNqaBtU+bobjeM2zFWB6j/+P066LChqIHwuQu5A2+m
lC04/jsNRK9lto/Ka4rcdrvX1L8uivTR2iuQFNe+VDqxvh5ZDEcIHk6vZinCCFANrv6Hsi8dS8A1
e45LDDWXDRLVXE/pq8AphpNsdH7heuir4whA/I0cr6fnXJD6JPGfroLUWcuE+rAPc+o4n5RZF6u5
denQ9kH0ZlKgJ/XviqMIDU7gPgtadKqqUe3x71k4tDDi4EHgkYkBokocY4+H2oq5kvQ6VQrWjMwo
fqPowKRFUBIbFLCM8LYgBFfHRm7Hk05x89bAlCC+1dZi2u/LK0hsTeMUwWCMFaJLjOmZ8x8KEIlY
4CstZdu2pt15KDXjL/XUUHNtqOpYscw7TJ8hYEoBr/hta84apaFGYKNUWcC1fnX5DvC8M4F4tfcn
5SC6U7tgcEnGQ9/sYREavs2NNf8gumGFJWtq+XId+cbiFDcOVxF8cj+wMesaxJRJdqbYtNVieKaQ
yfAMonF2qB0KCv9AwrO94spiOcRO2MhouIDkAFRvwMjzFHZNl3l7eB8/qiv2XTuO/PnGOq0mFma2
uhvrxCTJxJLk7X/QOmQx0FZLcfHMiQqj7jusLbR71EFldQwFea4PjNB9tzkLWgWjfTBzDA8mVBq1
gqkKhwbGkzt1dxH2CV1cXmbi3RoydLtxA/ivt+9adPM26ZIhWl9lczXr3nCsg79KzM/nOEFotWx+
BL5LS6HnGHPu8A5TAuF4NnR9Sho+y/jc0D6R2Qt/7EG2bl7wZHK4K+r6p0KlCX14vMLLKn3LTfBK
NdoCFiDp5+QHmvB7Ntd1L/1rE2O6uW1gfeY/4TveQkOnU8+t+bqnloz7TEinOwEWPMPWs6WnpKnn
19hIMV9bI8hR62PSmpfJtLMYywSEK7VPF9105RFe7TtWxEcJOfqruJQTjaSBvJSGXBLsBbB3jOoN
wIRc8cJtNbLf/FTM3uDG7DRLG1GUFM7nqst8rhpoYANBd3oakLc7iSXDIlboyJUcPamE83uC6rJf
vLfFu64zNKDmfofHTvn4dPuhA0HiAxUN9XeKfsDqLF/IyfuC17KbK2fmC0GLtRGMlh3MUvyNrCYB
Jn5nEzWJqfGJbJfX+v0Oirapv6wPDTCMr2MbhwXTydEZfoMHtZ4ecVKkIDKVjknM1b56cr8TGp1T
/dLpY975RoBUzowmQcrYdlNB1ehMzWJAewiruiERhyXIqf3orssApuQIP6WSChp1/1tr5BviYRAi
LYQfwEmQkORiHzDO+qykmz+NzsP2BYmhFpVbi5maQVirhZa+MxFRhtAqTgdqCceVYRzS6R85Nehl
OmsS7K+82rOhTUXBnFioG3Z2jnhoV9wC2CeXJYPqmJQhCRAKxZdRXZi47jkblY8EpxIw/9AvURlB
OXLQkycCg0xtQXofksF+U9ODlfLpoZiEUQrqQnVLMwbOtBI1ZGwEK41+Fhl9RBz8PbCDMcRGDsRj
pkeH/66lvdkDtysC7Bq4118T+ZKsYV83wGwp/85H+wgZL6Y/pOyE8tA8nQKO5FyhShJgWiwNHqsn
9bPQVkXRw3HCv9NRNHDdHGYJUn4tjy6/uEGGjAxFaRxAXG7M4GJDryzoPDC6nVNn0ViPVadE8wbz
/AN9DOOpm3ydTWb3nlZ8anC+hnHcX73jSdNgNVOdYqJBWsB4Dtc/ABq3D7N1MyOmZlMi/y82QT9a
7Fc0LFoYIFKXF3DipZ9Y4zhoa4RYJZuuNqW9Gq2zkRC8iPZTB0QjevlwC8PMOhna3wscvt0JDuZi
8i/0oW/i6bo5PidCxPSzq6M9j3+5lqdUkNOKkyxzQvfKFemm9cBVa7ED/oM0pmPHdNJZF4GUvsnU
9ILMLb3Me47a15EuCZVaOFVPKl928wUAXJl8aMEX5jiZC3l+PQdwTrvV656Np7QzXKZ/2mGKagAK
Rsj/RqGbH3hCXUZxrZ6E8E4ofWZgkmc1GIvsoRREUZPhxdFui7aEqsY2h31Jii3/DDTZTladGuCp
gp8j7q7L/qT5Fo6zt4vaamVrtqgUB9u3BSHHXE8yngcXldg5Qwosacwm01UDwiMJLxowUB/kFaLq
cDCXmRNjoAnMNecsSGqvkoXGpcW7xagBMQoIkbaGYOmS8WMF91OLCP7a6jrGHgIxCYCara9/C7oY
7yT12fVEGWg8MAnF1V+njgA5OboHxO+AWUzcispcAcLE6n8xWxtO5GveniDAK124p01lgT6tlqMM
cfuswVUsVrQoL1Qhg0NRfArJV7iH6Kkbanqfy/8gINx9WcvGYMgIB9QpDho+YhPIvgFNMRZPWQ2o
SzaDQcaB87RbfCWSweSU0VbwKK9RvaVc8F9Agx0hjiOBHNA/uD06hAZ0ESSk8U97SOIEgRJdVMjR
H+tUAQbjqyb+nGjFoh8dFuFMFUpwp1nurPGKlN1PuDHTP7e4cp0IyBimQZi1aS4tT4IQ2uQ67gRr
kzqxzYRiNaZ4lRO51DooDAKtQyNKaeAroMDIo1IBDceVKeE8oJFD/NEa5jqy3KnVwj2pB0Tw4LBh
94mq2GIbbiNssiE7N98ysrmMCFtf436h88jIZ7J1zD/xK61AVnWmEGXYSjlVCGS6aEf+F3YjJBAl
7YIb1G7kQXZZTv+3xOaKIdZIsjzk8lG9CGLaxGj31wh5sMA/LJtxHsICgCR2dM8eV7htaTrJX8oH
ZvZlifC3UjI6uetUZmL7M5hil/dCO3Z+JiNMxOoaKhSay/eN9+X47XSituke7OVGDIHtulQuyZ/k
9Ni9NRc6aIgcMpkZOd2nbWpowuxFxEf7Yz22fBE/fvdYN3SCtF/t0F6UQwfhSha5a0kZm2fF4nMR
vGslwkccHBn/eL6OrtOs/Zo26FScuyMASVhrtq2su51D4weW3kRXopqaK1/iPeCOhlpmZRsJpyUd
zA3tfuBUjqmFEQ2LH9Kg9QuFF/hihLoPIR+G5xRrNQP5rIQFcOw16tB0rsW7z70vrSR+oRjR5I2w
yF5/QGuwWlhzVwebUQxH67SJjI4yHdlT5G3/wjcUYPCprZoD6f4n6UAbSwMbcWXcGsgcDC5tZA0M
iT3jb1sIiP9l7jL8UjBfUx4u50KcykI2iYVMgF1ZOENqbtZkgrgynEsshi+jenY6ZNnMK+57INjT
2JGXFyyU2+oTHQjXmkcTyBa5Y6KwJtAEn5iGWKFMD3k+YpwZbM8MYxthdUsvX3ObIC9tkRbBp9r4
tEb7Tu9YqlVlHtHpBokaS3E4FvVoPG6xe6rAI+RCAR2MDzidxzDXRM+yFosjB89YIV/sBxOHZdRT
e0axQ/U51olqz5bQP4U9aI409DnyVOIbcxJWnshmuGOLpieT4moHKyQiIDXvi4eb67Egt03DtRK4
csVhb+MCXw4xHGDu6LDsDNMOwJjcjW87MYNPNJdtgj/c3cuEhJafYFWiQAkFa5ibND1j2Oz1h7vh
+Q88PincMoF8vXblRoHhiOMkZClzGGk8O7I8S3SK9sWQzLXzffJeY9jmpLjjWpAn6DyQL9ZFPdbI
AH0M+hlKaXb5kWVYQdeEH1vTmvuqgb6+JNqo0VIcg9ZHI1vMT363s9FKBWnPKvprc9PK9ya8KxyW
kgIBOiZoqdSnY2t9QyOYaU6VoqWkRUepKEmDFkRghVZWH44rKCjb3edTr4Sm08TacJko43UsNmG8
/a7SUNnosMxA82b2kn0o16K014gEonug0QexcJsVS8f3TmIm8UgmlbhgSca20YEB3kBllnOhO0N1
ijcjuj2pMMQN4vBKVf59GB2Wha+NcmAI2MAX9AKXg2PnufAYGu+nFlstKQNMBJJFH5eg8uDgvcs/
uIX/4UbViqH3z9r839b6zFFptqg7f3B3EG9HIuxtEGVP98eLiwm/qzZYD1GncmQbb1ABb40QCEwU
dOmHQgJo4G0MMLwNgYhLWpeFriULK4wkXdApedEvNTdmMxKytJX4NCucni9ToOtSHgo3eg3/NynR
NCCll3u/JftIBLlf0S3IB8pQChSWk/P3+pzAjCJYgg1MmMTaUNxQ/1AwLJ5fAKsWRx10PdRd+Y8R
hl7w+Sr9Bgyi+ckWnURsv3jV52lmac1ZKalJQwVtbWFrUml+q/ncaW4+USAqoa5VyhIXkRaoWiFj
Ha+UlFQkUw+OGkwpOYx6e2lr18ew0Ym3/gxgiv/jmOYYQsQzxuvIYgjE0BRCksdJxzOCLel5KqKf
kmHh+IgGurTsgwLYShVoAROPiuA6fSOFFuN3C6thYvQBDEk7MzzyxkW9aAw0MzwLgnJh5ja/UbKu
JYzjGVxS73TIi7jaO3mQ1f6+BkNACbPXfBQUP0A6LMgIuiWgb8NGJoUZEoOIUd/FBtK9TcMGQ50r
oA2n7ABbt4YbHGKxRN3dN0DAErVXMOL+Kbr609evPstx1ia2fF5Zu8RXj5wdL5XcVXMQuW/GivdQ
XkFkBoE/iNVxUNOMXn3ZlHVuQjKJm8uf6rc4Ja47hTDXTWgAW45d+hT7JWp2MEnrgSrbMoewmk4q
y//Qkuax9WdrNyok+mD1Kl1PSy6C7+gKY/shkm5n5Ps+Us2bpxhcV8DczLORGqp6iscUywtSpf9g
watQOABmqxSVcxP2f6HkpRS2PQSO1VeWiFwzZS6Rf1iDaIJeFb+oNF+VfuVuSH2hbZGLpgtA4g4F
dWDd/ThNHR88EIaQ2Qlbwd7t0PifJPrtUGToz1ym4zMDJwLgPHmrOZi/bh39IKb+umSY6RxsYfhV
XL0YofHMrDwjjRTZvXx6TboDtDzcuJaXVN6HtxdWWWzrmM/uksMYDl0MdoV+BO808NRgF4WCI0p6
ClRLWhLmFQ+sil/1DeVwKdfr9Nlu+aPPawge6SZnIMSd0ZfbWuvVQUKz637rBdQOCvHDGLt/qu2e
DrsIOEklNA7tmjdZ3hN2vNvMUlmaKo6TqZdSwXigbg64ogh3WTfWjuNrPIVkKVS7U+9/tM1+L8+Z
jgb3T7B6AEjKTKoH0+VerKnSTF4hDZdvyRl3lNxkIaaNxWdPRKfIH7iwLKVfdahhBjsjkz833CLd
SCFSCfCC+i5/UmnczzQ6maQ5Y7HSpUD6t8TkVHlIbThTanrmvqMuukOUOIXSXpPmbYcu4klVpzDp
7ZWHv0qHGlpRD+55e7SbnVLFVv2A4LQSZ+VXPyPYtDi865sbXmBIm+lyHIxIxBINOS2dC0I1iZxD
mxURy51A1vdpCXFCOYLm/zNwOa+1ndS/wJO6e4CWiilbkHYO8rSQt4HLAzrwcz4tV/2w5xTv9i34
8OagdnW0KrW4XX3R2Tnb7AE69JQpaLnsGxc+8WMusZ+lPvyAknB48+2iZ5wX+gu4PVs/t7QG031I
Y/U2JpS5HHA/TOIdWoF/LOn2jYmrmDP2akY8TUvF4OJSotfas1dCWoapHhdbfxpuUAiOkr9cZ2Sw
GC0TdlhsOMQ61GKHiNOfGN9BZK4uaiEZuedjQxZ6QyePWpvmNMVQDSRZYCHoDO5idYuWT7yI4pRV
aciaYXvUsfnWCAPjvDDUFZnrchUR3m6F6GNGx+t/3EAS1iKWWi3y8Nkxi1ILq7wEpbeAQxgG/zjl
9MOrbhfIgTLxYJjKQia2zBI6mEqfyDCIe1nfsuWepbGIHJymateIyI1fC93z2kiNJ0yHlrPQ6eFp
bjD5MjwTENoAibfKT68Zw0O9Cn7CWuXem0Hfayo2+Y6d7zBTj7eFE6i35VTG4htPxyAw7EH2wiUc
VJtOrl/FXV/2vkQEwf3eNE++fOSETYNDshUp1qQcqA2/U1SkE6hoo68NJ0Npq23ISFp3VNi0DcXS
3iSIJLfEjar0NGLuCIYeUhotGeaoYPLyxyhPl1kaFAXetLY22JCEPSDMsiaZEG/BbnQ8rjICZT6R
5LwdkkZD5R8v7X5E4oYAyAk2JeIngHVhVSjlQu0bVMCv6H7QJQtDYcshxNjCKPgMxvvFx2C44kd4
RvnU+x5mKgs5tHyJpAwu4mbsg2hBhrCGaANAAOl6kA5P9GSE5GrVecksB0a8/WTX/01D5Qiv7NuL
3nEFnZOc/tW1WpBVsIzitMdaU0PL3P/eERVi+jyLc7VuyZX4gn+CwhrYAOM2JHv0iUtWKca7uMTK
KAwXN3mYtL7cnFiGt+uhzBC8vdunWYZBgC442nrGhpKv9bzX3sLkGXgs4OKnQ7AWsQJ7jTQ6EX3O
xDjy+EZXheBdbufBcxt6KxIcGmHHgcW0cr2EbQNw944fKTCpx7bSxuiDFivObDw8//27I0cwd1r2
ES7CnF3d2P7VXcRkEFMbmeRdu5lQiobHiWdRL5URS24Av2skTYnXSGlM9VLIaFsPednva6KmS0AY
Iwkm93+3zmVB+Akwhudqh8uE3Rfy27IDgnf0OM+m3bByg4ZkFast5D8A6lZ25TgJL034MEmZD1nZ
tzUfZqoRzYYY+utclI9M6T9MgqTGEtJCU7Ii67NMt7HHQk9ZnClvmtu+hB0ipFC2+lXrbMuWi5Ol
pnNALsUyoqDfckFxZ/HmkNl2DCaYLsb4pr/WqDZ+RdsbyV6pM0gdduu4QbJtTAL6ifTMZ9E7Kgfj
WC0z/LXF5jT/D+w5U1RzsMRkmHdXSNwgYtWC6MdYrekfo3Nb2XnxYkDjVGdJtb8RYz8WB7z0mlp3
c6YTkERGeE7BPHHvePM6zyS6YubgMajU6CY6V4G/2/1XE/J25hAeYdOUJM+WXytOBvzhFDQpH99W
sArrhqN1IkZRUAZBKpFNQdi7q6hQj/AfvzWCEmA43IMNeHxZjM0WDxyx41uFXO/MxnkOEreFkc/q
Y3bjZtayjkaSPilUIxvPskyAPyDtSj6zMew6NLSAGuQIU990JmC2LfQ18rj9D9FeiVJdZF3Bgh1C
ALQ0xsH6mZl6aKQLq7qjvgBToxBmbn/Z0Q9IN05Q5iGvM3YE88X+prggfcquymnRm71J/cqu0+yI
axg1AEOg4n9k02YSJHeY/fuVkt3Ww5S96Ci2yqFmgmmlUZjBcOK3P55FN5aaiUK/4PpGRye1DbSz
nI+PLdYw0FGnDRauIkLqjwsQy1iE1dUPZhMMZfK3FChYxybRfAOIdE8MO8S+6bw/aMrQIAecIHu6
GlUe64m/YDo7TWr6iGQok+h/NZxs0D+1qIcXnuHQ/WcTCNZQgybM0domN4hxlZokzQsbMUuh8DvX
iuWgeFMp8r0cpS/pU3Tt8nAyuctULfuLYt34fcyFN7Vef/dcjOwlEjeQHTKdsy/t0mSj04+3lMPh
QRt4zFsxhHJWRlz+D35/riOtu8CsBgRDlSYP6KQExF/snMykQbTufux8QrqHh2+w/5gjNsaU4RYV
dpDeasfXlkVs8jqmKLTnQB8gID8KNgRjIY79ZD3yQ0oFxmFNh6BgOKeaW6zehBY8wjvPtISBFL8L
I7D6kwWEExMyQgUCDGj+F3RNjC+jD8lifG8/88x0b8//MCYpZkfeRtIvdnGAvZ3nsa4XRzcgyjgd
9glbYcPM8og7Iq1pNMhvXzdFTzCoU0mkEj55bX4KT7UZbEy0fQhnWCTxVA3CHt2gAqW8nrXldO0c
1fKRaV//1DVu0bvVS8cgkbPH+vyOf+hmgkceGcl93IbsJm0dH7ppfR85jqYb2zmlahwxJ8Ct2/l5
AgViEnE4vciabEAlK0UW7Ed90+grBk69aWfkf0HgOWib606dhjOAS5JZJR+uP/AaR2L6rzPCYCBT
a2WG3qx3LrqwPyWuSMkGE/g89h1REi9vfA5ZY6hcjpq1Sh7kiXjkj/adOa9WMlYRXEUXUmS8uxfg
n+b/2Es5E+xDwDnkIgIf+vCc5w/xYPwwjtzkN2E4fnRe1v8qvVZPHLTpi+KNeY9SEjyyVwURmCxn
e4wHIm00WU5xtDojA3zQY9ZZjUpuRETaE/hUdnntYJ3YUrV4T3lvm45Nz6oF32gz8D6AJT8K1Ynq
nvvBATZ1AOKp4Fd0zjkMCbZLnvmWEEkAyMTDb1EDKjpe8unV6j5m6jobmc2ROmZiE4BA0F1T/xH9
HKWeWsF9EQ1LFXN1qe7KWMruSdiYKqXNuakZfwW8xpHWe8rZaJgWpOrNgUoqcM531/8Yb+NrzV5L
OqvbqO6bG2VQ/BzZFvcs86v088U+LB/PQ68otEAEkOCOgqH2mI71I4QdNddb0LCXPOv4kU1Ore6L
7mJs9/e0mYLFsMRg1HTTo928058p5jmQxWb3hpyoOA663a06GuQkb6jxNpftmMlkdoDrM1GSBZpv
Y+BSGovLB1je7N16M1je7QJfCVXkDtYBkwNYej5DjZOdgxd1+FA7CgrGmQgtPZyQRmhelvaKk4c0
BYnCuVpt6UzmYUrIX/kRVC2fObF/tL6sIBTNFcVFxkXOkOQxzVnVizoEs811omXtBtNDgxpBsooK
RZCfGCFjwj8XDWeDTu/LXNEMGJjwE6od8Fr8QomgEtDYbswXkzPkRc//a1qvoSJ6l9HiGG7Aoeug
VmG1cMe7MxDLzZ/X9LtABbXbYXTILEXLYOHgrLZoJon09trrCB32LIxsW9jknL7wJW4h/hDDYtaF
lOzZd9+e5Y1bOcxR3JaOHPbSW2lHrr+bSlroPM+u1YAo0by7x+gHFqO90idFGJbx9r0mhaVsDsRx
CA6FXRCHkSj95nXkT9EvWjgw9kv2bjVypg/GMsk5y7tPv5bbud2Qp8/z6vRq0PQVKta0CcCHlgOG
abmp6hsb6qAUhyePkNi/JNFIjsVIvPOs7z63fygUPrmUx6b1agcw46BfkCcnbgPa5KhWpDpMtaoR
NkIudNmtdfiRGMROjGT0RfeYEfBqfF2TWvLzTdYu6yCt26+iIprWq/vxd/CZyQFcWiGXMxanKTZk
J3kD26Jr1M48KFv0P6EML8+O8FOxJ2aVTeA+cjvQNIk+AU0Bq0Jefnp1ZENoWRko+xYsk123E7LV
B84WoWtAKSeW5JP2oqfOJ8Jt2uKszgQ8eb6U/2OHQZBgKfDo2r/4/JzibPrQmLN/tfFU8wU3gc1+
0SWBwLDmSSL3MJ+09sAimnfwX3bDRn89QlxK/727G6lV3zE1C+raD29CVE1L5M8N0t2oZdnVrqYn
J7oRn/KtOZHLOolffNCi9FgMAQY28xgtF7ehpkaDqW0/Nw7Rvi8I6/sSMVKTzvKcE6jq84sqBknd
iHkvFDzhCs61gRac4J1Am97VJKn6/dVDOzArCR3/wU3jBK8yKSr9DPP4+PGdCM3U0Mbe5iES0MKH
pNOQseHx+SEItFZ5qdBPlLAlUPZWRU5Ayo+Xrqda3zMh5fC6fpLe1bCrKemawXZlt9Fni+NPV4OP
4XrOPPHO7R+3rJgwmjDASg7l3dTxIA+KNWUTO7NdkeL8tD0Zm0CSvsDOvtpHd0TMi9e8+EFrSDWU
kP9Mcbcp4964FBasiSvEUxt9n1j8a8RKbY9VHgfdHaok1C4XvBkXxmKvvLLA9go8GQRXQFSi+hlz
ra5NNMYWIxQNLZVCAGHX1sldp8Sd86t6+mdHxVFSJdqATKdAtZSZOp6/RAKo/JgKrh9HijGxin7w
KZ9F3AWFZYU57SLeHP87ZDK08KSrR4W64SJTIDu6NfTQss1Tu8OF6vdMN2287IQkGBmLLnrXrJst
0B2rQubzd/03mAyxUvUSKi7R/xhRhLKZruE89IpRn7zDE0G9n6DDF4X1cbcv6ExvfkomgXnS0yOx
+wD/UJt956L43n99JIONbQbGmEPJnWHmuvbyrZvD49kPdQzdLtbGTM9N23zz/KyK2ehssVvnLTEG
wuB1e4baFnYMqTzrJHHTpywm2nqQ7xNDwXbu9JQNuSHJjR6BIxZwDwXaJKUxmETryeNFWsc+iybO
7d090Qm9t8/dsJlHHYP8S/m3MVYHAOLblVfJuFVWPpp6gVKslSVlY92yYOPRx5pcYF7tM5XEWO+T
MQQ5A1EYbOZC5RRzjnMCJ7uZGeXi6+ZC4PwyfWehCdJlRVR+oCIHF+oTT+NYvKYxXZ/DvxULfvN3
HY5+sTmimMNW2GAvml3ksb76rRcSGshBKfMcBFCDypNj5I/+x1TTWuLuNjc+mg9I0qJ8ndD4Jxe0
x8P7LS6eMEncHZ/Srj1ZjyUBDrfcAyqoPUMZrjZ6y3mTiuLOA/8YsFobsn9V4uoq9XI3Cl2mrQBD
mbC7CpPSuVcFYDkilx3pevV/DUGS5PO+I8svIzPcBbk8ajOZ1xv7uM6sIzAvDGcTVClO5mXLz0kK
fSaEdbs6D4okgPOz1Lwad1CYmQsb5fOPgMfDuchHRHixGSeIsVsYe6uU1JvNW8lW98oY7Eh/mvcA
++Ob6M580ilOXsc2Ts3G6lpHAhkcDtgDatyfAETyw4IsblVFlJLS6luVcW3GmC1i5c6eTbhMObqu
uDKmZqlaTQ7QUTvLon4jLLP2qHBeLkPJglXFuz3mkYv+T0Pi7CZyAVvna9R16JEzvef93Sb12f4J
EMrreihHfvyG42oE3gerH1VUp+ZtBWnTf2/CzZRFbiWsyB93gp33L/ICM4qFl6kuwvCq9A3Yw2Wu
D2J5QztYd2e4ORUbcWHBoJOk8b70G16VAZR5PfklSli5HArsGq9pIAISv6/k8uhmPySTgk44HVxk
3pLJAlFl3WnrnfJVq/dtDNGbSNxwW8PTMjQocL0vgRX/eUOUJd9q3JAA+hX3LO6/cP0+PRwaKctU
Jw5BIC8zfx0lYXPfFfVZxor6oeOAMu7G4SfmAsHAyM+lnUlk3hgMTyjeuF+XVrqyfX/HqLUWbdFK
w2yveEoNeZih4+xqU1Wia3ukPxjtVUb7xjLxCJY0JxqkUMugXrCqd+jjajrZFahn/XAjX0gdNK2v
N2Nb82epeUl8SHU1wPZPPdrdM8jqBnavaSfTq49mkZn886qsnHtHbCy2XnLjUJ0HOwqSu1AqrDYq
fY7oaKxV/Kkk8UT9om/ixn1R/KLaczDDROHDfs3s0zclXVb4NaqYNbM5SDYJSk9RQ1fUJESmTqUr
yR2wE/LQ1t00/iyTPEtlwI1h5aIiH6JoVdKaL2cawB3BIFBjXLPAO+cCQGS5uOpMaQa5SMa1GSEp
VxoUNViyb+6iG/rQiGPpZd49wUJvKvqJtTriAGV0PtATbqD51muGgFdhGojy9zM6nVb+SVR2ldwz
Dozbq/TKJ/TaNn5KerZeu2I6oL4tk0xjhecDhIaHI0nRrSZrVD8/hvo7cQLDF31q/6wjaKRQZOme
FLB6BiaakfWrBL4AmCrG6l4lpAbr35yNmdW9aj0ICgL4Ykzkb1+QK6Z+mXV5TsDcriO6oIEeFedy
qxajcdU92ws0Rx2H6qIkCG9ebxZDDNuxzB2ETXIAEQaJ2xF7wlUUjjrK4iXwpJsjTFukE2qwP1GZ
PixFqZsMQ3iGiv/1b6F4xjMxVs28/xzI+9V4/G+0lbBlqwGaYjX5jq0jrvKwYe3V8oyI791J5Vej
H3FBYgZYAZjQNgCNmWIrm4t6EEbbHCay9p0e/HQOUG1VWNTSdidJAI82sA/HcSeFm6Rm9nSmOvzr
v3AzbKw4m1yvj5M+Zb9CKX0xRh7WiEYFQTNoBmzLSMmfAPiDovR9pEOwzO7//+ze5kYzUi+1CHav
VUNyrWdAzTQbzNJktJOOsH9zS5aM7i5DSaLLuhPLGepmswdlsL/LNmeq7yPryb454t3tPfIZqUBN
seeTp3hguHuZjhs08WyCvLxmsHsq15tNteD832IxUQpzJ0x+rCHZi7nDts8teAfuK6KWEbyGkrYZ
RbmIHrlIGDos2eMpRDTbaSuONgu6QsXt2FmUol1lgad0yDO7rrV8DvGL+Ir64XLQW5VS03BG1fjZ
v3jfKkC7UtbMxOTuYO22fTN9z6iW4XKoq+mllZjiIY5IvB66DAvxvAc2rUbgOobmM/n8dg5buJdO
b/lhMuXX9Sg1JlBI2buLw5e3SBs52dMU1Srzt/564mkuI1kJDmOJeAE6m4XrNamGRUbHnoWuhkrf
tOLXwHrEgnZM+IuPTi6wK6oZ+OtSQ+wlhBb2AjLO9BPDogmFa8Xgh3fWeSBIBMnPs8jQ9NNtjuNs
WfZrC+XhXFDI26vLMPTvfVNBI8molEhjVyYkoOcLShZDEMwBya3N+G7iiJ27u4GgUVaBxR++1wCt
QQLSLhAZ2gktEnObh2otS2w6CS88Ooi1p8gSfROZK1G/s51yvLjY+fZ4L1YXa2/qK1FM/LD/18au
jcLcYRKal+EuzVlXWvE9Q7g9iOMKaaUEa2kYG8CBgzkPAqPWm9V1U+sovUVoZGD4lgBu2FeeKTLf
CJrh7j+IoUGT1Ouf2NCz6Hi2P+N99xmXpOfJCES4UML5Guq+epnKmYnrkULIcySevO3QZnTpo+0l
COvsb7kRmd9GJNL/IFOeFYDwx+EWOt49qn/zC/cEgBSLopKMqBnDUp1u/Jp+OQEhduEhtvaLSx3X
kZB3U7JOUsDfUpKI8NCoKJKLPprpTkHTvad4BPQOE9MiuVI8IdJchmdjQwTsWFl9AjbqFZsJEtAw
1NoUGn6+BAAEWa+4uk8cx9nN09ykIl42BzKWm+JLL78mu4vMlxKN8kC8FOVu79Dv5sJMxfFLeLzj
CB2YWdJS+LApcOYclGV5z2M0OcUuGs9NVUQiVuNRlVwH/hE8X5Le8Jkq/JueJNcR/DU8hkfWyskm
uxBUj+yGtkf1ka2UUnwr7VkfA0CjjxjcE7hBK33Toyu/vccKS6Y6cRvThLCMJI/qBa1aiFjLrmcJ
8/qatJJ4IGiG9gQm0pXAA3GIvGecEgf/cXn62wVbHNe6brli/kWFLCXulbarLWHc968JqQl5xkY4
40QritCsladsuRxb3QQc1jGfgHaI4RYGim7HYh8gZVWiOjC8tTzYki7KUQNrAMsixRUQ4PhF8KK8
DGqVnDYTZzSWrf4ts/RUj9JDWPNi2RdO53I6jbc+c4UcrA1apODB0LZq+9IsgaFZocVpoQUxnGwv
ucDWLG8C7AHtcq9pXseuMmZANWA0DZSOrF7Li/UVeXAzgh7MdSZmAmob4iBBwaehShX0+g5KAYge
Xw7NKY7V4z2p5c2OOShD6TeNEeOSqGbYQ3xqzuHIhftlLhcvNpGTP55ZJ4lShgEhbmuTzX8SSQf/
G1d7Ul4Ju0Vg7TU6sgK+tqnaFm/gR1MpDZke/7C66kkgXjvAVwL/bQMTVDrLx5PXFfCg4I0zvVAM
uhMten6JCH10Py79bYWONZdOvJzkAF0pSpUMK1/UEsS7nIdFr6T8L1xtIf9wbjgG7gDqSzxcd/B6
9nzITi7gB5XE5Y7NlyzkpIRlYtXaF74p1Ru5+CQLrY9vJKJi0w7Yn3kBUBmTEVtRJKd+dlL4zPbG
uM8jwuer6wKRVQpoimXfzJg25vHEo6X2FPnzrFWMt1vYdPiX/pwMTx2qDfxH33cLyHcnwZibUfkg
5fhck9HPgYQkxoTD8CEGuV9FXBlt5XpzvHSlxUV7qd724xD0AAcMicSV0993SsAy3tDmZaeTs45Y
PaXUsOKiYR5uu5y5OcgB2Xlm2hkQKxU8U6Z5dxR42hwlkOu4HDbZzDuVrt6QlLKD8m5t7UwUO7/o
iySTuiTWySJfHJIZcCTXvTp0P6GdpmJJ8lRSAvCo/aXB7+02LhNjmUZ1FS1GTHlZh0uyuVF410bC
dOOSkChftg5okY9aUP4L22nDVngY1reBNAbi5YjxlLCXt94HIfVxauq2naG4VVGtdiCVnwRb9uff
nvmbRvFt4rlnIiSwh5rslHx35MJ7yTQaW7swUQ5KRtG0KkjDuQa1E/OYobO+0usaKTwuD6ORIk5t
T0J61VKf+zvNn1A9FXQI0fEMTEu4XSy5q2889vnw39X5HUFeS2kqYM99WC5gu7n5XM1WWWJtSu0D
5vrPUOqbWA9eYcccH00m1sNj8u+JS4/ygLI1FJCgFxYAap7MB7o0jo+36ti5QolLJtWtnD+ntBl6
s4Rb3LxNGEz/q5uV9nV32fsUxLVoBiupcvdHMBNMvVMJXQp0OAGr0FGlGhyDOqHQWyPKSsShLlT3
D71criHr+SmGEL1ZUkQ/MGcy3oWsrzfZVacbSvuRjRGUIfewIaqpMwn0WZxSGbpdrQvU7y78wrqz
IDO8bTmyyjQSfbgbHKcgrBozjRx6xCOFvxNIOB41mfdyfKVmXCfTx9gYCokPSQk1m+hCrCp+B7H4
2f6kROBw2zfFb+zZFJLyvvtoC1GgCKGT+Oku0qd9IA/FTtV8QV0B+Yr65xP6pUNgXBgIfWLG/zi8
2Q6VcfFhJIfNeAeIMMwGdUCWTNZ97mz+iAGNLz98Q5ddyCXSGEu93LhYyR/jXddS3y6CDWmiKCsK
3O9m9gUlJLfJT59ttxQB/knwfY0k5sWz3p57YayfOjOCFyhYh/0KgJCNcgpCpwDNC/H92guuo16j
jjxfsUqBsWMw42GrMuLnLtHJ+Mvtmtf1SSB6yKbLlOkuakNzl3PG9oTMg1o2O4gSNPK7w1kyDl36
sWRK+UBnbGov+Faryqn6DCogByk2rK67uet0cZiAbyaV/ngBdIOfUv9zyzE4i4IImOU3yeWAhf0O
+aGFYdVWhf6EOeezlbzVh5C8nBlWbsdhCIO5BW8ifTYFCqRSpzSXa5tzPiIH7EL71xpHHfrLB6u4
zf2jCRyDeGDMbdyYvuBgyxJzYIoJWtbN44i7JomnhI1lsxJVzGt48c/imViJFM3tu5RP6xrZ6JHw
Bw1M/wQGStqdvffIPNwDNaJLruqWLyxsDFsjekaWiq4hzUp7yhVYvcATaasSyn7JOU7IQTXZeWPC
KJGdQiomVRIc3oDjS/A3v5c4J6ib4eHSvUVEpL+OiqyioZykZgQBQipSY5lRZ/173ygYU8GjyQvm
pH/AqQcob8EcSuA7T/MTDlJlq97WD4eWNJGu5fPVirW5ub8o0A9omEDb4XwMWEE7xTfRXIR3xj92
B+i4247xe627rYtdr2VrnSQwzDsK3fzicE/P/igR6ga1KCRfADRMFMMfqHomsbDKpKAQmN2hIUJO
t8JEkfHItd6zbQz4FV2dhc4qnaCkrBtM6Je+vjNxn+l+MflUUjMvdzgZMjKoA4pglpqY57p25O51
CZYLk0Wz5b97gi2XHrhb+Fo5tdTjH7vpvY7pa/Ix2my9gpEvLIEvwncIIf5Wo+IRfzZypu5eAkIH
UoNtEImlq4PAXh3L/+trz2lKZ2/cV9xD2FqOkjWb+MYXsmOXnEDfqOcaDjSlnpey76pIBAlW+xHX
OylsmEyzGsRjb69nsWOykSburJiMY1uA7Z4ycrP0V1/eDpwuLAE46D3TkbZ149c5CLkr5CO+MlXB
z2/OfALsyvjr6w6d5gsEmt5LF30DVO+9syU1v9TMg36TaBGtmyhUO03Y4YKi8sCC0WhpQmYziqaD
5lGd1ZgtSqhl8nnd0wccq+w4igiV3lhbet92Wl4YTAk2fwugZF2hjxUdZpxKynYZYurdBuiW57Bs
e5chI/CTO4wwJf9NCrUH4MQuWU293HgS+8laxl/xWmHQ+VmXnsTbnTYbsUryVHxYDej6TXeEGDh2
3e22lE6ksrLNYPTltMARjxcRT8j+GTuSOJjparrG8ylXUszMWwTQeGcBClnjDP6fzx0DmuvHJJDI
P2/AMOPmuh/WBAGyS9QJwhL7cDKcaIiPmgzm49wefUs3kNlZORmK2KUfxP8Cs5GfLG4cuT3qhyDW
uqlFu2P5bC56jG4d88g1B2JKeXn49nl4Ean5bRL/Y6UJq4pe6lmCQTLKjuyjr1FR9Q/09waVstAR
v0miJ+u4+sxlHMQQJYCIrUakeCyyshNjGV196pS7aW/9SiQaUHAdRCmFxyd0QgHAytbkU0GeEBur
uJatJDMDT5NKiOPo21MCs+sPBEteYLb1c8I0GwMKnXKB6Rm4zzR6HpObKLuk6/lDZIvHuI+qsV5U
LtgKworinbJNv27cd1U96W9UvgenZZYPArzZZag/iJyjiw/YeF6WcwegJXYkC2Arxy50LQjidi8y
6UFOtP4zQ5pBK8SR9MhOcPObxanpJh72H3GvbMPNrExfpiy6x9tOOJICRcFW+HNipV53hParvwOS
F2Z0O934jDE6hA/zABKNXmeQvxaM1M9l9Niaq7aEff1KJvZjP+XoqiSJA0PBLKFz4sGGeKtmsU5e
asTyxKy3cIV1DJ2BpATFS1RtS92iRx+65pb9v3rdZ8Piycf/Mnzj7IH8ta17XBoNjZVS0s5IsCL/
aKcOOkUHai/QqvNevzCYlpCL5U4Joc4wiHN3Fz/PNQIVI7UwMhvhLP91OiLn6rt7DLeEDn06HlCE
80xrmpPkth48/M4zAibtngQQmDP7pDYnIi3djFQ5NNk1sFUe09ECf04iPtlkpq4QpiLrfahOCzDt
9sOVjzxwoSCLrNKMGnQ8mfTsimENPZqbZ+ZuO5FgjPiGi3EeES9M4D/a2XGhKDZ5QtyqHDFfJIBQ
8P6tHXFuE9Ao6fbs8IpDmQ9slLY+vrKpf2vSokg9rABdvLladymORuscMbdLiIb55HdHs68PP4lw
QITmlFUMa/TU1WSmbMDbvL2oCdGTkjcsnEbn3qAe1IgiVVIx3vAJa+/t2VZwFeODpuIwv9dRm8wf
HVXAbXWu5yJGi/5JIkdtEeHmYLKMNWGk0Ng+1XQqYDKgOJkJlq8u/Aua+wQlDMAZi5sScsD8szzn
8Jv4j6YLNxFxxib+9z19VdYKYRJgvtYzmYE0SOdWwlRUOCcvxuxHqM57Blm1uKdY5LGAsJCa9nHM
LO/B44K6kC8EJ5BR5l+wgzidOqkZAYouofa3/wc5F/Zw36Mfxi/JM+T+QNiaDafgd5ZDdB7yGX2G
WQuFPUlUe785JK8ykYUT9aktLqhVqTdgivnbNO3mziiaW+Xg4calKFGuWubmE/Ym18xVGiibpUWp
9bdWclHBgPpkgD02QXnN0kxQ9K/8Xi8tvibIN5vdcHx8gP4+fgKCc/paYg4Kqv1pyuzLw0r0d+nX
4+j+IJg96pw4XLSX8USz81dtPzl1IprE00qmws/jsQD5dJKmd+SmYrHlwIXgyFAPsJLCYCsYUC5k
pl6Kol1Iv5S/G1j4zVhDV9s7BWm1PiJelIHFFn8PLnR4Rig2mZVf8jYAlYKAJBn2fltk5GCKPzIN
V5GuwxBLmRBlIHot6fBvbPJhgPJuBTLnsPNGBXSmm7A6YPjc3mfEs+Y9q5/BPsbk9UiL/LGkZOi7
8V96CQqj22PdHZoQcAO2er4YreqMHWK+Yf4jX75TmlEQnSzYwrFkxmsp7St8hg6kU2lVqT/Jo38K
PTDji+66Ufbd/4JW5U3ZDi2TQkv9ykGyFXk0iSjGpU07N0+3/3dCXBmMBpP+Xw8WgiyfobkBudfG
HMwZFTVUAuN4xaX5OnJgb14beLPI63b9uCwaCfo9oi7bMOqZRUtK08KKIGC5Y34MjW8HWMebhGmv
OVcci2jXChZX19RKFVSarS13FG1Jyf8IZeLtlnfVRyqCIHPvnnavIzn6Un/9+QvYosAGh69UwcOM
gdvri67V/DM9gMfJMbocS/TBuKPgF/LpPr1h31aop7Sn80qajcpUwLagLHQDzMneqEO20V7WLUyT
0vXD3vu3050CAJRraOvRhqV2tITPyFX6GcpQMKv89NW83lODfmG6WQHclSydIKJwqM+D0InYocFZ
d8cn022JMUsoFfs4KQGVmVrfN+81uFNSulw4jRP97zKuPyL6/0Y+3CtjPZWvQnb+OPC/AMCtXD8u
6Rfv4ZbtQSzUKQreaJ12iHQluQB6tnYJIjbqKVQtpclTj1Eq5Q0xsfWF89BtXlJkW5qFEA7lbFdO
iVzpJnZ8h8X3aNwDzm0RtM0aSWgYEPN6QQ05gSCvF36vcl6Ysb1Zo5eNV4htHI8D4oJwNIIGKqzC
ZLx9eUu2XynWS1167c/Qyaqo3OvEzMTzfy7PbUW3pgy4LU3Tq6TraXn0DLmFGLaQcpXuk+PFqOWv
vtzegtKPnvbSdsluuLHLHBh4p2lS5oYwoqGGrj1dyxcDr3jaAUZF8nqM3EDj15e0jBM8lfFaPQGO
BNLgrSauD+WLtn9uWwIrwEeVxYfA0MLBNycSpe3fBUmsCokHjODMTMbL+byoyxRjLSAY6i7IGFK8
bALqjtqQ9jU03RTed3H7Kb6uy/7UzdKUFcDI/uZlyD9fbvsOrexLB1mqDJQ3geE4noiQad69Xahl
hz8jezo1TVfXZH/1+jZ253x3ydmtD2oR+QMISmpmxMcLu8QPDbalPF6B9y0eS+SPtVNdChIKzHrD
tWfC49/gtxi1r48VtWEgHyPc8EoQHA/4CQVnoz2xxJVnXDYN8Eq8J6/AjnkG9YKfzPSt6WYsz2E0
rPkRqdKyqUyZEY4ak96ItCzj1npwMjMXZoCnAMq5rZL1PqHS743XDFc/noa8Fo2dbx/CLkfPu0dD
Yxl7lWFBbsIEThqdU7Bqd8kMlCunHGyCJLyvBf/o9Csr0vLRTzt8IvIgTZvu2rPImNXxoJurq8fe
EAyHWqLMcy3Cnqf5AplaP5CISRvEZDOcgXIM5vUAXaS0YQz6wqWfbKTpVhsb1KGCpUW9UVHcGMzJ
oqcYBVrrGSPy4ReWPoxhJWKfXLDOH/p2eTDjOwxdHEWbTNXRsEdesBOgi4uxl2deAkZN18uUhdEL
4dhqtoRdZB2gSfwkpNBkyhDUQ4MJrOb1FAQycSFhUtMLkCkVA6w5FvXsmJ4RddKP/68rFpLvRjK6
3ysq/cDdL2Px57p65nTaDqBCUQmfWgtO1BOCzqA5LHhe561yBOxgJyxxqCRLTDlyv9zWIpcfa1Lz
LsRrtsv+Rnt5DzpCDZTkq6QB5zNKcdx0yDyHt9YJ3hXSdS59tk5yzQfUrE52j+uD2eoyAq67V1OH
0Po3MZ4j1tIb0Kjh8dt83BydZr3R3S3wAU5NpDV8l5llFOr0t6oktOyryfBYaNWCeXeHttepTSxR
S3uf8JfpR50LzNG9fo6aHtsAtjZuyduhDvXmKVbzeFfAjY2uXvN3laUWLfyOHwS/OqHmp02LaAq1
KK2mMVV4WBssmz7qyzarq+OIzsSM56QVKEZM80aRa+WUpd3L8WSqtxSPTGydMig31N3tgQvi5OnH
fNdJMkwjZJZO7oplMQOHJ/p7jQ3QmPwTPgKpJ5PdbQAmEFAJ2w3ZTYUpXwsB4ilsFdV7ee1AjYsW
csv3b9fWJL9vQ0nQ/FOb6YUAv7nSdl4wya/UKs83CoJCL8DMiNCuHYaBqcuZm+gUi8uvMmQ3nvEc
rXpFOpT1WdHVx4CmFA28yjcfZQL7qsbQDQWK8DqdMLAMAOlKvRWuRFXn16DYqtsuHZ3XuiebEOEA
jVdJutQuM0qn2FoC4Z2uvYd7Kx+63u2KOJd/uXxgWvMos+MLR7dWMchMOGW1BVCn7TJGHEv3WNu+
50qeG+zZaw48eobtaszOyexAq+cswAj4GUjqW+M3jJHci3VRxJu5DvegPOx5jI4yau9FLvKeYfMd
3xHZyk3XFfDbQB0fNQ8aGfgigt35iJuw5fMzBps2ZnJH7s12brO7WoUwVnsb7RDnjXlcODVCfzOp
e5FiEzKDx+W1ksozoFiw4pI0TXp+t8B8wtwo+RfKH9n3s25/ALZCE2pDp4cQGEshdu99iEDtwCBd
g0Q6D7X4zL83eE6IMePkCaeuR9NYpVwQRIweB1YLEUzFWGnrFC2QRD3Jir7vwuzb580eQ+d5goTs
EfKVhvfephtKkvDYVN4P6rFlKtBIibfrYAP2H8ZvLkoK/imAId9GFdpoLfxRdXLn+RKOPiGUBMLq
Of2sdm8IiMoq/kbr6G8ipk0oCr79DiN9ZKwp2HrBSgHDdFRC+6i+stavubVx/keoCQ4UtvTpS3Gc
MIC5yMBRuMUXXt+JmocRKHhEx4Su6kgeWvC8xHqwgK/MXmw/pM7JG8WsA6pNUXelNntB6RWGgsM2
W0Ko6N5dNLSXnb/HyKDhDrhxoBv69rhjSxUiYTGutZ/N4zELWIVV7aJP6Un7W1fVN6xFB2MAZQoM
wpe2fNLpp0hJOVkR3tnDjUDVmrSobisfzvacxDgGOqpJjk39pcBd3GvCOPtmcMjND58zLDZDsD/G
EBbAwE0K7C8KrQ99jCmyGvCZJjQ5gLxTj6C/eEnMZJUMNeUvvJ6hbf0ZWYaE5oI9i0Z/hZrHwR8o
ZFH+EfRGxuDZH4noLMJgu/Ptv+KqwTWRD6VMYnK9k88xQPD4JS5y/Giil1Y4cB10tZpDdhbfwpXV
rqdtmc9+8HELNcc3BbS+RcFOdaAbHV6xMAJmf01vzz7HQrKnx2aPtFE1YxYfT0ANoVmWDRS/aZCw
NZawSSt88XGwlVtLuWV7/I9/KuaJsRP/0Xo4y+XV0ILwIdNphxzWEqFc2mwbPSYBubhLpTBQHAu5
uApnXiV4cqpYL/U0b14BO8LdX50wZZF78N8JW61Za14Cr2JKCiaZCphNx5FB+os4degXyWSxehHd
EJERC85gGcNs6vyOx2jZSMlCNpArH/dY9FSfiBdUICim9x8aJ8ngTBQCfZkY+lFoOdSsjDW4CMAQ
dLoMGpWnOF1UUvmU8S7uHrPHuXkgfnl3gOuRThJJNymQSGRKWYuHhwzuifc9Njki/nIgUV8moCqI
WVf6eZwmXlTmyjFZ2lULu1aJ5i3g8F+EF+pD0pr0NU//XVWKdu/qhG3QxW9dV0T2B+j59DeWTP2n
FOftc7T7XUbsjm4C+QE0GF1ApmO/N79/8z5bmx9Bmuyr3foFt13k+5ogHFIJhkUfD820fCgFNY8Q
gVkbk7fVudYkK8eOtC0VK1RWnxhn3UWlOs2ijyrPL3SpO/wA+FOeJVxO7uVSMSOMDmnVL0AnIyne
on6Tx4gl2hYHVOmeK4vka8XxFxJQ+dtBgSxd7NMEDghTvztQL47FNXKUIwdUWWW/lV5vFuO9pR3p
BDLCqbw0nyWyF3L+tQ39eUKSUgYNviAYb1vFQDu48UnJSQLHxkgezxeuQQZcKBMWObFZ2oRATr5D
stLjrMDinyyWcZ/LBmsbyYDjFE3WUToX5T6938ksD9/YuaJ8DaYE5Z2OFj2/7Y9EAjbWFJRyetwl
tTgE6LDnAqsFF3pGNzI3e4ZE0CO2x9lO9LcB2b5oK69OSENyF6s1F1G+qsIVYjQBX6x8PXfCd/J1
yF/5I2vQwj5IipR8GZiLteFK2R/v57mAC5dePAyIb5mNoq7M2WINmVEPsJLh/6L/j40XHkGXqGKW
bGd6zepBOJ1I/5Ga5ClJ8iqqV8BLwi3EloOddErGTbKWl1UYkfK26PY/SRZmQo1u8EObDLTEawUm
8ThUYCDeNZaCdoiOLthjTV2sBf7zdetX+FMu0Zx6O30cAiv7XwgKiJ4OsqWR60iZeevB9JoceUBq
5NnaZ/fegozic03w2+ajQm2dfxkYC4vlya2C3itxqUPCo4AwVM9s8bz7UDCRM7xuH8RnVLr2IQYS
N/O/NxeGrIeR6DlOeCIOcOTfcQH9YzXdUcc0O+uzpQGy3hvXeCI7II80dQ6fGJ9i2X/UUuMfn5bk
cYMeqdzIuwq3TTnNvDFOW1BgMbnkLkDCEOzjSshVYvDZdyJFKjhnRL+z4cC43JAFleC/XlD+PXBh
sGiZPdD0HJsbaw/eTKllvNTMiMtSfPj1gGWf3judbjmezwCRpmq0Kpx44kRPzVOnpT7Sj/adqrA0
TZFt8QDbcEWZRmJcb2DSCLX8hvHbfszZwwZfcPixSDuYDgb89ecAt7djj1fOmrvNJZzgEsQqwup1
KnxSoIfSMHLoB1b8km0uGtt+1JtRsVxoywNbSB0lg7I/Gw774juOxkFFXfYtMkHtsIAX7o27M/Vi
wxTeO3Mcim3ppCb6YAuCj0TxuTR5vDe8c6BaaW0f+KYu3RF/7Hin/fQmExrh2gQFgoD8R9JAA79k
0hbAWGWGpIq7a/m6/maujlUrGbFIfm/+XcbleaSjYXxcjzCN8Qy4ToIjnm/tuGW1TbHu4P7oh0ow
gqc61bfKs2NWQewNcthgQjRMXfi/sOaWiHEKMpQrDaDxKyNt9JtqLfHHQhCbTDyrHj34hxbf/L08
ZAP8uKX4BWYXqG3mngDduoCLRfY0YvsvN1NrZ7v3jbYJCu3aRgP3cgMsocPgTCMBlAcTeTlyfSQx
kQt5A0Fhdmpah6wzC2sG+hcwC6mAMCjYjvfmROwoMFIy2RQ9HpAy3YcMTXnkp8wMcg+lPNyV8XOl
vq+dhkWDuJRKRNJqx0pFr+ml723TyYlnVhzrpZVfbs5/LTsChuNhkGYDmv2Pu/ZSuc4B6DsM4BIe
FkQvfwrgm8b8VH5z03+b6wOzVXnkBlu0ybXs37FFNiaNS5Eh9UxJGAShVJddLtvZdRCvRBI7n5Jf
p3FSovkZI3jQAXww6SCw7XPjvkWKcmlQP4q/Js9d7yawO8GTTl4t1YPq6PU5K+BSVuqwiBWUsrss
ZGp2Xvow3BNVGqSIkAEuRCqXmcaR3ggdiFThbqZK9exQv2JEoifizJ4QOfOB6WeSVLiW8YdV4Z62
5nysMcBLtcEnZnsP7cBJ3xCbYZbgpRmJ/7BtuxP/uGfb2Y22fF6uiwY3aZkvtY0CQ16dhqSpdtbh
H2pCeAeiGazB7nXMYZJLwo7OLYuWMrg1DepkFoep7xcx3gK1zO9YhAEopeYQM8CziZDKZ/BHGbl/
UH+dpn3pPxgYn/k+AYZBFQWeysYIuHHQlOIW94vRpP1fNjeAaLt7Fddh8GaaR2FIyrITJNSWj6tQ
J8ak18IdP9LiUSLGHbnKkbep1xPb3x4kEf4PvnnmaH8nJKYBhwcUhBGH81N6talRoedIG5IdkZiF
TF0/bWhur3tpREn0Icx/wzHaxKbKNjT79r3z0sECKTfbWmBOmt6v6/0i0bXFuKPMAUT9BN3zOdcF
M6tbSrahOzoc9TO8BxQzH03+Pl5Kn+q2C5zOeNcuRoi0pfYO3AuToww9T8ZfhFlJTcIGvU6CuNKZ
Wy6D5zYVaPGt0lcjK+X0UE6X9qYUxB0Wg9+Lr4P0gSJyd/wJa9KGP0sFE3l2j4FLpXKy5thk6Ule
gcI7bXfRKjzkdakV875BC97IOdaR+xdc4mr5TtUiKGrVXlAM9CBtUzAR8NSZBjZbTSyldu3qa5qG
iDGOH2mRUCoQpJFx5HDlSIyUyQXdRPgOZJ9kaBUAnv1UhsChAZGSurHMX7cIYtynIPulBu+Zr24P
XleJsBItG5Qhlk+XyWb+0fdEqaXTbl9URJMr3SjmWPmIJekW9Eh5T5MZP6IcV//jJpDX7v+kaE7h
4Z0qDtd/ZCIoudXZMm8GRtMVNeXnIAbvo2ezEzZti6bi20QrZ5QDtSpLiP1fC3FYYB92lPi28bhW
SGvOanlSa9tTzlfJAqv4aLMgcDUGTFWwqMKoyxTi+du1tepP0Fz8Wh6au2zF/x1FJFuMNYmHV1WX
UGeV++FOGsAbFkIz2jJ9jtLuoAcSW3AQ2wxnU9kptjexv3grbEirGMTtaqBwEReOC26rYupGD82u
jYWYrRwq0gCRu2FPmapKZcwahpMOO0K6+FNCyO5HKHaXW44xsusso/v49UzY+RBuYCw49DpFs6PF
59zWUzExeqQSu1p1FqEC9NAm67AnJ+Yfv21oKef13pKZahODdC7WjVcAVBmy4hAelOK8EQBwHwSl
i2kCY6St87E5pC5aYNWLdME6xGNFuxPcOhTth4IhAkDRDbWWu0WPgKR8tTn2Tw6qmjXFBwMDwWET
/D5ZZGbieXJqaAq1+ifZlpOQRYvu//Llhz6lmrjZiOzVnx8PShKRcF8/uFxkcnp53FqpUuisiQsK
LasAyDdENAkv35lY810PJA02SKjtpGLhk7zJHslxcQMpjOQK981wQhClyZNqXBpoRG7FpqPMSt0D
Y1z1vcOOx+DRMg2iTLBwoyYRWsZ3WdCYpTKvEIfUVjFSifdfZLk13exjM35vEmKlg8tWARhUOyqj
RGRh1gnPjFr7YS5iI+Yd2J1wVjVw6vdcFXUhXLXBmZkN8Po2oIeG2BjBe3b4GIdtNlgLe+XAv9k3
HUuv/upF1XoHSuXsWqxEyc3u6jhZALanmDxdH+1GhhbzI3NmRpUVDkYVjp6kLpQ0cM6TPWy5Q6Om
Oi5U6E/n6IqsCdjZtS9SaiAyk9Q+WhcKT9+O4a5MmozgJ8ZkEL0Zu9FJk76FIz01kF1h2gkinJWj
BvsjyKMLF1XaZns+irk30Tccj2VBx8BwS04N0U21cUcHT4AtjqVNx5sFmk7plgpG/Nt0LwQmzFVg
pRSvym2WLe87o12L45yuh6nSeDtPU4SEMgHQsFz3UIVGJhkH4fqLKM5v33ZDWSMKiJ37wgxh+FUe
Bw+TlxD3Fk1+nR0eS/Ei68YSJ9yG5dUdc83SC8FWQBKxxl9uXeimC9TzSwR7bu6KzQVeBAj64LSt
lK9/MYzSFd9igbzJGZy3ia5e2y4IV9/jPHla9vAc6GTWLzpdT4geNTBlbNZJZ+SFvyQ1+zZmkha1
10h0PtIgiIqqM5Ora02sQNr+xYMcWF7dXvRj0mSzn92CQrujCXfIN1TwaHYVmpxSut0kcaqzNsAK
bZ0d/yiUA8puUvtxDx5zPIX8HzXMTOx365TS7Tv4CLN5pOwzeh6kx489Ml6EfgJjfmmW3B359XNq
O5Qy3neaLyJoiq2RGhMz4bl4beQxXuiz/xpaQG3v7h+hdCXTjeZ4nlB6GzTkfLt0nhzDI9Ftt90N
1X3xsYD+qHSdZLMpezBtEVPA8m1/JmEDl5xHEnA427C+fDdiFOyNf8/sYepJlv1gMqQ4D9F/AGzY
5HxmMXZcy5E9iIqLgvE+SzZ/4bcyHlqDwuwo1v53JNYzjQfGkQOf0oqbkszFPCALuFrNI2SHKmu5
aaTWDh1wJs+tWawYaj1DWHlZ9QAkRFBINDj1X+ICJwsuR/fpDZsqC3xtAlglTPiiy+hcFK4yMXVf
vyIPJnd8DpMRFG/zRRT/xIzRnbmay2ZAWm+dhhND6QMTt5loVBBJviHT4LR9tschbNXpONbNbsA8
YaEtfd/3SB3B1LrMpm6IHb0dLV51VU+rIroX8kMUl6ti4K/20eIYOS1yC6puCPWk0Czd+JFegW18
tcmgXmhtzyrmjy4IhZ7va+FnMJYexnOwR7yKEfklwv/6Bim0LnMeRXqBsYk4W+JbJYShaRJXJZeV
AGOTSWzX4cCckpJr0oAjaWSi397hL9pfGtJAabReS2fHsoxeyj1LBKmQV8QiSvAM8Wsuhgb3R12h
Axt6yZ0DBVjJRallWgaNa/bCXxj1OO+GDIBA2cR5/ClR6zjNC/ww2FmgEz+vLlDWPfVNI2B33EeF
rZrn5XN6QBv5Mnb2Jdz3fdJsmhWOL9PB4+lUe2pmbiRYwW21BPOtBanKhA6/0zwvG/WPpoghyQ+g
JzSUJeORUOpu2FbzXSm23T2GOkVwmGU1u39e+BFGelwCrWS8CCbRIEbfba6iHZ4LIkQQaF5uiOev
HK170tZqGE+AAyv9Ic1Pc6vcCy0fEIjwmGiKk5DxINtkTrmKSSAAx72eL7f4I3GoPHt7ZERrEjZ6
ICLeQBXBnwu4D7kg/oZjfhNUDjGpHzcM2RyJTaSK8sVtjvlO2BFz1OtdjXC3D8vuix7E4LwkFgps
IVZdaOGUv7ETEUG2yKMMkUEOXwoi1rN3wAxrHg6G2Ml6ortrMBjB0yPJ2HnMQ8QgyYSs4F1WG1ND
N7+XV+OnXZzX1xV152QaeJJyQeyEPTLFA2vOnDnYLxgrhHq8VWZNN6aN/9Xcfkb1Ic2MGt3DdbOA
kRgs7YMCzhLT/I5pMnwMKVkeGtcO8nnN37t90Rb24agR0CMkPpFeq6RFlgGI/kgL9k21EZtJbQWe
XiXnuRZZEsL+a17q+uUflK7zs+3a+0u0rWQ019IGUg8oTR3z8H95ssiE5Y5osqz1MbZoD2qsuEK7
5mAvZ42mQsWiaM4XznmCZAyklZ+anSmwtA5tBAHUzXd92Y97DopNP301q7+IsQ2t3WrCsZrciyGM
GQCzoE5m2d8fD7wJryBavBAHHA6nkSb+a3mevgglBw4XQ5YK9zPsQURRFQFkWoqQLjrUzFwjvKRv
AceP94XC8bMGaSB2XpDyGLVnS87ld2Z0qKa57soULYguyS8C5v/dR8BZP/3fsqp/vwm8+8+nmLej
ofTpmIAmMEfX6vQvkjwwXB8/ZRmcrMszHw1aMOy5YL7lIICJ/W8qDozYSfFM9yWzcx3h92+LgTHy
4VA4seBE1GCVHZamP9pJfOVSONiATemQwRjWS10qOPbmrrYO/VRszMf9zTL7G/VMfoDHyyKtB3g6
NP+CjqPqauFdEzfuoEQ1dPyvOyu+dMOzshmkleQEk2oonzN+PvV2iVbvRvxagMGZuGCwcBMJ6rIh
/2JI8b1wcEz5RJEGOKKA01Wn3u14t/89bSRf1tOrTWxfcsvYibzdTKNhdUZE+puyd6eDCtr2WelY
6Gwgppvjz1dmFeV1jOmozVMQMfMwxA6VkLwZBsS4DSfU/iJu3yR8+W6tDULpMpkUOaS/7+ZxMwKK
znmDlYCwdG9rdpKmRAXb+RpcoOrgY0gBpk37wxptWeOltjkIM7lnt/87JICdCbo5EJL+PqLgG+mE
23PYJNv9/aRg6KwEw9hTRyDDwD0GvtX8Si/PVRq9cjPnYCeUPJa03rFxUkKKyQV/ZU40HIAwYJgG
ejFoUPXZJGKO01xyqSnTZb4+7smLZ32w7ge8NqTpFnwG9wMrUGMp9iKIupvWEuNtPLvWGExkkccK
xND6Ig7Tr3Qe61FzRs0i7Aqf/XJ5XVSbZ5g5jdSsOhv8zxuKtJY4iTt/bhX4hmp2J2hllOfpaq02
fre/v/1TS3DlYrvg2A7z4OXsGCrX918+PSiTQQFW6QYuiIBHw95Qi0YIO91SKDBWxcxeEIpBKsJj
ESFdP5IV8R31VnMeIjCVuciE9WTg1yzok+deAQMYNmvlbvuxcm69insrD67Aw0rsNi4RX4lmhYdy
MA+0HCSr4Lz+whTml1KixJwCFipTE2wJRuG0OTKAUuVji12AuyFQ5catYwL9rLf306sWrm5mlzgS
nWU9haY0LypmrzIa7cF4cUmF/HuamQ5aVme/R1xtREWopEjVPHwUcCESSFRBdAVQt9xunGsVO5qo
pPwwzB/5LsAVmWtfO5gH8MlLH8PkRiSf6+GJOcDlTQeEag4ZFp7n/TfZmhiOvSFp5uGCLhmRfOKh
oEaj1L3JC2C0cNHfxIHand670RfD2sR0NcPhshCQgCCekI1dkgArXOqJBu2pTUKpYh7nE87gL31K
nQ2W7XWuelXAcIj+Gc5D3SaPPM5zw8rk1ukxYZYjOShmI/NkmDA3QLUZDxoNS41U4nHT546NtnqV
vH2ewJMG+a5KsVIlyImjEUcxTDweWEvFIBnbO67caB0r3QCCSvPQq0i44T/kw0gvX2K4HdWZC+MC
qNEWJSjLUhLqTMf9N3Sov1KMb2Hd+9jJLQpnoDfj6NqMktQ5qu6Xt8Cm9IuxwGnuY0mEVV/35Kgk
EfgWXtqshjPcDBzugqAiiBEvRCtaHd0L8233PrkjU6dP4X7DjhJoKVlLKqvY6pCBcEsWrhoHKd60
84erwuQiPB5PNLX+TpM8ejGhxMfpKBoFoDlQ+ImkNt3qH1xlEHy23zjH+74i7WfYpVq47zJQQfI+
eXRkWtaEnyzrxORa7kR6dbU63XVLkQhTlTZUfAcNDzF2PMMQTCs0FNI6fnMQsJhWVs3XZ1l73cSW
xEz5q49tglP4nNTKjyuvOSc6Ybte9rZQBL6kLl5QcM6zMMohjP+dCL40iVcKcMezQztyFrwuawBw
LnS4Yp5ayXwycUTegFhXdKbH9kzTUiV2uLAWjiBV5UWSA/+kLUbcCGs6meAcjQN5QrdEmFnx4r92
8tdz3HhZ9CHbz/NYUiMVgeLvnrGQ0JwxxRglHvgq2c0foaotzA8rzif4oefKBwr3N9nbrC6mQKJc
oxVYjc3qm5/G4MzoNBhOrY5xEhQHKQdqa7Ga0ZdsSBCrJixpOVawqwp1rN1FFRQGA4J/bMda4rXi
+sS0bl1/6u4RGoABfY6YJ8zd9lGNJR/qLeZNomyMKxOx9CRW1J/0h/lzVcUoZsZXf0W+rZBokDU2
Iw105Qeh2vPDSFFNXHjtRgaFtkaBftQxuaOpOSA5Ll/U83VGUhuttLixiCeTVSmLTD3zUomNX7in
vO+xUrbIZrHc/iWKrZET1H83DERSyPnQUhQwDdVE5n4jhTjDgEiA4oMAMf1AUNH4Oufkw6nGciVg
U5HLuuwUafGznvEFhkQNwYdZ4eq/YG1KEW03AQhOKEva4dq9o+S0EMFrF47ZwOXVTaCodxJq90Xt
Hs3DUAdmVPVC/VwdNLAtrUAJjnagPSW/lI8hlNJ7tAYRshwc/+Zk86U6ClahunSgDVxgy26+jQG1
Jp34f1wLNDU7pwVOvrQULMyILXGWhruVeqRfo/W5ALcTf8muKO+p2q2iHPVWS6iynBDBb2yJzGmK
aCZg3t2pk9sASzYrbrPB+pby4Qmx7xRm+ouf6YgEfY1GYx6PsxeRlEkPVC2fOpLPpQ8iL7KUzuAa
YnBQiWL7UUzMWebP0JIHenyEtWiv4VyGYnn4AG8g2RWobA4usDjo6qQnkzzQoRcSkhnb3qK6NHZ3
NWYQlg6t00eOkxMD/RKiXxDGRGQoKmlzlqOeLhaiUGVBwNpBAhz3X8kJ1iHmSntFPRJ+ZsYaMOGl
Qgjq9Clw0vjyHaoL1eEE1cjyRu84B+nPSxCymno8D7RZ/LUIQT9ILroVfsB6/LHf4Y9pTu8BVYcY
lnNKT1JisKE4kq+ivC8i65VJIC+UxeLyE6s0a7WKWyMj6CuYnh5IyfJ3uvno3jeFDiUZUBVqRTrd
hFqm35LkV1Z+lN/ezMoigieWwekn4453AF924uMhc1FESDfefbd+mOeyW8YwaLRlbDhAv1t6fJHG
cXDThKJiqyaWstcp+TtmchHd6e3V+0x0GBVVfkCNJfjLnZCnLIkkFQS6wdDPtRfLlErmWZoix2V1
UNCnDNLX+CQwq6vi/Lh2xXC9uJRFsGK7iyy+3nyDLESSd1PCbytovWe6LfJoUEB2NR0IlEgcDCOa
h9AlZGhkrhoG2oq/gLHMSkQc73onswR+RyM5mROkVv2S/3/9hkSNmaXrohOCRT2Cc6v5YGRSKmoV
c7iDxeeuHfhx9lvQAPdIyxokhOF0yGqiIb8a62H5vgsoWTPMEuc8edQMkz+BboFU20LDHfXbTVGJ
Rz4/1q1Vnwc2vhguExmN1n9fI/bav6yG1yIFbzK03I6rOALVRdA8o5vltcbo7e/yVMKow0fwqzbH
ZYw8ujz9TGAyy7y7XfPX6mhxSX/3BewCOEH863HQKKSG9jn9H9R6A3pw05sba80hY4caqr9L3xnv
Iup7vV9IX0QB5Pfh3TnAHXcKNUBbk8NZMCEnxbk/pV0NBWNuqjwvr0uc3KetRYWKNdUY91N/tzW/
CYQfU1XJS7oFnKj8hyfD+o28edV2+hyUbX+DL8XxIz/HpNrIbVry1xspCHdh8amEEEqY380nwUF4
ZwBqsTi7NCL6umL9TETXlyS+5JhCOAsKQLoyQwhsw1IgVjJabqniGNYHk3S0EtWDENfygeTG0gda
fQq4QbCHucuuQByo5GxxvrTmt+khJkFUG0m2DSheBXzFghWd8ZV8/G/U1uP8tMu+H6r8c6rs+KGJ
E/uy6lxIb3evfmw4XTpwirTRAMKsc8QjdkemNzNp/voPJM7qFMUbjzC1zUHaMrTQbU97w0YoiKij
ycy/31QPF7X5f3tsXRXjht2IZPtJKpKVK06LAWhMef2GY0thqwqP1BezNSxywZXs4UsFaWupePmx
9BSrFayCGkmKwf8qf0ZMwBccXflOEXBEvGcSYSajZXLtvRgqlvaX6Om839SOlxgF+pIe2sFZs1w8
DVNmdYJA7JduOzYdekO2v5rxQ9Y/D1ZF7CxTijsMsxyt14vUpCbpo+fk6U27XQpZeSfH4i8xKqkS
SWsBitWgbtXdtms7lxp/523MqLyTPk0pIP4soNO11Kuh9vBay14o6o/Lk4CGCvEPK2GgZIxvfbWP
AQbX+E/tV2D/0OQzNRH2ZCIY3pnxVsspDqrQ7OrSQEPXaxeamcN8MU7auUmxwe09yd/91NdtSEjK
y3ouzyDUyR+xo0kn3i5n3YUzy51y1eQyJHa6jDVsOI343VDMFEHiKdU713FhNMt8L5UfTN3I5IME
pdIpyApsMQhA+7CZZMY1caBNM4YuoecpUxYML7XF1O+/2E1JKb+sl9VPhETAzx1bA0TkW23hnRiI
RvJGLDlI75vcLvVtL4QqLvz3kjbZR1kabteVkUcoicTBgPzb0nm27hMAJ22Eirq3Zw2j99SfuPgG
mZtGik9YuJPU09XBJGuvby9UvJGDuQaEHjomcEmZ/N+v2yCzweP8hZ7ApQ3disc+wjjp3p3b0Y6x
vGxRP62hXPOUvwzoxLAaTbFNusuq8a5Z01LpKpzLzCea8gsfZ06/h9wkrAD2oAvMrNjtnIfyMapH
PzgU4Ki0MK5lBBltF5MMxAXB/46ZnOfhY7Pe1bo4Nz6f208pfkTeJgrXm1FPIWegM8+cvXF+TXVj
+sKDteUPKcVrWobMFhbBZmCDREXTiOsO0UNUv/CytYinOq8gPOKukHWT90PLU2+L9A20KDWuzMc5
hVJ1hA6EzG1bH0aSzvLZzrpx5Db7GoVRgf0KQ1m4PlRUWmXGYkXBLXyGtv4Z0UBXwCHJ7NA4GIzA
zcCIuURLyz7VfTerYtZsHmvuRIZyXNeRd3yP+vS/uOOdXVSAqHXv6Cwf2C6GZYeK91SZK4yiK4P7
IwOIXdoDQWLwq4r1t+C8Xx9dFGJEMn7SmLqPXYy0k9cIF12lXkkgjzdu3rJ2gw/cEUXp7lL2HfDn
3M3FOJ1/C9sCAmFhG+etaOnsy6fhu6j96o7QbKdCcEpbKvlcbRL26hnnzYhHkAuMVH8uvgVjlI28
CLjAPdfpSkxcyGa/NnEjHjhrmG6HRb/t7Boy7onP+23kxvZrxWIxvQin9o0WQn1K3gVCNUB9h/0T
TfCiAu17S+7mKJgPEZd9wldcksLQqCmA0UeKY5J1+2tvLTU3FUS08nwozk/1cmZP4O76053nIMbg
hdOHVjW3oD3L/er77LpLAOeyYdeSYDj4qGsLxbvHTLejYjeWZAS9VZvDBIcgDvhOejZ+mC7BMtwt
9p/beBuYGbbUMXf23ZzL2Wb3ez8T7/k1pDrAx6AFI4mWAb5ji16BDdWGqAAPa9h3yD5EYVwnzuTX
tCtIFOffZIj1bX9+3zH/OYjxKKb2yucZWNS9Sk/MgXKjjA9IRWXlYzdMBRc9ldOphw0Lw+Y6vQ6c
P4hqiI4WdsUKZPWuE/kVWsfvr1DbKr3RVmnh2/BYQAu5hMOKlF1QoOgUtSVKCN8cLpEPyigf1KZh
OqWsDuiok3YY9BYyERm87x3xSjo4olMCF5e1FxCQ59U9a0ZVqyvnvj7p5cVD0BywB4cptCtbS0d7
jk2Kz4bOUD21fzRt1w884NUdtjxFi68V2/iBa0Wj0rOUF4GZyBjp99PrCRAqCA/PbT/Anq2o9ZXN
e3DH4BfEsMhNCWmY9pO6I/Ds1nkWF0cRGe1+Kb2OmZGhhzil8kjlIIykFQTLPnle1j9A3zt1trSt
hNc4op2Up5HF/Bw8xodhCul6t3Qok5w3t+1E4C5GVt1Ac0C1nRDwZeuYYeJj0wtw3P90xD5iRUHf
t6BraDuWaVQG9HGMyvhESl/I992LVUaiNGQPXNUGmlkcCPUoPdFdxaqsuYsvQGgvnr2tqmWSy32U
jPO0T3w6HBZOyXwuX/c6nX28Une3Xtjcy42nD+zWArIl8iERbacj6EFrddYaVWDHgm/hciZX9ob8
4AdX0pjCT/UBK71iQWJpi60cJsD5G8rJJoBAUIqHQ6iHtLoSGUuxiQpGv/7Hba7PPuWhd+uMCIeA
RvvEtb0Dzo0sGgNRjAsG4/XHpRrDOhAcZJ/suZokPFUuzF+c3X8XmVReEcbTsPt4aJCInp5Jlo7O
+syc+e3jCZ9dztVx4gkes1mH2NGb14isA63/wMXXTKqbR5dnV+kcnAzKOkGIP4a3kbCoDyOYwSGK
/31j9+dPkct+c2Gyln/nMShhwm4G2MjnlFyxI9jDc4fDyUZul6e8Ea5x8r7NYTnk8sP6sctqETRI
z4Ep0rp6L169QKjASVEpmbwL8MCy9zPVNWeM3mJ9nvCnY7nMDr6joXETVoYSpNn5pJ7s4OujZcwQ
YN+eTJXc7+zJopjWCEMxoMbW2tC4NilCo+ttDOp+GvYDEICZ0B/l+YVp/mced4U7ItBfoW85a838
HnCtIgXjz6mP+KyHCrGHYx2NbF4JMyWm/GVTKIB2qno3GqQcTv3zUytXnVuNZF7bvQrA2i+zNFgh
FFkKUPIoOeWHIFpGXoi3YUlbF76USWJjdVP/9DRMPcVcnmfSH/UU4sAF7p0e5+9yeCEiqmcvQFnq
ZgN5VLN1gSvlCZ6gmg0FVYiM0WoEVwiGUKSRxefVsjHJ3ZnjucpGILR1PuujpFF51uwA3PgopKqo
zgZJfFWl41uOiaoWheGjN4lKQDkhejfQPw62cOJpsCLX6uRFXASNnG6vsTVI2d0QY0XgLCs4WsgF
13X559zX3EbGrkvfsIVP2HfntfuHNQirHp17FUdiW0XnJbzc1aahUHSeRSzOx5CE7AwgUfhXftP7
ZvSjzkDfp+RsWRItVVW/moi9LnjkF9NkVBe3EGa/abaaRXYCsMZgzqcyD4WiMchQc9jHdClbVy/e
QUHZuc0elzTTIHxJMo398HQWxQQwdl/1wd9PcoCuecOBhUClXsWJgOT5xH1F7Wt7b4o1tYzmfcgu
I94qTeJw+Bnzgy5Zqx3ENhjDLlLVmTEmwqjgjMC80goVIJ6KF+HFMvRArPqDGD+6AK0QbvoOpd/Q
HPNTdnhePImXxinw+nILd/VFcLKCLGOTQLVQREpEE6VlXXf9mVxIx/J7AC7CigOA55OBly1CH1lI
/eo3oP6X3Z3PM8e5ltoS+wwVfrMEBZ7QG4MgLNYVg8fMck+qLbP5ygkw/nEgxTLTnbQf/mAmbmby
0dZImYp2W6j3nep5VCrJOmELqysvDnLj+GMZQVCCcmat62OdFk52Dp4sSF4pz68ryk75cOEHtfnS
ijr8zxRiDZdlI4fiF8gpNn0MmVp0GyKGlCmZ8xoqaJ3vswRhnqRDnp8b1HrISsw2xecWaIiLmIbs
qKWIe8aYIbFr9gWCy8UpCFCBLqW2ZvotAQbHTfmf+wgjkkGmhRFWcUxSI79p180kmC5IQO3kGSzg
17S3XVQ67CI4mtVOKmPhReB5xPF6qUTxW4udexMd6Wn/eK5y//7xPcpYat1aCUpy+KJZ3F5PZ5lw
Lyyr+OlTnRZETwmh/CmYoBYgPoq9J26QCPghm5ZyLGp9/0q+OKAr9aXx0vyXKK63WIhrd4fBSUYR
OzuDL154LJe5Z0ayv3nuFRZfnOj9hyodpVPlUfNIyA+gl3AG4KuzQ/wbs9+IsR20mKstiqol2ivm
8LyT38/YfJkNFM89/AjAUXtj7LiFbGYogoKmffyb6Npvq6rZjgnleLUv4JL31VZutQqThwaSAs1Z
aGp9GquvkIh5p2K6mIQ34YTnUPnvWp/sIXpwwRAcdri7IWRBkOilRZ5wZBI3X3F4EgFFsU1M/XmO
a47hnU4raGi/YBAIrteBC94X853l/HRWl0+U4yc01teZIqTZxSiVqOqmWhHr91QlHLoBhvTSCW05
kOJdWz1QlVZefRS4a0wruA4elfcpcrngOV8K/xwDzO+904QPTETeoZXRKkposFLM3AsQnPZRfBNl
GOnhDkoU4WwFnWOmBzK2o//dMoP5YwTbKocVBogelTL1ip/6B6w72NgD87kGI9UeuHa93ydWT1eW
/uY6aisTf0zCotoz6BVwfY/PMzPAp4082ciC8OMYbXJIZrKqAEnGLukdfrPnjQUz0OKitHH+gz6K
C5di7swcd214tuIF16B952s0CHXD6crP4VYbWq7nXV/7p1gXTOwYLb9TaTRrF8DhESqjzf8rJq9p
2Lon5tj7hIvFiQQ904s4FTJoC3tC1OiDMxskgtdx54vJ7P76IPCOpt81TGlZtdX7ZuWdRalGWzcH
IRYDKRejS929UuyrsC8hlQg+OQXkZnhS00dqhg/Nv6chKx5keBuDPoQIohwQS7bU4c3mUvOHu3TX
rXeSOKayhOyGMOZueRspuBcWJg/NN7mcDPI78q8O4MHJW1wiz72g4/GkCeexL/cUz/zxzEL/6Rz2
YmSLAVhv7D2dxy1zjw65odDDiOAqOh8oNr8F6EQQXmAj5qcWWFIXsB7Y5z05VbefGGhJ1lAoRrVp
nsPF8c7P/57Qlyh0h31cK6qf+P9lbPoiyJ9C560qOwYUQ97YmABc10zXy/BVQHYAJs9gmIBU+YqU
vGzL6RFkIEbGbC1V8NoMdc+81HFXUm2cbC5uA42e2iFzrlWN80ePGKOPYXzo9UCrQ4pPG/v6McWo
YddzXXMPzGkcTyY8Wqc3usXoqF8okP5PjY+cCfCD2JefAH6uc1gPqr6jTy+6C0UeOM8NntWrmvCd
PHSrZgCzI8cBb/gk2VWvyHr8wHgnnL/UifB/0vBG/VPYanNcEkMdSJun7gPnPVhGM59lukRJ8Cuq
jyxg4uIQL9u3oWiBcdAa38hoxNm73AwfKlFqtSSVwzjJJ6mYT5pKuECpnCr1EiYySjBfFfrJJUgG
OaIC+Hg7Yw2hWigfWaYtne3SzGWacGsGKubtOfoUim6GKCuFwwUbLWc7ZY3OljEEzsK2WUbmudw+
0GZE1WNswOdlzJG+Xe3Qkly9T1KFWsu7JLcOAgs4Co8RqGE/g5MEZDC7tsepKpFP2GOjpO/1Ppms
pXHHNDQ2oOgCx3qIYWDmxpUF1AT8j1p7qE6fVm8VL7bSLt69Q7cZQsc3QmV2EPLTME1r7EEqvpdY
nRhziF3lKVJkfgzAbFxQR5a3saNmwd67+laFy7UdX4Z7nupo92BHkSVvUHtu6u6OQYg4oqFs/5Vv
ndSQ+sthUStul75duYsUKXFKn4/WWsdKx/pAUCaKDKSDPcKecFpApfKj4HFN7HnenjGHhx0DmCu6
CknnTfVh+dqAQCMmtQkejPgpqKq7w3d0mxCaxWe5Qzg5yXZplD+puKGVPgKdHxmor2gPD1kpYFfL
xzOw4xSTnCKFWj8zpW3dpexDSBTcZCvPoC0OgDwaqNXgVnG2IsvV2KV1iGaEmjAJr45OIpbQFmb0
QN3pLOs1b6odBnwLiXURAEpFLd+LHKIOVK6k5UEld2EtOfc0qgNXomsQP+TmsrG2ByHXTjUYlYdu
B2Wc+coQwR0BgUtji/NTIRKjAbeZEgBV+W+eL8Fb8+rlxEJE3ZqbVAU4dwDTJ4JP6b9vXm4lptKe
D7sXGkMs+xOPeyJZrA01Nhs1zVEcIiHXbuVvvNFhsWWmCVVch3JUeLTo8Pk+zZQ57qx0v1sd12cg
O6JhVrZIyK26FNrbP7iTNBH5nKkunoFVJcrDEdAPz+A9BhjjMYad/MQcGgeXxg+PTmiowfPSt+u6
1+pcPkkDLOmznjQx6bKUgRHrX9gZHmdhC1Pwc0PqWj1WlqVNnaO9CbJz3H9Pf4i8kbqmQ0ULiKcL
argq2a4CiXroq8dGrCzsDA6psQOkWP7jGVNSdqyomgmKykkX2sVjXzIWZ9Hnce9XHVHJODCuSNjd
6NWw1wEABdXr4RCtAZXQsbErCJb2H4LFyH1kBDu4C8xhRcVEnIr7y0mbCF/yTcORwVaGm6l0pC/P
yWrbB5JjpT13ztekAOWhnT80ykJ9get3k5QsjJm8byKBb8Vul1dS8in+L6PWt3mCMlQ3KlX2+K6n
/6yahM+shSAP7r7bitOfEcPQ+Ataz/35JV1Thq0KqYfURvQp8xGRu0715ufTfkWxj5yqe3TzosX4
oV+IDKw0s04aa+Nzgox4v44Srp4CMUIYCh7hlG5DB3+vIiH+867LWRR6pA0wW7ZsVdHuXczplypW
mX3IWNGVEnpDaSqve9kbrUaMYR81DECtruoGrYoptlUoMou30VZ+lSsAy3slqVqNRZEE3R1wyjfg
ozFn69/0MI5lD9soU57gYKt8KgEuif41+vdNwDY6G7PDoaMQCvpfe2kj26HSN5CN8u9wxpiZvdQl
fus2QaRrka4E6O3MgXX6k5zYCWThtqPjHdci652NO7iAaqJKY8C5jDXdD1tgnQgymMjyRnuyKdMm
MZbZo5QWrY9K7cPLMskV//xlF+9F/UJHVto/NyRVEZD5ZdDvjLymO3d44l+9cexmwTFz6B3dGLm/
93hUkf4flEsn+hQ7QbpJzFwZp9RYp8wvmjMwETCD/2CA+GUyChEuJDgs+rKMIc8LMvuZd8veZKf/
2tHNCvucJqLIWBbVUuCa1QIw31633az1QVR2bsXZk43dOuJZ5I9yypYPWf6/4/oEx9/x0+crrgrv
oLyLAyzXTgSIIfkmzszyRyZVf4aUO6lv5qOb5kYlbe41pkPLbCrgjncwBH0k36KHyZ6ttge3/g1i
rFzxL+6J5m5PsGYNfYRC1W60Q4OoyZIA1h8kEko3KZ235sq3pcYMhDfCOn0S5yDP1Kl+mreITkf+
77hha0C4CK+9LKAETjrbw8iZdW6cHQT0yU1+TZIAIovAQmmTwc1kKmI22xpDE8aXzuuWuBaCAuEF
SqtNNTPhuk9QUPOjCwTwdfiTRxIY79ZlemwYT/K/udRyq7Z4prkObckTexXmxGAV7Vz/rhRFFvjy
uK5wFzt0J9c2gb14dUd24JC5iqFPHA64rxDsHq9CLl9TObaxyuziowWgwDSEJnj57rkJUesnua8m
zjR+6+aM1m1M4wpN8uQTYiEK1zGHiwwkJ2XcNHqm/lx4f06vsbv5nEqxSuTxGj3OJqaxZzShyCft
ldYSujXHOLCexIDMaXQ5jnn7U0qb8YWZjAix/Essz8CJaVqSkk0/qgT/PSZR0k4LTtNXzZTy9tZ3
nkrMAgh03ypFcXYLyOSser2vVYedw7IeLfx0PjDcSu0AH+lOxh4N/tyZS9C/GomlkZ2KecfCDPwW
LnKYtZbxTqz+sMAiJ/LDksHX/+YkA49iCXrLB14GqUaCSUF+kJmNdYyg3J8Cj2GMjm+auamuY3Nj
+0QXl+8AYP+XWgTnioJP+ALw3iE109YkfULwB49pV88hE3Mcy9/mXklKZJnitEjYNNJY3cfaaJcg
pOHODMuKjst3wOt/ou4UZ7CbprXt3pfbAyrlSRlnDRY8s+caSOuGLUkOXdVtUSSl78gtNSjPi/W9
BI/EI2/Wk7QjVxvRHcay1jORSznIbXv1nU1lsrTzJAaL7zJCEAnIAozKkn9LUAMfEzWFQ2LYO2Hd
vOrx28P3ZlHU3VYz8I4kbHbFPHdTcOVw30Vk8XtJmcjc80JxxVDtuXGBCwH/AgpIj52hkKhf3bPx
g+1mqdLdpFDggsSB1Plz7pKEHqwDd53krVcHx83Lgqs3Ev+Rk/80p5IHGPtU5wVedmatjZ0+GwDK
f7wIrJqjKcu0e2oRWw9AcCe6IQB4dN+v5r9QAL5X/sAF3BZwqy4bYAM18lCUvUCr9DQ5Xc3qX8Cy
NwFJSxgtmU5RsUG8adKJGpfAf5TQ30WRStfjvjhA1el9zaErvjJpk4mL10SUJ6dfbbSCMBYnT7a9
zGU28EMBwuWLG4iLEYUI1epJE+Gn5bTBUl0g5jZtiU1lefPBhz5gIFgc/LdeWkgOrrVE3acDqo2q
nrZ8vI+b43vtQhpaGc5L0zTz0wfMeIkmMgw3lHEAsgseFsXjmUMdp/+woFg8OjbuiccITWcTM62D
v1F/TsqJd/9v6gRQ8Ez39nokxPVOnEdyBrOs7KUhULZmFMGbjyOT6nr7NzJQilm3Q1g/0sJ5Da4U
+m+6v9RmUENcwTQv13IOhMj4x6PqMd3Am/La8UvUDr/gCYiLiXoFRkLqHLEnqWcKRq9i5SBBU66r
N9YFnF1mzT/i/xW7W2qiUnK15j5cU3c/39Gec1Q6R4hHwROcKsC/FU+zQnfV95JQFBoWITCNYfSP
MHEuFQiEFVl+f40USYG1fp6DdZxVYbLLQ8eT2YGRlvyMtPoaLqUpjagYnaTF4978GM4d8FSKNBHE
+WL23vYiaXPjxgDKJfA/nomjb8LTu8KdJK2lizBmv0QebhbVsOzySAy84l1wgcBW6xaTwkJ1LyQ0
8blE9zaHBLz6+8sZJWQ1KxfhJA15fJIdqoR5OYp57zk77+OFtqbqJq2YfYusuYp3RPoshotb5zET
eLnlzWykVb8fvdrdta1iocMA6YH2fEJJtr5za3RDvo6tQsdH1PR85O9257MsgEe0uMGcjlzRAnoC
xeosHnrNwLy+asO6unp+XN2ABNoWmGftbuYadkc50nG0TyG2OQ/6AAQocMccEyOyOFF6ODvd25ga
wMB8BXQ2x/3zHiDYFCEVjaM7e7COzRzTlm3J09VVoiRDT8jkcoOWId2Ul+kSsNDhWySj331JpA4v
zNdgRZ9WRvPW8SchmiHFSfub5xr+fnFoeTmtTZ22aCnTj8vOmb/xnTkj3AdY4AE8tt09+hlYQhXi
1NZTxAobnNJj/72kJL8lL5rJ4ZBvsPqszuo7AoqhF+LHNu2txtkSukhfQBgM+GUaoSJuXRFT+NYF
9qPf/MLtgbwEN71kZvf8DgqSvjNAJ2Y84/m/7IBhMBn0FkkauD+FgDoYJBRqqJeMDOG9ArRgsrpC
xCsuyNVt0PUe/BowjLDKqCmimc6TKRP2ND8LHBEpKKv9WIqBmfIMRaf3Mt/XXgsZoP2JqGUk8m01
OFf3UM3UI9sCMS89FSlwwDX65a7lrLPq1m3wCHjS4mMSQbNvOaAwNJZzTD41K9Wn6PZL0Qy+6qXZ
5VfBWZS/U7/hCuRb6lhkgbzCRNQAXLGxVIOWsiak5OcILJw0/gxAH8sHimfpBHRbKr6mn/VygwWE
2fHHadjKtBgpxZLVZ/GOGGokSfSSL4TO3XryOL9KRUk+nMulxHkhqDLWU1f0OaHH8gNwW4qWuz09
Euyh6BxL0d84MUg9SgweiF+kC738CUl+SWnmHRC/zBVqo5T7MAeiuXUsrUIng+NAdGnR2nLbDe0Z
+7uL+/m3B1QgYiTdDAwZ1VfK+0l9ErMgMo/SJKtm0j3mrX8ytvQyKVgBH2jiloQqr78LOfc8MgMl
Std5c+XAe2osY45gUy388lBxd1n3zRjKXewSCiOHgUxAwgl6oX3TJXflewH55OqLaidgWmv5ck2N
pvNT9Hif7FapCJvhFdwZgfW2D2d6OvDp/VO6rIa5QwspjdZybfvNiCope3CNPFnYkBS+fXm47hXL
wMnwy95xUllVLXjQAbaLGrmYawXFyX2FToA/cKM12FhyC5CvPVxyhiEc9BswhY4B0pcJqfJkI+i6
DplEeRnj8q+08TpQ1zEr9jJtLQLEaBs17Vot4RIJgPGJCcoTqJQuE2Eh1xBjzGQZr63mdVV38BgL
ScAjMMVimNn89OXsRtZDjvbGcniMTb4Yf7WuQyhmPUThzTzTukhsy0GYO4AVWgbr2ailUCEXpOh6
Ay9fC/Fsh4lk7EJ6PrsrcUslHvxT17+sIXzHa4fnyGVewjaRjHbb8tar2Sqs2yUNtH/tVfYstqij
mXLRE9wm1P9db23pq8/xukbR0bFXBQ9ENgYxkB674t1At/5WI5BzupDmruj93NH3uJRp0lA0cLdX
yxdEPfs/UAjDupi8nl0xBwWxhnjgDv+u52wZShsfR4xQYWL8g/wZIjQuv+0UyUJuW10xixasb4WP
WYajA8UepCDcJ3tN13ZgoM9TesZ2cV7gTq0iblCb3kwleoldcZRQ1JF5oLc8WbleXaNL55ivH8op
28e7Ay0LTTGs4aUnID9UnZrOtK6DdDekdXNZLA2mAGItVFTZ8jLCBLL8zpo8dUMQRLdxsTixp/bU
zlaHwCqsrWGcMO+PhFLFu1j+wkxoPp0BIyJqriSEQZuynyqs/FjZlqrg8BhR0mTFNKlq12mHP3Tb
h6CurbCPkNUQhxVybNhWARuP9h8dVg2JpA36XkEd8pzAUirpWGxmP52+Kf2QKFgwlhpwNdXYRxoI
AIdPm7eZBnubyeW09ZvurHK/Lh61uSTIYvylgzMRyZMzjtvd2NuOdGFs4J6DQ+jx4YwbEprkUR6w
WNDZ2A2fv7RlfBUaTRs8yXZ5BIrQsXxWDnjUMBIUaJzufu/CR9T3qEgkLFtlom5Dnwt5/yq+4T+h
5wcOxkrLTFXeRsKg2JMAJMqwT0CO1n3iKu3HgkqEKpt/WqrxXuCadmiPSiiwh2Sw2ATE/RLsFVgM
rsYBcmr37Ppmq2J4YXhuWY2YJKAtJgkiUAwxTWaOMfZ6Sjx5zriYUhMMuHSNt2UoVCCNP2V6GkIn
ZZq4oI5WcSEBiWHCxAXPFWzLiOxBH3dXzCqErhqa1Yu0E3H2gzjC+rgzT6WFYMlYGOtPw3EPfEYS
pjgL2e1wJjUnYhp9Ay2UICqssmMcpJdAD/RRNsO6/RbuBvXC79UX8poZj7WIuEMV2pbI46Mzf7EN
XaF8/hDl0oI5geD4s0ne4138pEdKY2i5I0Qjyj0M+ksHxbd/meVsVlUlRDAMir/hLX5Fzl9CNCyz
p2k6484xpjowbmiEbov7fdF1f/5/NRExJwIdLF9q0Jl+vEL6/W+oC1BgnsfIzwLcZOnqNdg7lM9z
leN/4SgK4PLldPKTvWlfNkJXgvGQ/dNRjb0rwzeZeJIbrp4cmkEChx8TuHmwG9LoWwfP80oCCvcz
ojNIKBF9LT5dwYXyep5NQbzUs1rd5QyikE/acUnL219+GyAYRCaJhYoc3HEEZ6+cFNpIIx83abJE
TxyWCpiJco44Zxj/UJzxTzqhMD7fHvYe8BLtK5t1DElFl/JtJJGqN+ODNIPHb1rFlVmNYaSTMVWM
7xNx9NkJ9/rRURmCmpBixo0YZ7sRxHkdvRXuoLGmqLrDmrsQurgD+ewn84YSI0DW1rMxE51kDhvg
QbqGTVx+TscdoFEQ4AA1DLeTR8OFfKaemyp99dLEz0RE5bgAJ8jPuLf2l0ecFFE4Ta9H+AN7WWip
uQXZIWNxBXVDgP1oDiuHXhZC5GL66Ny/CHez4dCbPvyxkt5bPE+QNPzmwljcFsef9h2lJstFopvf
Oz94BwZ1LuLJDyES0ENsLXZRX4wOvLqoOquF+lyXx8PZoJNJ0J6c6xgckIROjQHCcjs47BDGB3L/
i97M5rLM7f5bqfmMrtn+VNOlBRO1VUk/WdqbSEk9+D4hdcAGggssLGOb6gBJme9v0pPcXQMLgV0a
cCK9L7zVlBFvD8dFBA801hjzKVZCNN5DhqDtQhTJz6gfjKXEPrGaGY/OhWuhd23MJklQjjlyyIU/
cEJTJv7QIl/StJ45IYl2A5OD7y2+2qBwNZUIzTc02maWJXxluY1+uSXwFzMNDSHLUvZEVhw2/Hha
3c+PnPaxr4pjT5JzqwMn6abOs5HNWISDPNQGNdjrvH9dqSaftZNh6Y9De0ZgdY+62WD8rmtvu1f7
KF/VHlP0+51yvdOFxp0+rICDuL4aTIjIGwTagyFRg/W1jBZnQem8IweIW4woIY+PcvmSkN6oLcY4
z057C4SFUpAglWZMugtTi+1nJCviQXK3LgjK5exyCutZsDMsG5WYHXaOecpJjfS4AMUX99NsdKBH
4t1TzD1Nt88MfpBT50ln6MKnFvIhr2MOfsIye6naKJxvgysytPUeD9Uur+Y37n69W6gxTroxFjKz
nfGyirpFcqFUhgUD5yAk1AqWmDM3og3Ebt7BxadeNYoggVtH3EafkfmFRcNnRXCq1KP2kF+o0JJY
1hyoLStIOR6LsJr0VAL53TWZUq+pcZ1dp3Us+CVrCT3vaPTvKtPomS42g/KqZY5L5eKNkcDC5MqA
TGUBJxqgLbl7QKMf+b92tJHOSpiN3YCCOk95nonvZF7SKGWdJnDXyo0HTz31F/fovmBp0LHO0Sa6
DskQh2U29qLKs3W9leV55pg/vIheVtp+b0C59qrRo7Gi06ljvLeYKp1ix0w3/Rq32KKHbbZ6Ffr7
nQEeN7Km59WuChCkybxv5PFyc8haKJmgnVGk1qNE0Jjr+cWdhDjnsY5cf9FdAHhmdD7xL8oUFZ5J
AkQIqMMU9oLGTTSiDgFO4U/xMRbFyAqU7v4xcoD9titzbnQV04tAGNxea1ESS0X/U9B41Ldh1nj4
AaV2CPSFobZpB66BaHhD3+y6W1oJppbr7xmHgTzzSdkI8uISVJZU55GM1dyDxreRfz3Iax6Dy6u3
MdICOIAtGXF6GRdZVEfLk2fs9muggZJznAt2Ypfn8qVEu4t44+AdjXnsOWNzxI+0Iq9GBLsVbwCc
wzEkTBg6pT8IDIiknJOILUE6bGVwlBAT14mQpKWsASCgO5lXvBh6p2B76n9jwnwty7mcL6Ts1Y44
mcxJZifM44pBM2P6Ish6qdwMfh6CPBQVNZK/cYYPkubKd9oxDHKgxdJ7/sKMPsKeAI/Eoie4NQFA
W/BXZjGH3bjzwbY5u1K6jqTSxpP2ANWFcPhyP/vK6tPgrOtNhHqjKLjhggj5S1GfPuVzToHrOYq2
UqhQX1rYoyHINAsUCsZhFSpkUNqu5DqLQQKWhDxuXiIhUKA7fhuUloQge2PfSaGB8Gqp2ycQf5B0
YUsgyo5v9XpFdQmTXXmeNUdM4f5LZly8tHgX7pV3qq4Z7nA4v5AqRhATcShpT4z/y0N4lDKvmsMW
Wug/BvTpjkUwhXNvMsXQMs3NdPqxx74PjtTuI95hRI/e7Dx6wwm3WuvEfFLTYx7NpisOYGd4W7IY
uWBLmab1AQiR4TVuuiGoG9fpora1kj0Hq+cYt4QtFX3ZIgnkLDzyBNV/9mMxCPTuF17Ybda+wzMc
60B9tpE7HpqsK7cZCdTHsBmCDjkGz+Dq+3Jx3noW6iXo+UkcnAE15US0nOFMf3CA+ruwy3Jcs/sI
oeJtprCm1q8Z4KAFEMETfqf5fPJha4ah+cF7PvjTdwHrUOe86rRSQRc09+Sd5Wd5cPAleWu8kYyF
gcyMa8McC4ZdVZKO9JSuZunsUF8SSimX/wdCpVT1WFuzv5K1RATArGC2NZiHwzeL/uuAV4ukcSiT
yhaCHE12n5gfF8z4WVYaTUKPuOZC6/Yvyv7kC6zVgiK+HMrs6Bl5lNmYxYN0IOJKJcGnp8QIo4Be
BkFnbfA/UNR4w97GgnyHqWXQfJamOEcwXftMyX5iV/3/CoM/8fut3whBstMfodhD7H8X2AiqNbxF
JmKdsWY+uFvssO5qUMlkKHqiACCFu8xcUMw9GlRwE+BTtEmuUXAH3iMiJkHjdAtwXRMbPfs1s7VU
uXAOB47C0fENkc01nfi5SmczlKeupZQ+vN95sapeM834WpJhr4MFUOQRgNcvtYQl/V0aWyHl7A/w
0KNfRaxm+ou2Hm3DfHV1aXcnZtcHpbDfIgapk7CRS1s3SPtJPwt2gv+ev+WP5/xMQm1ACPJXs2iK
kqJEMF2l8BiH3rwUivKy2CvV9xmQpE2CGuFenFm0mtCbBRMUorYzrVohmixLJpd8Db3nrbiff/f+
1msKEtTgGnXhcpR7Gy+ORVoBg5di943+QPFZkpz+JsbE0AKPvYvZ/1BzsN5RMAT/mCrfKT3RjZ4N
ObFn7poeYwEM4/kBmFmii/XTA/qm+kFs97v8ydGNYe1+xqiTDQ0Kkja61Y3100+m2uWs8QGPbatY
Vtd87va6O3uuEK4ONB2llcpD1AdOYoYpVv7pen8eVP7YW/9wAOtYSbZ7LFq3yA9cAgZ2NiBc83k+
mvbsspwLCl7cld1B5739VPSwoNJN2OsPsUnSg8rNojRREFWuNoiIz3kbyELqMWb/jxVU7Wv7lUYw
X98b5dUKWU+Qk7oVi9hzbrynpPCZ6aCa8i58ETWi48D3Vj4apDczn82/f89tNmoadvPbLdzfSFpF
5k/iW6VIsQeqf2eYBVMFjLHXiRbtSJN6vc1EQ3+TpYdFwxtey20K58EVUp+VzO7P8gtBD1BFXKI2
+fJ6DX+JJmAlcZPym1p2jjUgwD2mI2jGfUtyMVzm/nn5XgtiZ17sljbbK80+LXFD4qprMvTNQBxN
cxnjYQdGtubKpeFzuJp8ZzMEYMY4YDqvQADPftwgW6SVu1YiVge52+bbJiulkSabIJug25fglPZ/
WPRxvH/6DZkkQdEWmKMtrqeSpa104eilEIrdmBraPN8Ai8pXUH6TxZWaW2FRTHeIAjtYCuoeYB5M
WraxlbiTkgGQQPsETQZhpqwJR+lzhxU4apJbQ7tg4KxiMT8DN4vfUTJatiTGupZt3lN3F/Y4RWIO
7FYeCT26vEcZosKCXKKD1s/iczcfL8fy4RIwpxQZmJFDM2x44PTpRofsS6ZywYlzrkDX1fwO9P6r
2IMLosaEfTAGtA+GChZasBCNycF/UUzkC4y1k8Ke7+SjTEaC4jXdHzF+zD+iystUgBGhdumSArek
Wh7B6RX0fBvD6qxkGReyAHd0W1bGjgXETrQgkGQLg/viAARV6g8HJnhQCtzPTLyxEs7Fn2GDw723
q65b2sidA3kLKCjNeeMxk4yzIjzs28xlYBRCA/AGES1KUrGo3QcuCFyCWPjZx0OC73OyklgDy2Wh
1QT3GPYJJ0N6IDDnTbapaZCy5AsAEuldWww7tDOKewd7enOpEkwYOTQcinAXwszto6a0hvfR9Og6
QmHAYDgjNIuqKVWhWNtSb0M7Yzjm6oixC0LyKoftSYtRcQfZzRVjTD8QD4njBKffbuY7xVPRwvda
K4BXce6eJIjVLbmCe7iTEigyJOa+atY69TfNUQvGji/68XHQmDIXvWD72ynLd9g57HDuuxWdF8D7
Z3LyOy2mcUfmQunELSB4C+FRTpOcmdVqUXhe7ckR3YqMc1HRWfoFVWzCV3b5XcamdfSyq4HjeJwl
3+LIj2bk+gfcCFuSw/84+hYtk1fNNDMD7bnVVkdPO+9sPQtd3ZLsTibSJiXVGBq6jVwQoKDWTaYs
8Tx6Ovqv4godBdc4HaP0uK5m3OVNnuK9Q2svVZzEz7X/F1Ore1MbGHOlVb6BGOnRf5wdw3TAU0sl
DCuapopm4uTvJ5+gSbp0JPJy8Fc8gWiQ5v7KM2R4HzbV4eRYhR10yeECbTKzEoYJrAxCnQNL4tvk
dPLEzv9YNy/fmMGb2pF2Gc/+xf/f59f/AbQnh2OU+WQ8OINFSqeba6lc1GQgMVRMwHtv7HMbJHQD
iL1uQUEIw0qxkEdwmnmdnp6+CZaocjnKxqjAgEcupxry4oKXhjzfxwNOraNFJ1F0fzHZYCfxLEdU
diPucAz3NAI+VAcQCpIp7MTl87rLje+0BMgNlijCh0kWonfBbBeZYjEetqbabvgJRQzY5jMPq4nl
XKShF7rsYohI5QzKni6Wd8QFCB+wM+Xd07M1QgGHW635H9R0Xt56H/aZMDV1qSHX/TMlBddQaCYD
ADMKnXlG+YdQIjMZK5CBmGXhtLjxIHYTVbHlNBBiZ73fjyPfiszcaqKReEP+M3Ole7ykOftSuCET
DMW1tYMqdU4QU8Tq+0y0YduZFy9QHuoxQ9WE7/cw9xd+vDMRdRioI5flOhzFkmOLCK1yp0SkTBRk
4hNKEJCZ0W0dKl7V/jDOceWKeT0W/wY0J7uMORdbYbymvNH7CWAg+maDDwFr48ccp6KGm6ZqDO4T
cGrM6FURZb1Cyy1ir4K2fYR96+n2s4xQFGg+IiQ6xMMKPI9X6/21K2+bO401+twfi1j3K3sy2Jec
Z1lcK6iGsl9AqYf5OEX3xxEYSNKM0Q4QOJPmkzfho41ePbhcr/9D/WNws5HjiFJh4BhTEg1f2Hh+
rJsyWsQOkeSOTLz+tffkOKAa/ZhWrJ44vTmKUe507uGh/0V33UHDARU9FI0zh3iJ3JDjyAhtfeaV
4rD2b/Y7Gkxot6BrB2pjKcE8fMF2Y8OQ7W80Zh7y9vgXb+taMXQMAjGCj2HB/QyJmEjEHB+1ezpC
4Yn82hpzESsVGNTvCh6FTWMpOs2qJZBJbrN1rcKw71rs4X51ELDu/b4WoODbcO2aYO31l4bkIxv3
XALgz6ICN2Da/82yXDKT8WQJ3G0unc+wZ7UuUB1vqU9veRlJ7TQcQzQ7805nQnHRiPkMgegIdDjs
k11ZTsVn41j+Kasdg6EkoeUblFKeFY2EcNQ2OzxgFNMf8oaA79A5/Os7kVgQhpR48St3GROrpULf
L5pxudBeSG8ALZokyF25wYarTSBow3O6h/RDn/irhORpnU6+ylXlFNGYZuC2NK+yFOnGhDpg9ObW
t+nNrVP6DptVgsHg2a6V2srl1/re8NL+o6pfNGLLKc2s5heu5N0p5wwc1SppZV2wYNMh8u8JOwDE
pDzCih3DQlQm7ofUg8ic30yDGqIYys/n5z9r956EGEwp6AdcXy4MmPHwEBtVqROVFnN//wYQv/5k
6CgYxn+Tklqoq6pUh56Rap6b3an0CMYt0y4G0L2jhPgjZLFnSp9uhZ9vR3jvO0iI+6xUDRWg3tqo
4XAPJx50LQ/RLswQXMjQznI0YHNrQXwIZUtuOlEAMJ7n3LeGxodI4lk8NRPt2kdxO7imAE240qie
zn6+JFdgdVtTI3MfnXnRwH0U2FDe7qSiA9KQPjkEKsOtHDhLZKcCNI7nX+S1orgl5Ku9wVa/G2EH
a2AenjhzVr1mvQwS0tPymGNL2yuqb5MbrfBA3CvSLH6iemO3OhDbGEmTpQ01Xn5arKBLJfdfXwft
GHTjVyrDr4utrrTp6+gUjpJmOE+WfEvGoQkFuNDUAIm2kXtVpAcQYO+/awJmXXO0UkqKi9JTbFU0
nLszzurIrIsc8qyUh3S2T2oShRP+lIUMTsYaQUTYx4Tuvpy8A3H9q3QtPYtyYilZ3nizOX0DXZpv
rBy8RLtcDyRMtbTnYMrxdaJj9Iw50+nltPSHmuNITcBbkMUtV3AzwFISpruApJonIJdzSBXhfYGQ
Ovnnz/tXZv3hpoS02mRPu850nAOLqLzqpVg3a5E6MYA3LlHi9WkNJqZnWWfucYYJEsgkK3jijBh6
8NRUGlIleCOTQVtBNLtho9ISKuU11msr0Q73fDndKrbCNFkGJLNl7wa3sDBi6r6uSgICpGb51U6L
mN5+LrbXqF0PoGfCqbxXdFnn8Ftofzz1gxGARjE5OXBni6jiyzxg2xsva7NMSLafWscg8ALq0T8K
h4m3IQlbDMfTBLx3KJI3AuoVJPxIvBFmGaneNQiSwR5q911ZWN8zEy6pFVRq7xGGwqNXuu78a9e8
K3IGG0Y3A7oBaR2LLPOml/dOB/XsyCjwcWtyc5DZ6l85ZS1wo9ZLbVRlMK891WPt4iqDK7tj54S1
q2OBhzqKULSNZ7PwSa3JXVkMVK3OVKAwsSznhItJ1aUwAoyWD7q/87S4LkHwJ+Ots1KXUeeCFuvF
rP2imt6vGjloSmfvS9/wx7tCtq8M0IX6jKmMumb8Z9LSVNYII/1W1PqCnMBzhySDcTQ/Lri0yCZS
cPCJp3j7jGTFvdIX0jLVFOrg8986cnpRK3XwhaS8ODjE4oSrJjEODvMFuTqsKdIagAYHTIncdsEr
KzA5U3/sdMluKDg3UMeoi31WEDI9PDq/qRX/65SS644v/WmESAu7GwiUrHMIAy1gXowFn/YvG+af
AJhh5c5mZUqTk8F2OucPL40Cwnj+GLMkvE+Hy9jI1/HJEp4g611FG4zbVg4+3kKq+jNGWVruHz1b
wLwzHfNAhS3iTnO+z5Dpsn9NPjvN8/4/3xS3Rn3iS3Sa/51X8O2V9ySbkC3esFgD3j4AHisx56VN
eRk+jk+PYBTs32hq89VyvuQ4S1AtLyOk4fMfqK1z2XDDnwxeyRNLjdyQ7YrTpO46zReqjiUQUYC4
kuWsnbmrICKggpN+9P+zHBPSfrDMTsQnzM7E7vOu2LnFWTuPfAFSUTeULZzg1M4mHVggEKr3Pddz
Ede+2KDirfViccV2RMWqIFP03lxsRoYUFo8vLss3guKoFUctPp7rZEk50lyGYuGlUL3R2IazC/cd
s08mtDh4lCoCd7KsSy25cYoZC46suPsco9jPWw9+NF7UROILSn0F0D7hu6uS4xWlEh3H6TostMOP
HNN9dznZz2VZbt4Q14fcRiZA9kszmC2qMnX5nLDQdzh1jTEsSwtTIGnGd8qLCSxSMHeCzFVeXZpx
3jdYItvTf4w+stkRjySBjwBfCLiAyN395C7h4i7deelvLREBlA9iDyyeKoPIR+UziYDh8uPhcW9G
62PJkhZbIvDH0ehTbuFhNqxC+tPEYC8M3SID7uhsbS/u6xqxM3nOK3CodTz8kLej3fS0eZNA0dlt
exU/MVwUVAadUA8rHjAElHvCuKkkqWrT4ZmDcVyLQHnVzVio3/htMpa1tT3vCiAoHvlhweDmKPqX
u7OMeKGfK2dnq+V6USm0q8QNkflTgRiGbLBvp+HFtRmzG7MQlekm3ljHpahO81hoNVEd89CTpf24
O5huSl4YWRKlAy5rB3nWkKFnC3SKFbj+Xew3IRtSD0jZZi22p7msQY9KnwuVzd9nt/qehVP2Zpad
PxLnDJomzjesqbOkLo4d0qSkrjCqZ/oaiDWkrur016b1BB+9Vr7V9VHWYaadY+c6UsRee51Ctkxj
KWVEdYnlAKcsGTGxWqjUxQwXKjffbcVwbyHCSPWRgoH3D8mnbn2reVtfEpGHxlap1p7jDRkBfFTq
s1vscgAbTS+Fmyu0VIJeqUlGg7EOH7IViEGHoQ1f+AuEc5J09Wj5JAPUG+vy8XBVgrAp3Oe/sWdu
Gn8noSrPN2zxgy84AHsqKseaDhgUoLTDHoxsjO4hkOPShNRrYV690WfWxuKosL/Teo4TmMgQoZi3
JBr0wYOJ1MNmiSNLZsAJ2MjvnZPoalurL02FwD7BMyeMFvOqirnoInEo69xhwYL2xOjzoeovlgiU
xJCMqfks8G/4qfPJWTBXbSKqOaDuVRmFXHukwL/tXrhNt48miFf/s9KlHJJRq42pSOTxLAzr7LJe
NI3OXKhkgNOSwqgHIraS1tI6bHSsWAmdZbCnsDFhjb//dUdlSAdU92BeIAL/PGCTOIF/CdzQ+pYv
r0Q1SXB11mc2yuNcbtLreeNFB+eeIxBWtven/nkFTVLAnIPp4pJNeEwOQXvuN761rCiSMFfqtiAS
nBpQr/u3hjSXnERRq21TsLWFi0EISg6imX0gSLkNa9cNalwMtoL21NmB8RsYHdCgTWFTuHQv5e+o
3ehz+qAaYeUfwm05qLThenLF+zaXRwUuUp0ulXoDG1i60jx/aprHwccOS9/9P36Bv2N6XTcf4y/T
S/QRIz8uwo5cYclWH7PKMPNJ5LuGCx35XCgKgwNFlKjVn3ALccf+zmzRJdxSDP3/edsODXtDXUAz
Ur/RTjDS923QQLY4MwPGIXu3wTEUZkmyfteAtpkgvtY8RhhJIX8ixoB4O516j6ubqYvOEvRMPt8T
QrarYUSgvQ8aElnBBBU+/xzyDKCCxXkFMF3jTmi/w6l2zMVbVymi/s2zNBSj4eMBhWCZ1y+/yamN
FpPzBXwJCIGEMv1qNGgbV2pC7ma6V9M6VVVHj80S04zgXhPJKYYKGGQqbIRUkoBEaRrLeCvrofOc
F4FMz2zR1tX13qxePISwLNxmTQRNLHLOpR/+K2xbJt6NYB+SzGxusRUZ2zTPKpgiYgIashVOMQvD
bqhhUGOBESLlmXoFugA9brHRs3LpMlOzRs7M/pcM8FBiNwJltlwlahxqt+iBRQwLCbcgrBSz+MPN
tP8iNQijJaorX4HC4nwGNKAfjxPr0uipsc8VZxC/l4u4hVLgw50K3M4XiO/bQ7ky2gtVcwwJdrz9
xUpORbbJZ4WHTAh2odUnQSF8CCYdYucmZgPE5WDhhY2YVXLXL3m7Y9naCFhgSg1byY0Fegfdblad
RSirtlKS9YLo1jdXKJW9BnLpgcd4bkiOQ90lT7vK0t2O8QIsdo+2/oYSPMQSegNWxeugAgpb7BlN
69SjA7JYMxd0JSa/GGvqOTmTuH00E+WTh2vO5A2JDwnvrBWJyA7Bb75SjPq3JoCfIQKCqFAYOZNf
cwBo+67NfTnSZB0JJXL6/CbtpgISdw5AYlGEE8hDEzz2q+7UIMIS+4HJ9dngMLBTTDqmNU5RldMR
abyyZGHcyLnyIVmt+gUKuriKLx1YdqkeYA0dyu49Ais1nDtwuzkAT7AR+xb07QazEuY6vk1orvaO
S78dWiEbtuK2L+eq6i8Dcxw5aKv79ZiX8e1AFZ51dAJtf4ahaAuZN6G0mxBLVIV2Ck30LL8JPklJ
RjMEt5FScyXAR0Yf4c6SVtC+qUNoGI0bBomgVdN97A6E049Ul00mn+cbV719Y90kY9tEJ8iR0LBC
F+xlCbWojW2rrXKWpbgImOeEJTHmbYBiJZiCev7TF02LFjcGROHTBdRxskI2oAwPWcbgpVyj3mBb
dS9hE7xHv4TfSkInjr8OR8VoZSLq9j2tgzS+I+jLCO48vYBQRyIYnlO4B8nCbxnnseljOlB+W5PY
nx4Wfezha35JEEh5/tgVMsnZQHKdvzDLb02PNv/4IPlCA4nKuScRww6WXbzYqJW7jphAL814+61R
c9O9wCUDgfFLCKamTpbpWp8ikkqRoBi+Y4nm0YKqg2T+5A2IA6DigLKUDfEM0nrHyBdyvgEOHABs
u42ZPdtsmDbBFqk/VpfXHT+x0HaVfv6LeASadIul9QylZrG3d8ftDzwqbK4q7ZBmGiT84FVvEtYl
uE4kK5+B8RXj7zF2tCCS5Ix0zAFiCFkbFf9KtrOHsIXIKToZblrO++nN+wssbuSgiia2qgukKlbk
yJnqxCisAhb/v1mIx5srVtEHqM78NNqASMCgU4RoBdAnPFRJfLHy1pgw0Xel/caRfkd8UQ8keRG4
63TZptMIqJJ/aNERELYk1QlmwAKl4Ate5LBMkHHctCsZj7vAffkmsLPdPPUBSPQsdRqRqs2CMxmI
Ai5RXCtpz61Slbe8pBVgSOIneUNv2Ipuf8PLZShJNzM78fzJlvI6ToujYrcoBXK4ghZiolC3cGeO
eWqsYBEBroZD7mwqLWwtlhCte1toloArpe6fYTDVHMMpZE7DH5d9Zp3J7rb38ISlwOaGVsyDlR9O
U0XvMd3xgYbVXewImfcE1YSErXgDZMue4cRElhdrKqjz4XGIFAIPJS5pWpDFeo2y3+r3QySbfgO2
RIFu1vKoKUtfn/rIs8BDMcA02deOuS9da6C18HQoIY09JbBPpSS2oacoOMJ3laed9vM9HUbhKQh3
zQ/6I71OUkbmG0zL+pOM/UQo+h7XmUKz9AG1YcW/y1UK9loc/n+IHay1BxDajkqSZNx93xT1Wavk
LcL0qEDS19F2gk5PWh0zmiqumPsJn8T+NdZ7M7g2utKaCHarliD9fLY9fuQg+AFqX6WNlBXP4MaH
BEbaFLQ19AR8xtMUWeIzhFg3tjoQ/xG6658dmN4ljeaoW2JWoE5oWtcnpMwUXwuR0toUeMjLtAbq
EAZbDADshQLWHoIvz9FJmnhjWvOKDJp8YvBC8ILqdQXaFPRdzGfqOYYHWdiYHY4YbtIbYmaCEkOO
rNVrfLCFZ1tHdJdl+RF+RWqyadXZHgn80jiZwTcuOSkRi4ev1iUhTbwnJxpaGD5SbfPvAJAqIl6n
YsM8OKaZrkbeqzrXUPLmUqxWuNIyFMX1sNElclkizf6sP1DBm6tRWKXlv49MROqtmKuB+81+puNJ
6OR7BBorRmTx7n0eqFplAm0+cZeEyvo83BEGpxzxnoxrM9gAmF3RWYOAv7H3LZTCJm9y0F8aWgS7
rnXbUna4RemqMvuhtEovAQu/QsqMXCOmQ27Kdd2Ik4GdWgasAfdPJcr5SpfntoG4MNfeYWMDjwAx
HRq9KXxjuq1RqJIxP0RdswqhX8mH/52cTYe2YKTirq1NJwq8nS+UozBoj6um/1oUTcUgxMYKx8gm
U0RaaSgJCfmXyYjcA+x2B5jCXdS5oOwgKmE723/Qdey6BRYfLtDhPHF/iR7QmHs6T32AmNedSM7p
+MI7qPj119IELu2SCNMiEe49iuoWjvD+jx5BatvZr1RxUAT7GiKjBLjt51T5nDaPSHyYyEgAXDzM
vfw7WmGPRHq2eZ9GdpCViMhwXFoOWK+6tuo1d1jxUwCh3zCnnp1rzL14w0lM7uh9Le/kF+D0Xmdm
ZFJ8YplUgOV0WVMYmt4Ab7hReNs/ias624mYl0+yEdxnpWwdOge+2ozP9oSOvmVqYnQqo4qn7yUq
LpBesS0FjnTtIn0B/sC85FfBGN1UiHD4cx4Xftfqefn5mUqxadZbgbpcHkIkNS0UVtTWR20/1TUb
3erE39zlzEZIMiHVi2h3gJU5TEX3flXTtjTMyx9EXODwrCyxG6ZFH9YjWHyAbYJMtfB7U8up+UIZ
RtKtavp15daEFT9cbdepw35paI002wXVirmBldLuHT8mm8jhIlj4c2PtkaxJEttDT5DOAH3HmPxW
5Tewjg0vfOYFgnmbeyN3oVArw0nffIP6sbf4OEUy8IIXjQcV+8umLnoc2lumkME/pf0I+LzpOHus
UrDe5dwumQFrSb/jCZE6iAfdquFxRphYpOayu8CeILvgU5D8fZJLrkflDSl+xHW5gpnGXnUl7CmV
d6sSgmiTd1ACKZgDLDn8YJfFS/74JvS6+ndGk4sAlYK5jYUVYPrKz8KkVZY31dGl5hKEXDPGqKIs
DUcbKOnx4f64OOWQijayxO04yzz6mG1E6uqE3mhNc3yizSCqJ97N+AphsRIfgC1ksOaKslKNgpsR
60tEWXPeV8wR3b9ZgHhijvmGVfLk93v78kaAWasalHo262Jka5KqVkXTzws/tv0dCtUVb5R77xSx
+oanLYLDliuDVwD39fUZP4WsnL015X1tvTAA5vyashD/Fqf6lCRC4teBZd1tJAOl1JsfA9O0+o6R
jdVZREVXIbwoJCdZBmj4HfZuu00ycsNSwR6jQ/pKSvUcylXBrOgJgYMGJokr8vejJdqDXxf34La2
cLzDr9SGXnWlw9ofy2rSygYoc7ocIKVEjknUbYnEMecKXMhyGunDfoa0+h0RoAK3zdzyvrRjOT45
qKu+Rb3gGSYMCrZpbAvjscjbeWHG4mL2XgnjU3cU07pxzvulZkGucQqnHslXXHUjYJGlxmN5iiJ/
ietjqoQUo3YXhzsg2YKPS3VgvC7Cl/RTa3wNk07/q3gu2Rspc40LLxhH7GcS8HIL9mpFh3teU8N4
KqIpzGw4ILfaw+1csOTtK9Lr8+dCXyAl5krD4183AGguRi19L9uRCjuB2smudIui5ckQxuHu5qz0
UprmiPWCskFCQQngUpfLIpEKdq0+qV+1BX2HxcHbJ5sNIW0oqaq05cipfRazArOZipoP/QgzUQlv
m/u0fBvCc2XyKhyN/9VOWynGW+usIA+En/cYa3RqquAVddK+GsbtGAQkfGwJNYF18GbWFzjIVMLv
Wk6uX6NhRZJRvQHpyCyLf2X2usR5cyKkK6I0ah44q3wdwX9a6tWtFSrcdTgAX1lsF57YLS4gilrg
q62iJBUu38/cR6yEoPDS9muXelq+ioIK5tI5CROInfr2BnrKbcL7sjEJBrNzIuzfsBaWN6ffFSP1
Q9Zj2f0x/QDiFebPT3JwN4uSjiJjYy0pQ5CMktpVwdircwXOKnC1ezJz2E9L0uHHte6F3etEzu50
viHkpFaFTSZNKTf0JNAsy6mYS9JOfOjL51HcHfZcwc0xUS88XERABA0NueR8E5OO35fxHprGiO3Y
H/NHDv+0Pd+RY7+9cMM5y3NA8PFn+AUv2Drz4V4rk6WBT69a1KdYJk0brbAqQHZj7HMrB3odnmcA
JpgY9EdJUilBffu50j6uYajl5lxhi8ylFAiEliRNWQjkc4lGxXQ7byqgo7exPHPf5CmzKZO+MzNw
c1rR9Ox5fx73xz8Mc7neVP66DZYfaEk+MquMjmg0yGYUAynXXV2IwcQF9PBLxcgT2bSgoO3Iodzc
BjNBXkySp68BFtJNnW3pF73f4vZMBdujSI1BY8I2m89GN+ZL00D7WKS29TINFzIZdtBP9Fa7L4oS
dQaTmCjcAenQ0BqOGWzgDSXCZN4XqKBmRyTw8iqqh9IOisL7ZnvlL3yIIoL50JKxVRzjZMtNXf0B
PwntfcJRMpD36xQJr2FP1KQXwLhkciY65fI10M0iIpKLJl9kCjkm98EDR7p1Ii2vT6lQazHV8HOe
0f+N1oXnE4g94PBeWMypED2WD14Cs14s4B42WncjBah3F/Q/dJY+QIEW0FT/DSDJS4a1wL8uhBii
eTVZFFLIKFvwU5zhW2RACH+hU54/DrEoQehpCeKOswzHedGuanBhrWonZyHIsSZD1YT4An6LZ4wn
Uawe/Fa9ILPK/h6pl7v1d31RpiOHSBhij3vmbdsC7IQtZud/+5XFfSmfP1jnMdRQbvbjhSlhyYps
BIVAj+7V5BW/lYi5CMw1y8T5VcN6FJaQ7Zhcf4TbakNLWUs6oxSe0tA8Bni7x4LJb/JuHpg49OE/
9GaGShXx6KnpMOkXrKtHaFxrm/sYAmWOqnIczuiZjRl5dNIK5BuLRhe6q1GZ7ZbJINIxxJzRvs0Y
07zrzgrq/taHDpAhnULz0/LXwcxjRUVhwrx3//D89TH6YxRmKiijpFkSHM+wFk1GCmteF7YHD3mg
bBHqmIGPf0Aj2L63hHqP24dZvxhFG5GM8U4KTl1x8SYcWql9BF8KH4xBeC6upMRnE7ni19EYk7tb
e9cr9dLaftGa+KBa4ViFGMnobmwmIdUE6lqe+mdDdFZTiEkzMpESlTANXgbRMfeO0+DNiQ/jFFCB
PIgNzsVEPjYa0XfZzzZ3EKaaeqO2TCDtIlTEHbENisOpCw7YI/S75wIpzsLf+14IvK1prLXfO3Up
Lh4eYSKppEFWnEld93Z3YJWR7rCtJl9THNZniUPMSiEIoUqUiecBMkLQl/0eQKlf0zW1n4MY/ujC
8pS+m8QuDyMEvrABTv698xLAf4W16J3hMwibi2TGzehVcBCSjmUhTm/fULGJ7TlMM1HPvkFXwMi5
eYg9EM1u5LjEEjkfJm9fBu/yjBQYvYZLbmx4G2gQSHWQXhkTlQ26ve1oZvIdupRGsDfHe6ZO7e/4
gtBkSSOh2Lb70EFhmodDrInb+LsBps1MJ/vnggjGqQQ0SYrTSFziKhlgHf0HH6oU8YIbrDrxfgO1
sOHaypG/sYifH76QWYOZfgECQ4ABniZMqIo8Gk7W/2af4y/aMbDrVcKu/2ibzdsmg4TP1diWWQL4
E0w8sGzUvOglno4LIneAZtSkJvQKyT2QVHy/UtJyVYVBzPPeuA/bR+s4sxYjBYBLIKO1t3JIZS6L
DDOEEKO1naDGEGbaI47Svl3vuIAWGM7P0zcvJdWn6od+8EuUz0g3NAB9BHOW0/prduGkBrBos2hV
Jeypl5KW+VLyIP7g+1AcW30LREtMDUncieagJ5j1Wnzfdq99aombVRJ/xAxcuSAqWcchAy3aKHuV
h30pU5eajTWlHw1IRoqEP+28HaqMEgdr3M6hHBZCKEa96Ki6GJ1vJFBrHuCrPtK005r8xQ1kNfmB
EYlZYMA+v8434aGXo5dov8ZGKBddKAQRk/FUgBVyJuYdA+1au1jLJDsvh86ftHNoeUZhmfX4kYUG
khNL7QAVBz+LrvDQYFkV4ubPDIYRDCOuqqHSQ8FAgoejJntHu0gOUy1xNKe/52xDm4KMO0z2p258
Kp05C5FKajRV0ZgDvpuZ6WOU4tw98E9piDw2eDIEXHWh6JnbdFRRSfaGHLt5edhRR58rlSZ0vLSb
jIrnaIFtsil6jhopgHeAQ0bDP2bBeSeuDeqbc3+i1pse4/7sjG44xXtK/KDSnRd+c9Ttqf3F2MMf
LoX9tLg6zDuwg4/9UIB1VimOtpKn4qu3g8O0tlvc6cx0He7k1ZDa+bNkJ7CwRIfDQDRYxF+e8z6/
7nU1txJteh6UxJ5KtaM/fgk5FKuoQnF+tJi/1+3J5GqJVTiV1zbrGASRe1pJYlCyYEuXVjW+6XiG
537zJYh9CGPKEGf90uPIbB53Y0IV7cVABlMQGCzqQDu79q5XR2MIWPwaywvw1V8LcSm1FOH/xSmy
2AM3t2ZcQvxH4GJMohjt28xO8Sxdza1XqKzqhhP/YDlUuORLyY3AwnNyfO+FrURhO2Ac60UvQEhx
xpEq1PAicIVnpiclC+7t/ZKbg+0WDyI+23hECn6pmYz4FLgcjuTk/69izRo++t1fAmbL74WV2YnA
dGKH1gQIpQGWLV1GwQI3H6Gf6tO7NJIwMNoGwOO16ceE/Epc+Dvw+NcwDwzil7JbxHZkws6oWt3F
ALQdYqolVX3Aw1Elzf/of+A5NTWZYKyVyzGEup3W0vjHT4G7HyAOnVED17Tt19DgGDTk6fcua8YC
FLYBTLzxdlu5bcojJBHRN/tmIOO1Fu0ALUf2mM8fEQrF6o/kc1e7UcKYxjck+Iy6Ewy59ivdTOLf
XdE0VTI3z/9fgCxQ2ULxZZ/ci+q2MOwwdE9mtMpC1avduzrnsxVtYebHf37EvXKNLPnSImJq8+fI
sB2M5mj0dDmTeFKrQFzd5DxV4U1ltEsPb45T/7thCSUX/mWZs8iYOV5qPz2kUW2Qm08c5HLCvbvg
S9XCpoASRgzwHjocqloBla9I4DB7OI/UiFszRax7pPB82Qo2tciUqO6xg9w7vf/oZWFMAm4onsN2
rq2EAU2AflwI8ct6PUQiqcFbQpwyu0km+02gG77o2QhsJUdawkGjDfZQWOqJS1+NHZLrLVaUSYpU
qWBcrsCnQAsPI6pXq49l5FTfBAHlhy4C4hdtZmlJFv+0o234WY9EKRd/U7XTgD53Eje8IibO23A+
4uBjqtwSN8yWjA7S+J1eTqH1aktA8EBVSZ/S+T5mRQmia/JDNmTDYCy9X2Zn5wbdETUosL/3JD1k
kf7fAv0jQG7ieQ5YjMxQXgdpuaVJA0EUWANRa47SIJS1FgpiYqfSgwP0SW/R56cBP9RxrBw9Jvl2
6ctas649XAM/8WNmam/WkwaPnkjxwv7J41m+gM41mv8dOIjKrDcPVce5unKqGy1k0NzTSO27XHR5
FR5O4ZppaH/fVnsH0XZCjYvLvEAtny4Cbyu3P+6TUrw9rPgkeAgQm9Xk2kInvPQiUxAuz1j5HGYb
8MqeMT7IJOhFWJahjmr9NBMvZF8vGythiw4Z3sS9oi+R7vRRAs7m7tlUhZUNV+hR4hk3zTds5I4o
uDLKiSyZ/uD9dm3LEHlXomlE0iIoO89C5IX3jhYWVlIl3eLcnHzpB5S3tK+xJTAp1SBdPhzg8w+3
kCgaS2BfBHuSwV+0YRFH4hWSU/MTfpqhqIXo7yS9vmj4DIwTgAUMjEMSoesn9U2lzmNhnR9W+AZe
GyF1A6s4RpipuCKZOvTudtKG5SnhA0nijVY7oPutagTygg6g/1eUY/0TkL0cyq0Wr83PEZzeHKD5
O9kGq+73DIzOvHYhYbYEt96RZO96LIBOr6PNhcJRaHHMUtvz5boCMpuMMtAR1cL0uuyZ0mV96PFZ
StcVRA/C+VAO+g05HKh49PkJ5eP3H1ajcq1wKIf9ZzRHBuKJMKtFADK+shPMenyTFMdFL6DRJl6I
zBPj7B/E4kTf3+5xitLfwYMIq/qMCCeK7wjPmQ21P+7z/4KG6krUSSsWCsne55WTPel0fPRkvZ8O
tC1OyE2vX43syPilEnKBVNHtzKYFCx8jA7po0kVWS4VXMiZIZjRp7TB66ckFhh7HqWopzDjogYfS
BP9BOCmOesTdYZ1yBE15J2dT3MXr82Wnu9MMMXr7L68vCarue/mhqrnLw97cVy9vK42qKe7Jmw7Q
xb4dTwA5/IgcsUv+NlH7YtqqtXvca+Ka/Fxwx+Hcpe5AWOfn39gmm6h8EXDryA3tpCTNOZB6rHIs
ZBg2y3YwvnsN2AbPg64c5iHO6ALvStCosCkiprmzbNnDsLRvJb0/uadMVbsp/WqYObGE9xNn8Slg
2gT9BkHq5qMs3M0ZkP+5981vFpbBmVTr+yHMpKpEXX2A52IeyjJzw5NQfb/gDIuS4eSMrQr5GLuj
Gq4kJ6GzJwKL+sYg+IUk8rONizXFf//EXEjB62ypRuDv5/0sauP6zxI+MxVoi4cwJp8Mbwu+LER2
/5XS1sV9uWfR4ZJO7LBHSUUc1Rbaq1nYsTux83mk0CRV9rD5bFGSupD7mw/u05zqDs0+1SAihH/2
/zyCIfJtr11+rILpDJt8VQap1UzYHAFSO9w4Jrp0dVrYCyQJ7T0su69g3wcNQ2EpUAudxFpa3Dm1
ggWJ9r0OJHR4fUY0Xx4SOuRRgu/7UbLqUHDXYAWlq9Ek/GndZlTWL1TT0yBkRre11Cw28YoWMkVT
94Zru8UOLFf8ZLQUKBBqi29nJU2D6Phqp682ErZW01gLlouIZEknRQQFKWi/QgGLj/qVGIuyAAHI
qBoiTVav9Up9JYguUTexIZEU2XMav9RCgUCwfoV2d59cO+e75UtkEVuY6AALaAiJTNkCq3faapCK
2SnDhSJ6wz6Pw48joDtDwWSuOGQpdo+zW5XJad14veyU5DuayE5ghCapTEnybpV0DGK5V5W31S5S
H49vvW3T9W//mtItc0tWobBOyw79TWveYqfdeJC7rNDyCLYfpJNV8EZQqowufjIfFH9CCauclmQB
5oTBENomIcybUIEkOebq4ILud0RQgB+1VL4RYEXrRRDEIsLFkIbbBnScEqxW5b4McOm3G+kUKUEb
o6Fw0v9j0faVYwQO5FpB7LoDBusH50gVUm5qhnvbavGbguNTft6O+VQRaAj4irVq7ZVtbOUIJhSB
c6dYyRzjNS2Q1OpHrhNvNZe+Xgxgwr4h8R5nqOOJ5nd3XoCUQt/Uw+VMu+WmAcdU5gFhNfZJgFnZ
hz6j/0wUDLQdvkyQryWF4+1fhttCy+wAotWi81iATfNJcSM/vIpWjzIL0b/Tv5Dj+4sevIp1OV/o
/4zjZmR0CVn3puuDyV4PIyrt1I/FwZ3LRZyalrICgi3e3/sbLRxaaHvFvvIagQP6Z8vvXDiIFZGC
U98cV4qOw6cpcbJ1/66ZjTCqzjNAPBV1h71SUEykvo2UwxGaFTp07OtYilAWTGjEXh7Sksxyb8Sf
H2uTCLeydpmF9LNzl+dWp5dc7GQPZXDfB0zYSMZTLkwKfX0GC2RKC1ibB81dTQ2/mYaOAlHIBbez
NGZpGIuXyyByAS0ZrQqNvmda0Egiushbnf6aBflq0PRAAZuUbNow4dDUndRUTcSVG4szdMR26IKr
4rcqO0sQWHEU69JkgW6umj18ljhV/l92nuKrPgIhoqmUKKAXzwCNmjH6C5IADi307bv9jzJDojAo
QfqR6ID/RM0DvgEIgoc3ofi00L46hlxggbwepW/SEIsz+ORmd4XRXEUTeSoY/KLrJ2LncQDbgDAI
ezqTpJlbWrs68jSpoVlpwVcMUY4ybGX5it8riX060hRzPiIR4RbGzAJAb1lyHfMEvL/PDfcebPh1
rGMGoJHehyUXkYPP6GB8SYoaE/tPVmJQwK2dHXOo9A/sOMLJyqqX40HTN9GN5OnnGW7ybcE3Ut0w
hvKvXLpcmibzp2ZPMTsHg0VNtpcsEP3RyOHYlNT+Fd/LqYWbMnskz1ib0TWbBAHBR2u8SAQs18UT
7BT/hvDZHL+crvDsBRqVTorBcMIsKuDB+bDHF25lVVcjBHoVkjm1gmmRqX6fLDXzaPeiCjBoC3+O
oykl9Kh7rpTWoEBJ7WG6PdKduJw7GjNsPwOUD5Zr0YVa1qQmF6PL7g7KdQaGxeW1hLy0Hkkqfgj/
BKtLFPXIr4S7ANCaeQVLB55SlAPx5lIcc/FNioSoRR1NdBFr/a8rBiFK4rHbHFvrkY4vK/97dVcY
kxKeVjGKd1FTzWI7djYk/rYjAUeG7v/j7CRI1wwgGubFxA8mpTeISctGk8dYBksnloYPc7evm8Bk
hNd003pHukLQy4nK7x330eYGQkCrL54dJBKOkzEeGD/8fU+tGrXHSeq5NVX/qh2CuwLuw/A+VJhe
1KFAYnlZWbguqPeeTkLrKhslvqVqWP92NtQM2KgUYXJPywH4lVfi926mIEaNei1UlneIExRh7N+w
TlT/YR6SobYQ8zwqlP5ySoX7tHsQYRqD28Fl8tYV1gl9W3pwWCh1Ha/zjRWJnJDVUVmOWV208Bcy
SjAbVVyepfnIFcIYKcbRas28qEjqrSq1Lp+1NhEfY8PnbGzf1elEYFvUKrXY2L55ibImD2racFoQ
BHuyXI3tu89Q62Nf7FAxNuq3Ns9KMyeM4n17A3l52XhwIUhIiJLcZa4G48IYgmEbhcCQ5kiZYlTR
PtbXsX2FqeUaO5UtoH3H6Yz+YSvNZF3qsZVqV01H4GFQ/sr7KxF4LaVqDmftvZp1P57lsXl13rjX
VHrP01ELvUnoddMzEspk5f+4z5tT4ZtI5Pinl6pK6Xw9n8ufqVF+/qoUwSjgNotsTFWRcGILomo4
04GDQAvYpDDRDL0TlHLmrLdCR5vZ47v3bTMWFmfXpR/zmoEnWAfvsYc+ILHlYbFgwdN6b0ncIAW/
4/aBQokUNvzF6+V5okfBNLeh5OnI4a00yYAt/E52muR4OjmGSn8jNYs/ueVl2rcYruIuHf+Np1sf
ki7l6Qd2IPclJj7UIQ1KxGfGKyTa1oxeSrXFRYSFRgVCUiy3ZuTodHTw3ZbFu4v6SmI7dmBh0CVP
+tal3LgqwhqdCHHoTYRiwXpTknHKEQw8cxaUI0QqSFKk0ajjE5Hc3jDfERA/bCWgLJsRevDcv8py
m52/lzSPDbGKdnQW0ZTLnoyDrReAswVYd/WfwCFFvOgpIYsbhIvs7ObhNkm/QsfEgdPCjq2hQLcB
bNZpKMNMhdml2pny1PzFioDjB7TgMC7vknJJUZPdp+KYRkRUySeZ7wXDIJbltDVzlZVBZ7clp6PO
47LBnLBS4DdRijLRPpVDuKHEDmFIvC1uSljkm3HJyZ3ebCLH321n3qgCWNwOiFjpdNi+v1OnKZuo
uHQjHu+ko3Y8JEq1rM3C9e/tyKjTCGXsok6+3+Gs8VTArS1PQj8IukWLy32A5nBYjWuJ4fEj26p5
sEWgCfF78iMZlFZLcWfClgA51X4LCFnE0wZtAs9Epgil680nrpYo1Uj/clypfzUSWDhyTCf7prGR
M++DFQVFIbwU8B3+OjWV6FIi4gbW4stedZ8wWwDB3NS/XMEZIAa5Li5eRclPaWqoOAGb+13+PVMr
u0ggcz8EI6ESiEwg+rr5cRDOaVDj0lIbBfd4I7VW4oNkNP7g07CAZzAGXm6Nn6X00/xDRISeb0Iw
Y5vUWWkgH5/O7+ZY2xp1VM2tIcIjIUxqAKO6QofUy08/B5pEvh8BMh3NHxlYHBuNNpfiw43rUzRU
CB/rwW74xvhBoUxhWhas4u5Yl64apzFTerTYYOEQqAcjieD4YSFpBkwbzHEc97pwswqajSHC9upv
mBwNlDSUEdEaxQPGRuedsj5X0Xy+Biz4Q06xD1uprfwSxQmnDn0/G5usz4oV9CMdK8lcNVUDLBlk
fThZL4UkgX2qggKaMubVXPc9UXp9pJf7laXprkNf7AHxiVlALiWDM60yAsO9iKtFRIBEFJeOoHDY
UkxRrfpea1qN2/udGvHdZeEV/F5pW8eYw07PSmANqeo2qnOK6eeEWCa5zYzpfAXybvG+ESJnBi0B
ATKS/OueZMqFnmNL3I/lVC7RzEMaaL5cEPEfVkV2VKSWBC1zOn2M7p7MQSays8mMdPYTYdulpsGV
oquQ7Hu2FlAxkvo7M33ypIzWyoqsAkr7rdmLRmlRfVMUDSqXbymjS3bkgKyQcTYo/G7HLs7PbYi2
vX2kgEJR3H+wPW83l0Jxe/60cJt4Ruft7fro/IFz5kX3pEKyVw/1DawDAjz8l/IPqsgE61a8MiQB
knjq78biPlqalwdUCwmoxjmrVrwpFGZCnRm++rPJA9MnRLvFHj73saCOlUlYyx6+sPkiExg3y+oe
2U4f8qGgOX6tNYmnRoPotstoCzAJDL9+GdNbo+H0djyGayXcTXcsW2IlX4L4lkJUmsrvPOtW2czv
1/etnJLsq0x0yc2KEOmfUVO4HhILux8nYnfBlDWrWgxIZvjT0uDEI2e5PfmPiQFJ6C9A7jDNjKvE
jfqCIJgcFEKMpu+9R6vkmH4DizV7h5TOKaPUBRS6vtwI8w5fSfXiYG0REVrEJ7xmg/siICJR9RJH
2JXxT19ae+BcVszxSO6BXlPWJ6RBsROshTcIp/q4LdnssbReME1yncxRBtiqLxxVc5oICv3IrLPu
hsNlNbCnVyy3lBaM3824AkWUuP8uTs0hGEer56dxXn5Swev/5w1d0zHqPaFCUsdU0HdS9gFXEGoP
qQm2NdJb5V/o4CPs3EUl6klNWxHeTQ2Zcw9gGNMNQ4EbtIUKTuc1bZ2v8Ck3o1GaByqVRNGN2+oo
qYV0X2IpRtkOAWGhzYqJ3CMqL2kpXgz0+AmMUH6KV75AlvUiFQnldh9dmSVkyEcz3ppAIzGh3BRO
7yqO9yghSY1voI3C4Lf580vqt746ot5Ua6r2vL10XRAW9gBC5hb+DvycYZlmQiYkOT3QecDkNr0m
cd1bDGsmE/J8EQ4aoklvCcGaBRe6twAw+WBFOr/Ip3mc0a8X3oIciZzug2rclnt4COlLdf67Z3eA
2BikZtajMYesmw5UQ4iyn2tsLyHWZHhavk1IwbBV+82p3LtA2YDt+hABsyVYvihJ3o0nsIbb290w
eSDze5vNv6vfG87TLkbi6ytrHnjd/uStXwwg9hJcDMSioZ3oNNMKK1CYvnkr0WjjXs/BD84qrNPg
0w5kVYHjjfVZnm8LsIShsv6PL3F+U841qI1F+TnR90KnwCJs6KjDk/Kb1ymEivxvRXoE6fyoKqPX
AiYIEGFgU88K0hYLxMslHVzdtLyrK/q05N7ShajF277Tf0cEzHzgIcZDTCkhACDmSbJPsbNE8C5g
YGKiH0+/q+ojedk+X27oKEAgoxUY01aegPFuMrv0MiIM8fSo+pdK00aWyPXBbC/P1AE5Qi54jxrM
PoZittIimR0BsNq1en+V69c8Y0ARAapEaEZFmIqc5Z0oVuZ/v/16JCcPbdORy9LqiMhLFX5Is9Xp
dWlOOnU/J+zcp/7HYUvwLraA0PUhJt1To+9gOdaRtYF+ivE8CgicA3JXRKizWROgZJ9v4VLAdIyP
H8MtOJGQzSQm0UKTCvzFs8xBzcq+I8KXNZcKoCBzVtDvVNDj3gNbKBOOTDtJfZr8GLWjtmo+H0aA
gh/gQesi1IgZ61R9kL/wEAgsPLAsG/HKuIpDJ2ILwRZQ+4PJYRDj87PYTrpEUVWgoBsKKdXtMJ5T
quouWz1IILPV+jJiJ/LSG3XJ+7BFO7VZB+Jc3r2ICDwJMpWu1MbZrjbtxb3V06orbUI0QSXTa61r
pnRpgaWbek9vQIxvZK0QIylgLekO+RUBJv2qYdsAw2LAwZjBXz6ljBof01otCO/BfhaHu1ZRrpM+
NbmR3hky0SBbOq2WiWCby3n45YCRq9qu/aPL9rCB7cpWqTwqvT3T7fE3iE/3nFcp5vY1keUGlvE1
Tg7/EHf1fxooyaEur2RzVgNlMC72QS5lGUkmkc0bqtIrfOtZ7srozmUwFdto6Bh2EcNIPyHMG9G9
MzX0rwC9aF8d5QLqKBEYWa2GIxiorSYTZf+atad7UE9QG4XAsmb3uiO50mq13m9XPxSUZbV6WaFX
Akog4PL7cBmLNKiPKHhL/EyE6QJYZOjV32gOBTL/pinysdcU3J+4dX+Qzp3o1ze4Q8/tlCcVSpUK
l8hcr6Hp5ZMXQNK6E0sCrXXvL6HHjoH+Nko42EwRitSp78OJ+333vyvq6P3qFtntYw7xlar1yjoZ
VXvM9p3Yrka1O/C7BfhhHs+OUkmai1mLQ5vK4y3jM9uMUUlg9zgboQWZqnjncSmKG0NwRxb2NQqn
IOffm5gpJx79y+nyt80lXxpMlMCeuO31UJV+2jIcPiWs9vXqGn73nI0M0OtL9GGuBQQzxC+EXSeS
gW+EMCxtqU/v2aJFlTjx1CRLmaWDy2Oo8EFLynaqx2Yy0a+Nz2Jecn/PWV+yykO+Q1YT7rthmF0b
jZLYtZ7tDnpPtI0/NbblS/KaPnBShPKuN8485YxfBUPgpa05GHl+EfXzd56Q9W503n73r88H/bgZ
QlyZA5cy4hKMfFZ9CDzjDqye4jgr8pupCS0WyO9m0L4eOWJAixyv2o+eY9Jg+RXsoU8iytIezpfM
W/n2j2f5DM4F1W8/f2WJ8fI0zPepPBV+EcroB+cpUo1ufMDYGsRENOnN8TaT+2pDMFXtrti9osqQ
FXfVisBlQFpyp7tYFXAlQppqJ9Cd8Vsk9NSpIw7IenCO2J0wZGmvi9tycxRdJvFv9w5rfFbRV5mo
/NsUoRLpkyKvUyizK6+3ufLZbVf8ZLtA/0A+awSyfJ0dFZJUwQwYgeR7eKXOBJzZK+TnfoLyhpXw
OuLNl7zZMaRYZTQOPSsPgSaJY1QlJdUtMpkYn87N/kIYlwTyN1VD2EQRGTh2m3iMCnglv6uEvBfD
9HkJda4IL6QbE/+Z+zcJfLfn3w8h1ZynTUEI9ZnBUqloBneib4TQ/PJZLy06y/pj0fDAs4XdZepK
DwhNBmjc06uAjKLpsXNdOd9ivEbOnoQpfkZauDorrMQxusRwbjZQMZ7GAMAD1DSmPb82opa1G2Ws
v0Sb9tij4afQEB8j6nSIM0uvd51ecWcNyOgyER1J9zUqa3L4gW1k/64y03aNw4A1dmc+zBnzzc7C
2jPGQ0FBZ2hRURRkDeJcPy9Lh8U4O6W3HwO07HinnFPWHw3MhAsOYd6zuiqpSm9oCFWfOL3jXmA7
YLOsdvspkQzP/TVj0c1P2lcCFOZLTjcPm+2lzV8es1uBokL/KB67CDUd7jAwvgUefgwVaokqFjPu
aU3mofELwAaAHZoS1/gx/vFi9qhQ6L5pleHE8fRKgviDO0O2PbaQN+0DSfvM9pBrIr+/7CCspCiX
gIGv/j6JLG7yVuGexp6tb30X22iP5Z3+vFTu4KnQVj1tsWj59eKNQVLd97ld3CECcZKeDwTg3OSd
LCcqC0AFNuHy4pCTe1RdsA/5F+Xrjl1iv313YU8lAgVqqPk7fVi0oHzTPIBIyhOfNSUOAOrUnoAb
JZYBcfDhbRMzFTfBwUHR/VXq9SUAiRFRzcHyLmQYrJEE2xg5rrZ+cuS/+K8vNLd+hT9iAKzc1qfz
uDtBNp/CFQBTix2p6H9/0lt2EPOSr4umHGpRABAhcRKbUbwGFzp9Z7mWhIoCOLRTnPWiQwbR8cU0
eFE21CoFupotkLJxrjAtbNunLiv0keQ5LJ4SjrVkuli/9xrKCiukaOXbc1td/xMMZXZFHkRbMxSy
dGrZUtnc1am3Xz4FeLZm5ZrcoFp75nAa0arvvCY2Gic1fr+HGGUChV2EhK6WWb/juK59ZY3gaY3d
SxHOM9xpxqJiX1KNQpj9wnNGD9F455NWk1Ai1+a24CnvRb2//gw1VWwc6OtgcWY+WdjxDnu0e8+R
VNH3teNV5kOiVt4kqvoHqnCDy11U3/iPbU8MUvLQ6q2/u6VpkzTCgUBn/LEe31H2fkURjeKG0FWn
xB76UhdntNtq8zWFWm3GnQa4BTsdWaIhHebVdHwU3QBysIUWYrQ7tXavfRjnzfoXB2Ervuh1/TJd
CtOikOowzwamMOUWmn+0egdwoa9zeYTze/4d9cEKiSCSYIs/HmGWwSPrjLYaXjmW2tf9OdDDEnc3
POE4+tQgMXgY3fl72j/pzCmhXMOwJJLPIktsA5NRLEPn2BnaWWUed+esvm6oBKyIlUpo1tKvhe+u
ILdJVGHEuBw7Jvz57Px2N4CLEB4aehbq93Hh599rEyTHKpc8nMqgh4oQuXOde7bR0j6tH/R9sxVO
ukocW6ipxAnrlb2BVbGFWJISZhVWPIJEpsoHXEFUV691ZCc4gdz9BpNj4GXRaj7uYTSzGw3RPilg
GxHlVhV9H3NG3qoXjdLI/jMKOpxpJgtKTBB6j0zGdU3dOO8A6MrtEKJUXztFpRPH3oyW9v59GWZS
kMC9EDdz4MT9IaRWSpMuRqfjs4F3vT53Gfexk33IMZTLi0/zJHIsRcG6aAj6hPJj3qCDN3s+4yCA
lsKQeuiozo5wOiTpLduRSttoLi5i96nkx60tLb49RHBfwwLNOGl5bWU/6rPzzQebgnjIFgdCoccS
aIre5uS72sA4KCHL81lyjfUZ3zD+x6oI7RH9ExVgM4QG8IVsB1JlI6K86JI9LpQqgqCCgWnp6hfS
ZNosrmbxonVge4ZgmCBXf9vUarezWsBF+ruTYefoowBhxngrCIYEjm89jQ5aIkseQMMyOvBGLFP3
yX6Rz7msd0Dt1JM+tWGd/mOCl2c4mgZAuI+8v2uELAaM92Ab5lOb+tR80LMBYRDRwKohfVRL965y
Qh8AmzBi7z2UN/ch11J/asAoNvfiRMlzKMxzfYYNN7lLMCR3IGCdxAn9zSB99/1SRB4ulbKnguBX
MTr3K28S4rmzd5CLRtyfTahlOj+3BGE25ze3/L0+QPXQx7dy+JoipMrHn2bj8VJ3C7JoEpW0W4H4
dzuBoDCNY/BMQwx0Jdt0Hok89/98azNvupKolLu46lGkidJaXCPFyXVsIN/YIHmQll/oEeZxZfNd
/EdOW7rkC/BuhCPfUwfBLp43q4oJLSJ1R3gYouHCC5XJ4KcU8fdQX+bFwYU04lKrdjQhZFE6j1pI
biqw6rVmM1vfvxXdIb1UGsi3VgIOpDDsTCSajCAZPxUo/oy1/DEOikasaOKwuUYRIl/MUdNUBume
4yxaYdokZNR1rErQ15Q9f0Wrhg3AQDkkG1ubG91HX03iL1AmIX0U4S7DuohWmHM8KJ8oNvPwIhWK
dzj0VJu4ID1vLBdYrg8J7l+zYOSanaWzV7v2LrNCGeU7J9EGzmTistAdc5ANF1Ck50zgqH6e3KjS
MJm/Ru5m7+BuFqcp4dxk7d+Dd+kmsUlAcZnFZNeJNKMNhxIGyx/VOt5+uxvTJwzfNZydC2Ph8zKU
Garm+OoUhfK3wGlH8zAVxWAqoSXWXTAw51Lp3w+dmumilqXV/Jimw/GQVaPwSbRtFU5RDfxR6oMk
4P4mm7sHlXg0HLjl+mLhNaeYbEsjqjUm84cTg9YEvfq7fHlW4MGaQE2moQh5XxlfyviSXWltZvga
+i9NG7AFa1BCE6Vxw2SqJf2rhHkYWoKSE2xXc6GspcCq/60773Dei3rjSGkEBSvidFrD9RiJZTCI
uUU3NZx8wOPfJIoLqwMxy+rit2QRKDRXKnizPLpMdQbH/d9uaGe/HiHQJeUvgJ+Y0Mvx+GgcDPzU
+LJvtBaAMyHdue1ihPmismqVxoiwXuaY5NIRP8KWcDo6jH9hAEuKQhkrd3dVB2uPPGlfgaa+2bAo
wME8swmPKzyFnYWWY5jokW0F8nwdYxr+dzLzQUwNVPx1dhuPVaDCji91x7L+Xup4xusVVSd60uGE
4n9O80TAGoY4WlARReXVTHBVBSGOL9/6r92d3YNE8fxcJIF6NIKTfzWMh793C+X1p8bTjM+aGIzJ
ePWgXS/lMNcCQE3ct1DgVb3eyiINK0C0CGCNb7hJqJSAM7t2t/fuowjUyJLODzoe57KVuneDye0r
xQDhGAvCSPQL7Jch6cI4o2Q68jZuq83xgLEGE3h+z2pUyVwqav/ArhTAQOrNey/tImw/cSHlXnKz
07oqjkdbF3a2A4giPY+1+vKa8kame7IIptUnU2bQ5dlLlpItw714HrEezt10Ec0RgxqNEJE9JTWi
a9ttb2g10FD80ZOrUwT5/jm3oGC++g9wiQd3Lq2yU9qqSmugKml1zhHPD6jLnIKclSsTCwNGFKTu
NwYdXL9GzSygZeyMQGOmHuyK9mma0GngEUyM6Vzy3hB68CwIbHADO7er9EQZNCC4lDjfw4/iQvu9
zHuyYWC9IUavUYzsTZJb1gM5UXLJwFhUsE8Hb7EAz69bAEwx7vsxJTZ/raUUe/wgRrtSQd3Pmh1w
YIBu7gPNPX1jCTq/gEkBieeEXLOngHw53CsUhgUeCFm74A1udfIUMt6gSuu8A3UJW1QOpIIXU/wa
iNFivITNbKw2dNA/yuwaczyFNNfEP3SWIDYwTK+E0SXbsh2jY9W7Cik7FJk5/I0k6e4ghZT/oe3a
p4Gy2akN2pFoCz9I9Y4AnQH5ZjQ1vmMzF2ftWBP3geivtXcJ6hDN6PMlegiYPo6fhsSbfSus147V
44ePZj+ypXU15zG1byZ6qlzjVK+PbzOzAaXuqsimE3sNLAuoNEptdFp5vef9TenJumx4/9B99em2
eifKxzw1XgbBQwelttQcuQmHQcv1ycrsqx8HCWOVE3Hl6876ocxKrVWHVp/D4+QoOcUwDmaDO0ab
qPp4M/+5LFUNAAzf3BD4kN4tgl/lQdEb9qjorbXqQRQzEuK7vWBKcMFZYA/wM/Xmknl6RIPdXZRZ
8TDx179Kop+KnhvasdVDTHT8FzH9BpmqHDrF9LNkCf7LjTnRwENGqRxdwWoajIy64rNF5ZPB/3ta
tO9ubSrKgxXRGWUwDLYOVAQh8lvSsc4eDODkiMbzx+nIRA2oFra4TrJ3tGfhQGE0q0Pfsd5FbtEP
0e0BFNIYHZ5lFEsC251Xqsridp28MUgxeIkCcgGuebrirW5JgcMepCbkgN8yEmyO+QDrvBlYxJHp
ogVqtG6O/UMNrtxTTAPVpvxcF/M73c5m4sN2GyqV1Nf5u5lgG974mxstVNGq52FmvRSkad0qCYkx
5IZPHu+Q9TUeEejwFaIahSdk57HttbczDLh/Di/0uyTMJ6M8mkZ4KtFMYqcF4f3ifRAaYq9JDtCl
UMnBd2A6FNnoft0UF0IE52tc+iKvNGRweQsTp8vkg5jwehOUnY0erRxCno4RA1poyjZoLka9Jscf
p4vj81WVDiYiIw4gscLrv0yvaFWI9sh44W+A8l82BZZvTkIpNXrFrWlcvb7WQqh7gWA9YbVFeUSu
Vnq+qtFvtjRcWGwFERRManyp79IpmP6gQ7WCWe0lGfzr9XhTXMKAoOXHkaVdd+yLrF5+CnLBnVqJ
PSJmhds4rAgJnlbWInAT+B+cDUmPR3Bb3S20SbaiGPZ+DvVc4ZwBpmmEHH4ay46PAPmLMghVH5VK
Xzsa/GCFJAFxd0vP/d5kiO3EMYzVtRJXDITRL6s71eSfWCDCxocOUbFbCccF3JZeo39677WsUDeP
AOmgmwYsSmLOaM/cL1+L5u/gZAU10dCLwTPrmUjSy7x070UWpiGAC5AdsaRZ4HBLZ4E5IHwJWH9t
ya++JRyOEWHTjPhZYSp2yvG/stkA3woTlxMsRXnSml6E5HqFg1vm6KAjEDqzdXXj/uZKZQV9vOdH
PzCtnQjquI/gO6m8EeKh+lJpHdIZ6cDkV67kAS81gVtcNtQTY4QtQBdRF2TgjrSrCw2F42LVn6da
5NDVv/6GerWSuZ5UAhmL8tYehBsRtJ33T2153CtZayY77GHidIAUYKip4ycUaYdd8VrjCZX+K0oi
FkPC+XfgamttLPcsGxXuuRjT7zWgjHLpp1U6a80fAOFtkIROk8rW/t4OMYesNhj1oRX6naKCHdwq
NXQnNpKPvps0bUbapcGTV91uE/+PtTJY3paThPapBKSSoiaMe5F47UNPi7qrrekgd0OkvJt+kjc4
ZreGTS7wtYhzZYt3yy6sK/NG6GtZjyUseKcobmlCTbO/hZmejPTr1H7XwflTie6MmOvdxmArARKu
w1rOMgt4Y2Q2pr9BcZIlYC2dmcKFZBCf0W31BUHUHAeVBQNpRNCFHjNoea73955iaPgf6VyH+tS0
I6ZxP8BFg5NmF9IbdWcm/ugB7VaLwRvDCMVi0cB5HHvFKBP/QlT18RgVimLuYC76QBJHw73XVaYj
Pur4DN6TXGMPmsMAiktU1Ydj2PmSWC9SWnWNoXiI0BHd1LdTwYlSRcAuf9M19AWa3dbfPsPwbT2i
0EU/40fymXwuNvbcsNniAHYmBmDZr8erxPHpoOcWue/B9f0fzO9L38ZA3xPnfVqAreyWTeJygC+d
kug66BpCJ0sFMyXrqwXr2PVMhkGZUvt3BeObcP4GvzgQT0PgkAgQ/QFhdUqcOOJdLT87K5CAgvMa
hW9skThChV/wu1LAnpvZPUfB1wOJwsPdJ/moN5pakHFjyKql2ZkXa+nohbie3g/K2PiGfpHKPt7H
kMRgwDM66LNvWkyJg30hrrKYptXfEgYjCXxmI9Hux83UgHpocOhaBKtj3mSd8sMxd53EBvNwBTzw
uiLw3x9LKg+6yUHnJeunpGbZ4glV8gq8x530ddIMR3lGHaBavZWzUQizVtwQzuw6VgQTqrO1UROu
VufsJJEXPVmtfW97ePLS8qbn3LiaokGdtKkbLoCPmJIrqVNQLeHziaursP9igoFTiEZttLc3pK6N
2onRKscXscI3pyIFC2rBxw8p+dMbHxxbP75GBf8gsFEWVdjR9+0QC5q2JWN35SmExuUAD0lHvENn
S3ODWH5yb9vtE+fHPK5vlV31ipKflCqA5Je+QLJyP0kfBng75cKd2AHnIffQ38c6R0NsKYyBWmWP
7S9ITlgdOWYk6N0raqkNVavzYSqwGf92lofhFzOvQyt6QKdpQy8p2RZ9x20yWODMawRqoDXUQBsd
W0f7v2oJslowYv8g9rPYRKuLXcXD/Qhc5fnEt/XhqvZnM/iRRhiPqx+0h26uScMCDADL8S8umcC+
WZBaLZe1eX1n09tprICSnT7d/YZ5M6is1xp4yy9lSGye5A/3vHU0wCbEprBxFxqLdv3B7TMznqIC
rd85Y/7pHcpepgL3R+20pUKJVQeLqR3SBO0rtO7TTiNE2zXnhK1yQ2de8MwIsVXEn8cguV9D3af9
8gLt04WQEwYCLEswKhvJBq/P/+yDoWBoVPqa8cmowdaylUixVU8BjZh0mlHztAeDzZjR/k09tx8N
BnUbH6N5DxMrz0WQgZ5NJk3Xyp1kk54socYAyJEVJCWJPjZHa4WjJFp4DWJ/DNKMEuOg0dL9W+Q7
gFpypBWNR6unAt6SKhgJVdVLqyTvom1iHECRQ6BLQZytmL7Mbn2kAmA0Ncqy5b2Kdfp2Wx8RGxBQ
x/EjCIxIZEETfYFm6fClKHxLO8Qf009nWQ3O/3HtuRORoOgbqyfawI6OqUBbgjiP9G6s7GcmCj3p
fBC56j4/wUHmFgjId6FYFb+yrOTwK72A1c4dn+VKnNgyZNXfUr6Zl/K+NXPr9XFsGN62JURoAoWj
Oji1SI8/wfuMNb7SoFYNJU2hgGzSLI40R1zWVODza9HnfrxRtsVMD1b+4wG21Rj36AA5S2eKxCdT
Yls1CFjWWTJl9gZiufzJbOCIvKTH5ec4Y2H5CeY83Kzqv4KK36gec6v4tuJWQDshdsch21A0c+Eu
kAi7X5BpwiEJyiM074iTBAi4db5m/5SSgX67Lvj0h35hTK30YafOgngk7hia1uer18ZgZ45GT+I0
WiVFuPm0chSZOZaQ+gNKOqY/u2VDOsdC9bKi8g+fzmx5TfXJmGAjI1fYf3KUo0up3yxZtSAnUyZK
4lBrC7adIWW7tP8UHRBCIxAN0azcpo92sDf8e4zImVMGr6gOKAt5ZUIt/JQp2CuZfvdB3a34Dki4
pmzmvV8hMlK4HRwwocfNlWaq3bdO/En5TJ0BlHxz0QoyQXhhuDpbPf6unjJ6ckgzfCH+5I+8o9gg
K1Q/zYzq/Jl244Gq/Hl47B+ebdZyXszHo202br7f/Wl2qM/QRTb6o4SOgSC8jTwcat/zOvZrZWPF
jSt1rLsR0TIkPEMG2lVKsr6IarwP+lU9kVZSxaD5hy1N8lpOoagHQ7Z8uQDqYC5poVG9WmDL3Rwr
OlOsFKHcUGrQJrmQ8izMlFvBLG5jtaPZE3qrVRTJBD9F+qyii/lPpv0kMVxhA4VFxxm+PrPKzRJN
Xw8nmrfJx/VSPtum5q3zkRU+mhwMcqD2icePLxBPWdlZLHBx1wj79vJxkrMp+5i1hqeUQRkBrI0e
AkI39APz9n9w5ylJE9x66rnr/SL3GLyfgGe7gjAJAfaJu+Y1lSrraRA74+LBbv3zHsigwhEn8xd3
0mAYaBQfgQQqbmSBlo76EW39xcf6+iG81elLNecUnvW0O1yPkVykVQhALW6pxVx/2W+8L7k1A0Yd
l/rFJXj47YfBr2ACymk8TR0A0Uek/7ChGq7tNN6kRf49J9u9eYsOiU7R68hGmEu2eHTYocb0BiLx
yiwIfWbMinML5W5zPJlSEJardX35WDWi/BZvvPn/XRoCjV0MzW8LorRfFQ64fMTS76m8uf9+nzdZ
tbwbBcBaWcx7u/NYHnvRCPm8994dd4ZMp95+EFP0UrKvTzyn3rXDr7D8ZKGAWdJRKAczmLhLGBxj
y7IrzhEhR0TzBC6FBlL3NjSV5Eb8vfQPUHf26dNnAotGoKNNcO6Nm8I/VbdJMxSuvQrLidjo2hrH
G+RPLkNZ4MsmjK/s9Vy5HGIokwb7i47izYtYJguqVCGjsZsAhPLVIldz9yJjaHlh05BrqFHqBgKl
dESB11g9wV0gmHHxhR/nMF7SR+mpac4zAAerQoXmT8P6uUkB4d+bPwfT/KwA47hYuuB7/qEp4jIp
hTTwLwWarxN0EjwKkBh4+ZZkiKdZe/bvY+gXFSGsUTPLHvb3+YiZB/YYkr8ufqERJN0NgW0TZKzu
L4fCGREArLavqq5FZEgRs203+X1Rk1ZGtyxu8Q9PP7lriSYyyN2ixbVUVSZs8HlkmaUEO0vUCApn
Zn/gQNo8QyMpceJA1ZRRRso54IUtYz1LhqG8IEkrzFZ8Sn1+TcigUXjIzl1l+KF9Ss4XNom7mycf
kq+snqjtCIL1d2QQe1rELKg8DLvomwhJiF2N8sv1H0PbMSqnYQZhcMZsH/I0XJRof+hqVRnMoFYb
9gBCUj0PyLNwMyaAjhTWWhKhDb0o3/Q5m4yk8xnM6LfaZGaT5bJ9TgOgDsAjISxPXTO+FGVBG6xQ
JXlrWXFvai0xrWEMMLb+vnyaPR4k83ykrcfg81bBUTzBPq4Z0A44MfW2ZbheaiOT6dikDB8RXVop
84rZNvVbDHYOGNPCbPREzxSb1iyjea0syZ1kwMV3Q+8DVlxbBLWczSQ7Jtt3y+NYiC/Byfi2dsKd
PdTsTUGbyTuqjZdXZmiXzohM3i1aEF4r0Hq4io1lyQ+oyEZbW/Pc5JIeLB4sd2b+rAq0p4kFGOeG
3pXajI1bRXxwqPNaVcWu4fMHnzScGmiAx8rb8gTz2PLoD7heN7tzgzEZ9Y229aPNEh7oBTFtv6OB
6GxhlAr5Rh9S7A7j4+8oqDK8sn0zxOHaBCSs7+johYuRtu7J1hscfsaJ96lvXXvKqOT+JsGMglwg
yEUpk8pNeC+76Z0e9rAAI7b3AFcjzDI1OOqhFaxAk15HPLqy84whNouWRyRMokrHebtAr9ZhXfhq
YkUO62sDwKmCMYz/wB4rR/auec6J0tWBgobJ6PMVPBScBUN4CHgKczUzlDEnwdeIGpwIxY/3Z6ej
aGzH+eg2iXVKCikSKt7NSAEbherXw9ru5oYBBLApIl3TzPfrIkDxRr7GpZ5V/ab4GnM6Oe330Fh5
gdsfZrP+/NnfJZ3K+76pVz00Twm1ytP3GQeM2FWGahzkLGUXnnZJoA2OBhiSu9eNARM5/uWyyJ8d
ELiEczNm7Lzl+9fwRC86R2/MiBmcu/OXyhqr3jrMzzGXRBKXGljZSVOcGcA+QSslWlS955eyKiXE
wOUnz6hu7442S815Cbld0JF/v2F6/1m8hASuIGYFruKp0Z3fvSqTHL62aEFUbycJhYaLTD4YO9Ud
muqu0RGXcqiyOhxnNQDwzxtre7PBCHO1pwsKAWVR+hrPpGqk03fvwPcFieMABrJz9u+hhxCnVOCU
ySr5a7ZCGOEkzbcZOKMh+O7TKJNBFIuvhYK4tcF2Tl5+dAnWwHlmR3JebeH71KMseVFz2BJrIHxF
9qgK4QFz8BH5gOw1vra7IJZmDukdihM3zA4EaK7UqznXn0yIpXYxYwGYE+G8UkzJPpebFHwJiziX
hv680jH+79GRIWIZsh1QqhVY0ErXUNo8KrB7Cr1Eidu259i6fZx5q3CPXJS2FGLMGPmSDauaQb25
JiPHj1bVLlh/S6vR/MAxySTZy7UooB5Rgmh4KfceY3CgYJC0c/r/DB/ZEv5yvzOysbOYPRUDgOO8
kjPWIAatG+UwMiFfuUdOVMrgecE/W1uz5Lftplv5L7ARhyaBVeOhVVeEkJeeMTqVrd3jvnKt188q
BHfQj8l7Cq6QNzHt3N6VkiDyXrHeLumkexGLAyd0c6P9iSbQkUt1E/0H6B1h0SxjGeo+EKSqmXaj
mD8w4f9tUDEz4HbpnaVsrjvtuqiM1cPvyoWdJ7DJxs1pXjQijxDay1jy140GYa9HkYjFgFk9/rHD
rKcFzA5N8OLfuXxb61weH7SZ+CCrfF+n8u4wbqdJMeAbU71Jxmr+1JjD9zOBKUZwOvGCxyekz+9H
CnV/U8zQkmbageZqWW6ruL2o22HxCE5B7Eiip1wCiXqbuLkeUTqwYkXlUVF4Y7OsCrNEyl4rTk0m
9YI/wty3WTeJBsYZ6IZ82Yy2IPdNuC21EjbXycKZ6XJwyPsSWdtmLzeHSx1lufMyahZxqJgRaidD
FbBa9WCRAafvK1rarwgsplT1LoEBHTJulKWw8S5lhR3h8hH7+jA/NVvQpzyajG5pru8F8KuFg9ws
XxFuGHkq6mopnFFC4HYjz/psEH6DxlDy1vYqUsrLOsY4gDDt4gcKdiSHKb4KAesw8wt7RhSTyyeN
5yPDagi2QjdEnLoFlCXrgpk3G77b/dS4aYHBXruuJPY8EfWRwjWNJUpZUDsMynHB1/QZpmucKHt7
YbaOlOjUYS7CLS4JxCJ32ZRyiV9SapkGKjPxnScNUq0NEJnS5SK7SG1RxzqIP9AZ77iFiBuw8rHq
ovSlcmUCYstYqNEy/8VFhLpCivof72wXw65a0oYAhz0JJIAeIGxrEMGpN+ypy8GoAJadIEQtahWC
HSlPTKguF3vhVCirNdKv8CLxZxSbowKE8VV3pGxa9eSIDluPITP9llfGM8TnY/klWLPZ3ogB/g5f
NU+iEnfdogiq1ttlDQGLF2oE1qREq3jHZ9uw+13vt1mspe6ho7fHZ8aAO4GiTpxrhd0LwiBXBAnp
qFVP1sT2DglkywRvZY1Qk0D0JJFBi1cG7fqkwV7ubJlvlhYDPZemJa9lvT74Q/OYw9HTc63wR/LC
Ej2BEQHCDgzuejK/dmK+Oa/NmqcRXrkOiOFLo+8v8Bm7IA+7AsPlOqdp62LyvSw+4tGHi7lAfM0F
XYjSLBhnow+b+ccg4/um0Ctcd67S7eWOEs/YI11+aPHwDeC4Q3Y5MOmpZ9xdACWi/PAAc83tHQYA
P6bzYdj0LsxqDoctbNL6g/AsPeMyXHqS+tzXFlVEYAQf6pAIq/JtXca4JEoJ0WUZhooe+FQf5bvX
NqTaOF0wxH+S57wAGAP/1eZ8ziLiwEXeA5hSh++rHJZtle3vixrLHl/jKP2zK+yD2iriIOlHlkIY
xcFfnM9fp6qETeSSzm3ChHJzsUB9VNQQyvltrft0tzX7i7l21yUjEBSmlF0iGM0YNsWy/k2lp9KB
+0fUeTdca0bdPyDt0mtcdU2AEDuxLf3PgWCIgrTDUG8mc2OCbrIfLw390cDhpLcHjb6W69iMeIrB
3P7DTYmxGCkVddthkan9hjp/L1AF5jpUazTLvJZTWtWujwsuXKnfXJfOYA3SQ5rs54J4A938c1jP
AUHUG11FNdvtSQlYx53YhPU6UurP1AEp8yCRqDWVIvdgcor7rtY8E2/p3HHFLO6OAJDU3TXLzhky
t+eW71fBWfcqvOKK8T9W41LWcv5atlFnDuVpMB4BJMxvbLouT2rRJRFKX1IAHXPorohZIlatPvnV
V5wRd6WKPdvHY4tpY2jdGl3nd5oDosy/i6D1aodGkotZ1EOP/yol/mNckNjigq0BsUJlo9t+6RR2
MARxXeibGgsIXrnWchArt1b5aiYubXFEMlDEgAMx+RB8eAW2IIz8dmzJZ6aXbk8eJImMAZ5U3iV2
kDL0rEbSPRWuxFgrnunIpqOsw9mG2MOhatTq1clQW6JjseBom8aFpSqSFQSXWQPiLEQzxVKx+hpH
w62OfqkksG4KXW8vxBihlAt28J1dY1X3T8zhyP2OW3qGX9ShTY4Dmbmhy9IEIvKMzFiPBqdnWKNt
hH0lx4x7Qp4wz8KoW3ap1MLQNtahiX4uBqikjYvBUlM64sAPn9E210xZf3Wo3dyv9eaq6NA3VcMG
XFZfq9IARBaVh0cS7vVKM610u5GvFjF1dIg3xHLvufib5N1IMYRh0tbUjzXEukMxoGGe5P1v7AJX
bnpa+NPgVJa0bk8gMKJQ7W22suGxFJmUhyAQnRg6yldocz9B8AtPYwrwwZZXjak9gEb8yLOvQHSH
S52/qdj5C0oX1VruKao0f3FBC8fGCSOHHHEwevvF7TDYazyKoWTtBKrG8lFlURgqvFLr+18zSguq
MgReqhpvPbeqRmhsSRBbJK36QSQnTGuksWpf0635LK5/YyypdZUwuYNVS/xeEUkIvKdpNRZqeYGo
D2RygZ47KoP13zqmk6IN3H2DrwllSuUP2AU/E1mlmfFyw8Zz0dZ1srCchcf85EdVhN8FF0DxcE+L
8vWsgJbkPmAwOIxc2x4Iuzzb/3rCuBycDSN7jsWuxzpY6U2Re1bNLS0SfvKMODr48cBUSTh4xQeb
Tuh+L9dQTmLg2kdFiL7G71PjSoUZq4nwsZjf+/9DFfdgTvnFcTt88gYcMQkPMlkFc6teKjQ6MnRx
CJa31ZlXMstvuCFG207F3QUxUBx0dqIxFcPNSEsLFMBC78HT+9XN5QjprFx5J+prH6YvVEBXNcdr
kTJCT21jS4pSNOp/4z+WKRD9HyUoCNuK7vSBpVmVPYZfv61mvJYwQgSIcrfzNUcR5lNuptWPFFmx
HQkM3FxIs31tWOLjECaKUZGSsWTI9Mf+FtlLqjbbI6h2IEZvZ9+xys6tIhTLZQNTGXJ+S1ypuJuI
vf0OBzAu+K0T5Hck9kz4TcqqoU5JbtLf0q+HYb/BPu7UNqPq+I3UMaNXuRcAaVDqVmIzzgdCIdK8
Pc7ST3Hjdac3WTkkyqV7mrzX7DRS56nxT4Bk/Snya4vKzMcJO5Eh4SU12TKO8Vju2tbLd7Xgzozv
tG+Un2JTNvoZpMmkuaenZFybjCp9r+Nx9C97rhYEEcBQNmErtLgUIJd+QQgAhZb9AqzWK4/ieQaW
R+tcvv37dtADxur8VooZ9w+Vf9OJGkrGW9OLg0BVoUBlEyk31aDavSrp8Thux5VEKtESUitSDyKv
5rF3JeMdHU3702lBm6Sjq2oNaGCEM2PxwX4WnHQL3iCTEWq3RAlZvD8Ru44uM7Q7hs3M+esLccaC
zsQVSQ+UCzHqY4BOqZ4GigUlbotdGF4JHe4IDZL38ihB5IvU76BjzyO/DYg7DJUFI9oITDoZBY4v
jJF8Ya3FFU5DZDInEFbJAKfzk8d6UJvWRtyEVWUNX+w41iiZWU6QJ/4vbTc1BEQe9eASVOnC7cIW
acuQtGTbRCdDoeYtku02Z71meXUZEbDXea1ztk/8UVzyalWfewGG6IHMASueSSZM1R7r0/ng33OD
F38RhNwgM+HkKmsY88TBq53tuBzfWOC+fSr9ANtkM167fA70fZwahz1zgGjVx9wTjd/Q34GZjIHI
2hL/QEsDiy4NSUen0TGngqqpWcHY3b2NbWGrp2U7iQAxRXH6yy5LhZSoohVp2vptz2UbkoRSWy60
Qq5sDon2GS7NALpyycSNn1i9BjtGqqi4E/s2HKj1xIDE2BLyKk/0DVufEakFw3yHgkm2Nh/4ka4n
9OrgZ3N+Ad7oVA2zEEPGfmxardrtXdv+B4w+gAl6NZOzfdECo6b+Gzx0xj4ZzYCpG7o5Az//0/F8
Uw/SBzVR3r9jY+Xc4MbZnJkMQfu8+NVkd6zXR2fi17VEqkOeVuCxYw9IuVtCN8UDjKxcRuk/MYfk
royBkC00gQh5rf375gFX4ZLKHQEDQjJ7vnzGlTC4vHE9EdywbLiZqsCPfPnwHKEEXTzchpAlqwVv
JJDsv4vHPTSmUOqZpCeMDYDcy0/1kxYc3pP/WaNr+wZov5bV/PHgpmRfvM93uoeZgCq6wJKugdBb
ShtJU5BMn73SgDaMs75+uKQ1dA4fUmf7U8VmdBY0r506THGWKkpsH9PZyK0+/NZi5OuuG3dhxRnS
DvYd1/S4Yh9+KVYQAz22qRjb7cyGKNY1pth5AvqeFSCc6g8k+Zi0h0f88LltTPYsKbbI9QihJnm3
DFyYDGBJROtskE0gZmDAQjTeLvNv8YGGD8XsnnyULeE9DCEEh0KK1+y0+CurXNvbJ/oQxe7wZfw5
p71sNY2VcESwd8kh659u7qghL6MYhKzTVybNrVhdw3Ns4JPcGjyfde43JODifDFC9WIlzeSzT7RF
TCovHnASoQ2RK8TdzVJgGstYMLKALPmQyhg3xwG6nyabT56hK9Ei8Pft+1sXXjt9Tm4t1gNYjaCm
3RYpxMn6TJWayWw0KLNQ1jhxg9/n0135AATYT/VeIKfAIXu5lW31hnf/hegML04ri40ygs3Zjgzz
h8cIwAhUkI1Q4RqRIGLRMAtKbkcNR+zYztyGoKe+z724CiFhRuk+rGGqJdyL1zDB9WtSYjc0frSn
hwk2OlwQhuktCmPiFPm9QHoDXxSmp6uBpjuMdd2KFFb6OVDxgEClQN0++DL13e4Wo0H9YLynsqTA
ll6PmEugT+hPrbUBlcUF4+rrtV51tIyfm6t/hnQZ6z/lETd82FX26tLwX5CQHG7fDX/B/s4ZQ6v4
44ZJsw1GpIIfwvNOE/jY5XVlf4CBizQ7rl/XZtyUfBXTOkFTKhK2QIzF3FkJbvJjEww+fYv4xJVD
gQUkuiIEEtA+nvDu4Le0F+ij+2xBvz4x6odPdX5drhnkfpT9BkstbREpsYwamFk1vxS8IEtGMSMj
S9EtKfeuEZgMVxNy5N+C3IqFjy/oYPsEdvOzmawmmyfZhd28rX88jMcf2BHkUPWz2PyM7crwvg2z
wmqIKM+sKfO48tWeREMmBWwg2U0R8uxUGn+Pf3N/y5y32KToLZyviudieo826suhoqOKNqqD8EzC
FbMNzueR10eXos1aMi2bNc9w9bS50VdisgF2oaEwtyIz51F9eVoT/tZ515OtQZc1esVgi2qiDAnL
2G8BwdYfeLF04nbmeuFegS6WzujJJ6OAzoghf4rzD2oyBCTm4W3cOIqyrd/niG4NgRxUTVB0ENB4
hHT+5e1MEWIgwLE/11//tU82NSwrcoqKTe8rL3G6JDL++Fv3oSUKxpD5KknF7fesaf3k1VuKPR9X
Zyh0siS2qIU67mbkqAcmCfLcn5xB8hKdvDToeD9/HbLIB+xjDguF4yhqpWVXZQXp4FhdJHWz+oYR
OTcj/dmTmCLgfrXqiZ6IBX1liVmRUd9lD7OUNoLGkWi/C7ycPP/UNzZBIExlisC4hpJlg8RWfudy
GzRu81m2vzoeF4TFswhOyhZMRtfh2ClkPta0Oci2X6y6Xk1gPFnogj5NMGvEkdDNbhYx+NlLzUwT
GwzbW2rakMm3XiAa+UM1UtBGIgE/hRyYZaepTHZ1wHpyd7Ss9QQu3hBxLB4F27GYlZvrtLFN6x0L
/7mN8rfnTLHxxLbFwJum8OoBQu0nJiAO2l5jFAQE4UnfYQaCn3Km5Zfm7jyVwtNeQnB/Ji3qvGz2
v+clQLyiVgLA+hIGBS7mu9SoLQ9icO9uX0SLaXxdTGWNiv/5HtiJ4DDor5yuRwFp/p9Uc3DlWZfL
H1OrRkxTOR91Eim4WOwvrjxhkQUq5CctPU6P8D5YY1/PwyxED8lCZQa8iyH5FY40fkdP3T8Cy48j
2o3bvOOFulGbDguEH87Og7Q3DwrOSC7myuujOrLHWOS8n3ugT6l0xCWUfEBjgptAm0FjaGHzWwZY
ttu8l1oY98sY4WaSaG3Yj4BCEG60hm7WlAQtMblQBXwS22WHIbVsESeTFtofI1Ty9RRv+xCv+UdP
Cea5bnWQW1Fpzy8OIqL2iQGH5UdUUQetttfl8O151Npx401hN5ED7HTX/nwnGxDRFmaIqGgLar+2
O0IQSWmxhAwWf61xyjLL+f/eYgkkRZXKCTpwZdd7phzKdLfe0Rllt2tXUuWnRXIGHSEsGhKsdHbD
I04+zSd5eN3iyYVU3pdTiJicTM0g65ppFh3/DCvkwEuRTWcJx/eR0D0rlxenCUrZ/Ec7BCQ4/nVh
UkLFkh+BM8dT0+rK5UAYoRBoz6yRSumz3QpE+HdVrMdRnSkpHYelVqBe9gQtdPGTLJW/jFESIHJT
qdxnydLlODRqjAvH6sni5DAVNxZLzhh9N420NDkcncphMFZ0Jax86Oy13eIW96gl8OE6E+ugIgbU
LpBke4vyoxjyvMFfolBRa7yFjLzKCwSw+YE9F36z+0QGsVzJFWrS62YuRnz0g27AK1oBEQjHr8An
HLggssVuOxA5zXBy2vvmWc+A8Ejwf2bPkLX2ZqiE8B5pUydNjuLLvCDYJ/aKPP+2QUZ++Z+eyXcG
tyr5xtH9g7Zwgxy8Eg2wSxvQ/8+mEVXG/Mdlm9VgZKHX25vzrD7s3T45s5dun6Zzj5w2uKOlK2w5
FSiU+TC1nKNfm/tHweRNMzGQfdaxWlRu1AUNQV0+jbSvtjS8IeER3LUZl8leDOKrEzaetvo0OGq/
1RchRiSFbPWcofZLxluvvcCn6Ttq2vWWBMbGfa0ovOCAwq/PMiV2tfJ8JgfQWphEihXoPjwTfNnR
ZY2BJGimaWhRqquzB6M9fO2pIgsE7TGPHR/gvp0iH3eY19N98VqqstofghZPJLoUH4danCInxwTz
j9XipPZcCugZ9/3FgJ9vHcdkYv4VQU+YMFHoFHBDL/4/c55TzPnPMR3SliDokeKcmMRDMGgDXZcr
UeU1qpvn9OZBeFbka4o9+LCIATp+s6q1jPvC+uxXjJi3z6CG07/7MnNBa7Lmj3ejGyR1iuk5FMpx
XXhzynJ9Tvb5KYLXY/Rob6d4ALZnMuVBS0FdsdxLHRHudXp6nqDLZ9UPPmWScqVj+d9e/0U+XKbz
xuqgiNJAy5n1rzQWut3jWXc/ypZnY49meiyOK2GCExVGCK4gFia9y7kEvAQKPoXjPUvKJ+6gq/gU
DYT/xgD+joIWKrdEveke/mB8zShM+KQ6YGu1+XjoguqWeGe0cmxJb3+Hbs5q7oY3Gb6g17uePAWD
0QgawcFV4n0tQolu/LcIhsS7QXcAl945Ka1PJFzpp2aye7QbLnygNYA5Vd1XCPtA/a3LvPrmfdAz
RpV5w9AnTlhs1eNJsM0rK8vcflil8PTJi7ZeU3UeRLzGditIihN2Wo6rRDA04d3w32+Cj3VNHNkK
24zmMNzktqFB4XgyAMcfYyVhWeYJWrNFiocdrOcJJsH1LXK8uEn8No9/hXQqIfaPvV9xOup6qo8g
q4FMbbMPXRjq4h6eJeUuPo7/Q+1KhrJ627W84U57TNLS+J+SXPIkf9+xqXQPRHdHxpiJh2UyWpB3
ssa/yoMCTGwS/43nkPBSFpoQVNnPNGjWYXr65E/dPUu1k0JSa9Ka4eaXUbN5pVhUhV/S5YO45/09
7+PqCGJRc1thYpv8tBYnLfe7IR1DL+K0uR3InTfk9YmUit/POw34asGte5Lh9OjRnALNmX5I9+iv
FudiqT3NyQNqOba2zqjQVt6KiOwbvm9IHoubBmn0k/wUcOKYui4gFY430OlFT0uvbNUxYS+Wrb29
mjj0DhcgkTmhpgwuvwz3p7TrE7Ry4SsNtflWRNwnHzr46QAGxvH386YtEHqqZbE+sJWwWGInzl0B
wohk4AVrNqNZXR+7LiAPnRMstT910xj0kAVXinGSHnF8BBYXu/Vv82r7ogLihEME8ybEJBkUNET0
Bm56zre1jS/CeKQoHAbd7i8x32lDaORwREql9Nc/RMWzIw747OLSVPPwj6oxWuO7NvUuK5r1tsNG
/+1kzrMi1V/6LUQ+WRz8IhOistDtcs0cecXM5f/6t/N0wtZYPOX2N5b9m8grGoCGcz5OaKhTshlz
5G824ddWJ444oB0xa7qHE0qaQH0SzM4nGEMddz1npgnouTfkshTYh4YAVVxxIij51m4cFG0MrWCR
OHzi6NDNk5IN/l2Ylcw+4GpwRlWdoIjbpSFy8dduQs7+1w5Zqc3Q5uI1+fxWdc3WtqDLnVccWy6o
i7rMHfDzODaMoKL/xoJ2OYMlnGWwUTDuO73eH29XddOKe8g1F1WA+T4UZyoX0++CyZRWGchRHXq5
KUpLB5eWFPkImPPY6oMX79AZ5OlZ+aycGo7hTnphl9oniE9OgzYvTXq7vO7iJBeyAmFMmn6lbleL
MG2es4WC345Vr1IKwUbcRLCdOudQM2KifSZXbRCl/665BAKWcAL3Ws/3/jedvY+bQB4wqePOtiJp
OU8Hjm0OWtf7homEp4Pba8u66whAt0OdZ5B19NmzJqvouNflzvnePrvAx16NnrG73s4L4OsCAcv8
vjBIOkTytLltrHes64sMybSblOHO3DViLtOCFoONHAY1mHAQmqTczR0V3qHymVYY3m4t9VLMM6u9
/KYM3UAyP2WHR2Va/YGqo+j9AIB3MfABzh4sPovMtbg6y43at+QRoMMTXqHjAcWy+/3JQe+snwA1
SOuS4+YcTOTSdzy4BNqkbyYj7dBIW+zUtdrfQbyvpqXsp7m2toYU/o77cDCkq+MkyeTMZ1URn9gT
2gC1STnv1Hkr9CkDFMMu0jqXeOpfwPnTl9bNcVsX4NtQy8U9gYyJ5Gqj8Sr2nMlQwWnfN5pYHigv
BSzuLzoQGbO8Z879K6VI55M0PYH3cZ1KADCAo3Ir51D6Jb/bi+PdsgZILY3UjfLG3coKnFo4vJyO
9rcKlG5faKAgl3pJRQuDoEnj7vldvVHt7coSXKJD6puzuXdRQLj21qW3JVCBPe4Z+hyglmYXaIf3
2VWOD9FBP7tP75JM2pg+ru5INTRXKSIAFbvXTV7/S1Y3xfGFlqreFI9HsVrzAXbqVQX7ndsyXN+w
FUr1cBUrJAlXVw7lXHlLKcYjUBQQjZmldPhfPB3atSMM40ly/SPzyN3QvZJrUy4I7Io8/rLchyF5
8js8bLTD99uDD7uDTDAmOqi2DqBz8LnYW2C9PN0Bykzp3DwTGkdxMLs7F05stqzwuHh45w5+/sSw
PGxKYyeEt6sNqVX1CA6diolQMZDrCW+6Or2N21xsb9RayiebPnMF4UurnAEpqGQY5kw0aoJXbVcf
R/WV9JGV3zXu0ZcCVJ64WImBn3cuzzZB3QPQdDnlVbM4HbRI8uwi3GxIngS0unl2YFnDxa12SnmF
efbrHuT1Nlh3LdDsvcjVUQIZGgrydHvWWjXzqT68qsMKhJvzKxOoJ4Xb0wGtJkLOVzbpgfcXWZq/
MkFnltmznOO6vgoM2/vayMv4XmyL0JjGVOm8a84k/yc3W25d1w5L9hSuoxlGL0M/j6k98qrlOtpC
tOOzLO7F1VvM/7jpB5otLUEbSv5Vo33Wl9McuFatAtcfYJTO0L91KqO6EAeFajIFqN0AMB1bNX9d
gFb8+gNpGL+hU5yAaVicgEAxozLx59s8/DWhaK9djaq9RrCnkCprhaAB3YEDL1UbBiiGPf4gJ3Xg
TBdzMVldZptdssDMdLtNhMoDS2GmhNJK6Sm8S0nyH13+Skqv4FxAF3nAY5TFTX2Ckahry9jHznrg
LjNqK3M6K+Rar6eZANbx8M18yqoVR3Ay9ocjR0RxxVozEUMXuo/P/df0eFlgSqGYuUaAD7Afg2Jr
rEeRkcLNcuBOooSlvc+ly2aNonIZJuy/CJdX4hTI26phS9PJKzKYHW/brAv9S38Q/2fKVyrru4og
xGzj4OKH4P+kdvCkV34DHtQZ6gw5sVhemrqjL/k+4Lswp7bCiMiTfDwtke38lD07+RCh7sOxogDK
aOl9JPwFcbdqfu3AXioCtPhAtahWg/gffv/g+Y0u8eVWgZFvFm0jw/8i3zknR5hiSbsNPXtaWkLo
GxWSCvjsUWgkmoSP0KiXXqJ8MOPZogtDi7cUAyfMv6O4WkBp7klq1cC1P5i+F+MhIEBWc1VstHNm
4jjNR2mhRSKi6B0wDgbHqzNHbPKwuNeONg0ea4IYNWPZBf2BTy9knqwQz0/zVi/JBvKr4sOfBExd
xBxhoFjvgSVVWPkMFVQjuSsnaHGEFel4sJp9pQgnNMneIwimCboubOfDhCFIC9PXpUBAJfgy4yzF
Qtak5LMhM+FZmR71N1QJBt+MYDHuqESLs/Qp+7HD0FZt5ybUTP3Go1aHEuf6CLQtw2FfmXMaLeZA
egdM+mOIno3q9WuESmZsIf6yeZV68e8XEeS6ojxI1MjREhudItp3LiQw56cp8vhqUJqxqgSS9Aih
V2Yi32q1Yulhl/WMkjb1uADszqSxREZfH+5uM9SnuuyFkmsFImA2DsJNSNxL/G0+jEIuunc0FgMY
tngz+0iyAqoepDbct60De4hOT9G/2NdN0RWI0GCzTtbk6WgElsvbw+q1MiXiACnmspUYYSiI2rZB
Rxx0NN83fmrLb7E1FMQ0V8Euif2FXUqLi6PFwUFKKfjnLwzNh2TSq0aVlsDDHazDY/UmULj9doGN
UvOkEKrLlw91yh1m17B7n53z/LvwP05LATRrG12KR8KcQzv2cwB3YWYCYl4zsEo++xd7Qxh+TjLM
s/DAQyl6F+RE7gJ7md0XcuiX9R6hA5dCSBs+k8VR3itQCy2awGJzKUwRp0CT6kcK1+mAQMaKm1vk
jGgVWRN+T7abeWCSkmkF7YHbNDvz+NeYHR7GhPkXqbwQId8gXrQ6AaCEOz9UxJzT49YOhp0x+X7Z
9aKOTxh6SgXO2phiDKcgQfc9pbFq5Mx4J7SQ10kfjNrLBUc0zztQi+gLtAjj6DDMDKEclimjDK+o
13LnDb6H9yEUpDE7bVeTNiVHqAvxfBz3s6noFrEKjKm7tgGlYJsNFCy7mzG16x8hhS/S2G91c/57
e6yQNkuHUI2NxcFtC9UGgI88jAqzMRbk8hkvR2aSXfH6GqVwVfRNkpjoD3iVGxWRjtgmibS+dws1
gqp/aNJ5CoHXH6uaQVijF4cwxra2Xj8kXAwlr3DPNB1DaLCHG/Eucmy6w/xKR7t4vNatYyyDz3uE
PYxf4Fr742tJdz2uHeKa8wINw0deQXi8DfjofQ8RAsVKs05VphLLhHucQFeyvz9UNR6vkGIy7eao
bsFHPqvhPRehcWu+KWZuJkMLQ7vTMDMYEAP16cggF3LVUpur8iDOHR40XRVVZme0qLNMKKXUDJkt
MD8XJ/5JDR8kF+NxziqdhDN+OQ4gy5SZc1ZblBIMalt9mZJruj6v8gm/hzrVdBTfmEG/kltNXNFH
5tnQ39HyOXrDJ2aLCaSBNGMK7x+Sozc3ombnvJAKbmMOY4peq1NBp3BYjeZSfTPmZwnPgYpM4ccl
iQ24O+0Lc8rTFsK5LAL/irlvJizHD+miBc4RHmI0MZSJp16n4zgNqpb39SiwcvgVrgB4xNfpC14e
IkMU8Mzegag4GSyigfkor8fbbqOiFsREKWfhyRPpxEwE1ZIu0sYOZOf0sbb1yqmPccXKMcdrS188
MwNjiYCszO8HHrv6KBx/YPHJmEDIYxPt1pAXAb3Q9XXfdJ4wDenwxa74Y7u1gGrhx5dBjNtGs9Em
aioKIFlceFQ4gERUqqJaqx32LOBkH2cKV2VBtegJUyXQygpxXQeHAEo9yKoxIPiz9qy6xyzHsh2y
SSzhL3KTb/N9mjJSd48snuuY1YsuN4GiAuURR7ubZMOHXGDIpVYz7m6vUT0ufnWhsopHUIqLpxFw
alNv5Cly+gPSxFeD+oaYNlWtCd+Qe42yUBabU0vAbRB5r0D3PluON8gI7cO9QCu0LAJyW5Do6fKl
Hi33UIssgLL+YgRTQLn2u3IBPre8lZQ6L8GprJ6dZkugsfAv7BIiy3QVzvVCSbX6igMZM6PNSDhP
IPnJHwh3+WXu/3EQ4CrxB702da/JRlrAuYVnCnZPSImr5jVVz5dChGpBmQZBf5vUEzfjuYTK8RWb
X3yZpHxk01bQh2rRlrqiCWTBlKkBNGuUgL0Gy9/KVQ4kMCfO4DFBS3lPO1DTz8JNIosmvOfzTLAL
oWHnCca2SoeOnvuqG9Y027OsgsEkZQdugx5uyzKKyhYjXiINpzcn96eFJvgr7E66KTjPCeeJj3XU
KBuU7mqVfFEF2F2S6Qht0OsJnAL+Ui9LLzCT2oNoMeu+c4jk7oI0un+wA4l1/NVmcZAxb/KEgER4
YRrCDP4/cUo2DNWecd2VUm8BKX9oCs+p6XWiks1yv4Tr9w4c2HXibbMcQMgx8Er75YcH0uu13iUU
8Noe3NoztgNTCrUOrC6ZBQ0hYpQPZpYDtxIqZBNEyzVFwse9riBNm5KeRzUecOViePC3jk8b1n3T
FI5Qmv0hL/9fiIK1CMbVsQzIZhu/VJghsFsgdsoXygx1cWBmq1cnX12+s6QBHOiZmu4z2q+ZyPMJ
Ae7B1LJ/C0PGz5nVHSjJA5++kSW+eeLtdRcpxKcxsDgqojcKx7tV5cIG7FKjW68QgnSHYCOn36jn
ciWtXacrkslnUop+wyVaA8e8FEsv9GlyMDBwIBUog3DVzY6CeiJmTVGWcuHHsVn9kzvPbswC+JjY
X19qjG8D9gHcwphXI/08gGSo+l+Pd21HwgPXyCl9bPD9BzE8Pun0mON9CalMomMLsEZxeVggRHx5
toyC26VUHKR/S+HwlBFVHvVTXDMIhpWrPcDt2EmO4Tak+OkiCYKkrnsUjf215/Z8qlENE2C4jJGv
AWF/3CHLulQrwomTQSqHTQhmLrmEdhWNzr1+its/k+lCmV+s1OwwBZEKrz+r0Q2y65E/XQT1RzoS
1WAQ/nshADt3rkwetD2pjHExigwuiGSMP99O/RWzgMWM3x/G7JpZW50LCa0ru8ySmX712lpN1Edz
pv/BJ+dsGarnxRg5WYrWPIaRNM0pQaE8F+76SjpQTBq4PR8g2pdvVzIrFsnqG/Be0yl9qwiWuyqH
Xr0p7bD92wB2l7dYxdUQXw9oKhdEqIVpPY5J8TYJFT/RlLUq69uquShtlz9Vo+XcUGQvtw6tvv/A
vfE9F0uV8Tx4xZC+NQF+FsXJx/Lq2nFajuYJ6EjyrnMuhfe81nEQkGmEw26TSxYBPvMQGGkgeJsC
XwF/CZgeoQVwFyMF4qKl36I7pagUhOioQo7I8pqP0jyIvdiH/nTkOz5A/mAnsOm9ZM2B2tGP5a9s
l5DIUipxg6jkQiNFLrCQVW49ulIhl7tmlqvFE/yEvK2em7hsZJd+duoYo1lUMTJsuy4UD4wSKq9m
YyqRzM/2lrgh/WNZ3Ja6N9h+GiYuXYLHS01p9EZbsgpzWHNe9jYaK2v/wsehphBSD33x348hwwJa
yXydNPrU3j7j84d8orIt/r03DY41kPKKq/vjG4EL6nClsMZKd3jP2B1wQf7fUeSfziNw7FBiFzFF
cyGSpOlBUC3ZMqPqCRQ1aMU9YoI3mObKX6v8wWN4o3C7hZ1fEbDGI6GiMB8jjXxsqsUK08jt0sTU
ga/xLpjHqCJ6FH6i+6m7Z5QJ8g6U53ybSZ8nNlUyMfnwe0wUTH4sqL/7HcRhzG3OGovNi95MYV/k
QwqYh9+OUjSSYPh/RP0WqHE/7WYScl+bEVJ6qJQXsj1JfNQjUJvv93Q92xMoKS0aqNHBYHIg1zvt
7/8D9dWrUjFSTOja+mrbM/fHe8oUBbnvayRIP2J9bwyRBFz1ikfN6DL4UwjPoNfrYUXVw0zdKkgV
8Ih3o3mIvpMDNnlDw7+68r1UWAFZcOjknMAtyCk3MG3jJpFTj6lU1lLzFM8u0mJw7xoSGTBTR+nA
p9hw1hMUecNHwmW2LkJkfheic6JPZ1zFNTxTpi9YR1iPYn5wrotLSxKO8UxzMrMdCIl6ICZ/nmi5
4VeyTtAO1HO5dr8x7hwF7kNlaOhnozkaS/uzIbyEv+OyjIE6V49IviBS4c81mVhnSlcE5vEGEElh
slWGZ904DSWoOdOT3osBTHlKTODNo5Q/a0ZaMcVs8SenfWAhEIfdvx8kRnFvgFzWKF3ETeKXjrjE
XvYmPgUPrcbO5MdE0149IGGX9SyeFcPs1NHw0bMEgWA3zDmNtim9nEgbUwzYKfRsKnkKvZeyAVde
J68vFFpdVHcB3uxDSj3mo6d48JH+kxCoBLqBBmlwsYH43CDmqswdGgPLT4PIuiGiz6KVDqQ6vQUl
wodKZ3Ti3E7u0k8b2u+jYzhgE+x9XQs36+3ERFiFvq+lZSn3BUbE0vqKqnqrWRLD6Ccr58CK5t6P
6vHLR/Vxq6jdCMQOEwsatW8NRJmggIIy1AFrCLTsUdtQm88z26GE5Ajj2A07uZKvFbZISz8g9OvF
YI7vk8Xi37c55ffDZr/gFBP3n86CGpLT9HwmOq/dwGwAmC2nHuOHMmcpb2r1skfoBhj+nLqUK9W/
SfZa+mhnZT9Yki2vmTEp5Ai3HV0pyjvCoJEEgXvGQtPe/upHZFgrr9YJmOI39i0g6hV265IhRRBZ
xA0FLrbrdYomqFc+8VNOPYi0Kxe5bwoDUwz0vWcPbkmWqBYEOLiE1gFT6d1FZR3NV0zqZTIEbUIe
S8trTVb3uQjBXyQ5ByBadR+PF/gu1F9HNYDcz1zZ0TOMcVg3b8h0EPfjx6/YxKqeuUP0CD8CJss/
J8rWnfJcDpogw4KVb/4i+UP8QHSgG3vgkFKjMd3qlJr+4mE/sLuQH+V2mUfeQev6dxwGkxGF8PR0
jfRBaCqKii50lyUowrigQqz6O5M1k/tAw5YjiEISRiBDriSjhX3Z3lwKOD8nBYhl8kxKaGKrbUgo
1vzr1V4+yVMpAE6K9O9N10aHiwjYlZBF0q6RmKoz6qSJ+ZMjI7Bd1Hte9QaRqmpyImNouQOZ0Svb
TgYxYfT9OLzXady414pDiYslFw7zqDNQj3XA22pPTwGe9vWpj+X6eT3BCH+bPCcC1oG7O2dDkLOW
FnmGNcNrg2FGf9G8SyqBRdYnNmxQ3UMmJ8sIgzsgi+NxwNzxPLmhzbM9GGQ24yIzLrLK8766Gh5H
zSpXGM0Lsk7HOi4/es9yqu6O0iFddWBVsCTrENTXpLlULGcODohKcIRWcso7skC/I/cIQ+2/9VlM
ux4lz+Deu3yUmq98O/4s5Ab5Y6qfHJJ96s7F/IT6uVkG/tH76JOTnLUqeIaJu2kGMph3/F/vPcAN
ywL1i4TM6Q6t4Uo2jlHlTHFNl28xJig3ZLfbmwYoWCmTxnXJbOS4UxqiNWf5jQObQpUEQWCL5Maw
Bpv/82NFmGjPwoLanWkVG62vSmF4dg5+xuwWvmnyt1wzIun3ep9EGaMGpt7po8ZlMJtr17DDB0Un
drEdOmP1wpO9Ih583MW6Ww3xGcYNw5biCCapjddnwrtGH4KvMz2Aa7VIkNSdYAyRDuArFkLDsfYQ
FFtsYZKxxKUoDC/K2400Szr0lDUdbPyfUEtQNl0uBC1Z0dFpDtUWCzBwsMJiY0kZ4xfLz+Z0aiWO
E8qSS9whrfPV+D2fgkd3I/F4m9Q/CmG91zdkxPQbhx22a9ZwTN4ucHLtqq1YSWPdHmbj8jVsQ68z
qOIbJTjF4bkwocI0UmTppz69Yq4pcvgosBSfKLyIILzlJ9ZqYRRl+KA0LGODjU/3zduuCWPdijvi
v4AmC7Js9fUT0uIfCtOqGeLe8FZDZ7Vn17Cz98UQH8zWn0xf9R6tcwwBK+lFEZL5TutXw+D6vQOZ
2jIgXgWATN/3Fiyk8xiHS4cZx/ATE0fUCZCxbmIomiy1w6Myf71kuipfmTLmELIGkkfubLUu1WPa
6cRDzjNgjRZUQ1XvrJPkYI7AjM5+GjorVOGv1qiqBNH8KEOqdFxrQxgFk3q/z7lkKAK16VbQao4n
j1GciDt3kmIscEyRGjlIXCH36BmeOazyTMTkt2/T+N/D1edIWhTWYv5jcrIeVPkK1N7IlBLEV0Kk
cr+BnhcJuOkg/hsisOhwzE+wTbjMmu57g8pEQ6GIGgd4qw1tC+INN2O+qTXj/BBnvC67Hci3wJkc
CW0sXiQNYdp6lk0zC3czo82kXOgvMHl9Sw2h5OuTAxJzeEVdJjD4ufz/Eb3KtPxKlqeIijP9m41S
Oq8KTj6bxhphZAW3VYnuidopJEkWt6mNB0QUdJ+QXWXbs31g4BIUF6wUQHtdh4niRfqty5LctWWQ
Ts3DL98anNzO5ef5UBNRA01MC34SKLDFEOwmGQ72JpOov1AqYM+PBfEznsBMvbM76cn5o41XTu2W
VdSPNugj5bJH5n58+0qv7krVxuIKhomA8mbqV9wYhnPsqxv0g2Yj+ICphbjF3rPCU4QJaAmG59i+
FefZttqQcb8sv2ROvFVGUfc2i1YwHibVHZSx4BEq66uS+PzbHAvc+yX2J2pNsma4eoaKIrODLfhi
//YLGf+UX6lNGVOrrSI4rv5TyMSnAjHqB/BMq3YDaSP/POdxa2Bsa+nH+G5MG4N9G71E+NVPUG/F
+KqLrWcvgNFNRpDo8zfIMiSDiOgzJ/mvt6vd5Jyrga/G3u+0rFcPYZvI/GiorijfZ3w+Gxm/H+9O
Ivmu6kT0MNAX7SPtY91YCwX1AF4Qs71wWwXV62/KOVOGpIE8PTqetGoKRwNmGySvQuSLxyIqquK1
uNmfRlzMv+y9SUYumGR7/pmEE58lmbLGi2NXX1YqqCmQepk3moY4o5s7i9TmYN2O3bp4SqoyftrE
vYu0Ws6PFx6kwBzEboJkvclAxw+6sh0s9PMiY/PhsJfhexco4I/GZjNsEoC1Ls57ycxhDqKGkjr2
13Lg9VqpJ9gka2B3sqxRWU88DNr1DVZsG16iolGMlGrncHfCQT5s4kSkCyq+s1nKyPjzAX4xtTEn
hxu4JHTJS90QVNiGaEpakpGRAFolLiOjk0b5/qDSzS7sJgOTlKgo+elbZXHW9PUB8qkJDFtOT0Fi
dYTXvsygI4PLE9yFgmV1t4147dNnHu+JJ8ZbwG/oC5m5oQx/QPr4SBHKBGF/8ef6cYCsVm08jNvi
UDVdBJte3bw68fpmQUrlc5q5+IPLCaIo4Eq5i2qcxL6Bx+25cFZw7VAaqWtsSDHgm6FCWjrgV8bR
pYDb0nLATJsKU3oKx3GkZr1jvy3f70mXFJez/USl4+imIS6gSizj9tvAq6EMc6jlheq8hv4R+JzO
5oIvmSCmLhzyg+1RI0iI1MHV78bPEDZtorWJw4gh8BulHguCboqnK7OaLX+TRf5pClyvQ2gY2sKa
ZTtsWRYr6atmcfFQswZE961ERzxLOWL9VV17hza+VI+OHgHw7ZMNg/NSdsIwqYhrPEJjEImgUXXp
/+DCbAQ4i2CL4qaR+6crkws+N+BFn2TW32Othu6CjChYX/vcrPNAzbZXS9VGzUsNkycXnovhI7iC
gBMhBoNcmK3z/P9UF7FMNnWMoNtno4iLzey6mEKL0u4EsQzWubiPwfdQLaoFIGXnAJMZf0IbTEeu
m7RWTsyoUTSA+ZjrR/ml6oB7Nymy3SdRa6MrXwaJHQyGSAHXAfBGVeqmZ+QiRoLMBaRDIqRqR1+F
4ksZk/HhxK7NjrPU7bZuMmt0dhpXRnUQiRLSOV1o6GpTm3/k4EHyQVnhXDtIyz3Pj6pbyPxsR1/B
TFyPjkSm7TbujEitPxMgop6trK7ny6oikqUZm8Yq/zmTvgd/SNx0Gp6itMmnbS92jOpbw/CaA18+
guEbMKf5+4dpILPFd9vtWLFabKdGFwT6hVR0NjZWEbpaJeiV8etrMC4Mjei8kjtIQd1HjJoxYnhO
JM2X7KvBPCVYzAhrQEy2fKu6yMYBQyj28ZHhqyoWAzbot9vj4RKmT81oHsocz1yGQvhqAqFv9i+d
6PQN+dbYmQR6b+rGlGkmTm3HocwmvY4aO8z2WQ1VyCMWLG4isZXhF8kQ+wPvj04OtMOuD328vzD6
LW5w+xNdtrdDGEFKpPulRfQdcQj9eBqlBJRDw0KGWixt4gdrq5PK1sy1F+J9C5vop9ARYLYK45Y8
fOi0TjGCfGEG5NSTmkgDlWDZSbRPsoPMGtR1wofSaLk43YHvN239v2oD3jdDNU4TIa62rA4zWTJ+
FRcYVYQb8J8pUBnMpz3U9zVoBocNzp82g0wcgvt/4MfmLIQMb47eoOF9gX3pspIFfYFiiBFFbkdR
Yl7M/z+4bKhX1DdHCi9Q6ct5aH2UmiqXBSB8m694NxxQMDC0PgRTeWot4BHVMt1fCvgmyM9k3XBq
tWCkdJnucnWltn5M+kLUsEJcexEAPUQ30KSWY3YqzZnM3CYK1t1g5gwTxR+xFDGYLuoqPDihsdzC
pN9gMCrPe3MJWRlgCjo7O5UACY4bSxwvl9aOoXq6Wk6wBVe3hjVK5jXTSy6JjriBHnWCLE0bxmLr
NyJqb7j6MEzd5OrmQmCbIpyfEvjp1dWRd2tcPm59iRgN2fGkNW0wzuU8s71e/8L01eqSYC8SqY7p
+utsOhMoIqbjPl2SkRETN3/E6wE15lUCGE8TD0OEkH2hM7dqZiv1WcjCE+bskS+e42QNH8ZouWvs
FoqpB8RRG+pS1uYQwwsmmQa6YM1+io6jFOq+VdBSxLRDM77IfosYvwtA2T/hQkITHni2PDFQHLAw
Lfa0y4KGZHYs2bttWbNtEw95LpeEGaNq8MRR3hOy1U6Anm0B4/LYcP5aEA2ym/p55+bI5FX5rrHh
2ETf+f7b+CCVMggB5AwiKE4wmrHZZt4ZC+Q0B324BPZuKJjOaHlEdq76SGUb6VSXK8lXdC+fA83Q
CvR54Jrrflp1iVZfxRTZBPdFbJ+UK4jjDUm5+wbFk1N+0ROWmVVtTyYR/j8mGtD9GnprIhBi52Hq
kEB8MsXgBGdKI27d+XClPTei3VkdhfOs1QyeLhD/mx21NsACNGKpnSI9obbBlREjJyKVJhdhZmBb
8UY00bXT9BiL4zHRKUwo89k7/3j+AbqyJWuhVWQtqextvX5P4H7rJRVEd9zzZ6Rn2rKuXMpBcy3I
bzdAFSbfJFYjsS7NBnnovrJDDqdY0ty0FBgn2k+E0gSBCNrxW5gEUH2I6KMT+Pet1A0hvy9+7fDR
fgfhtMzxZtI3twqNgVCdwMXT+MY3F/1r8ptK3CO93tUAVg6cY940MhdPgGCLG49kBAMWb3VgGUx0
3ASWUh5MWONykXHZPya+n2vX+ascuCo6yZwymaZBZbLUaIXJrHHSAdGiS2qD3fpBJweNuFZFvMEe
wYkK0P6YFkuQsXTQXJ70WsQfFJeupYuhIV5ukDoHjYjv1380PDTZmqEOVBB3rb4zhNMN9GSYpMoS
7ver4tH4i1MuaxQ0Z6fopzNJ1LLvVxrSO3KRsHhXWRDzrc7dvcj6tGqblJuexxwAmY5B9FLKy2cr
SKv3QCltO3AWcPWyTSAzEtRR0mjHTxD1Q8z3yOKDA12m9BuqC4VA8nfXhkTDPv2/0137vxjK1wZ5
RKgatlzJUqpCW3jduVikz0fJbQahrixN+eAbhl3qwDrpwGUbSolpAg9opzyEnpl/HF1xt2Cvs3vI
JpluVwuG/pcGL7FSI8y6FeKAADFjJYv3s0y/U7FwBahTp8+uX/Mn7NffATrghhVdsEK5/jZux65T
tgoHKKgJIRnTu9ykEhOo5I3XgiGslk/ouBvqktsU0jwVSijRlXL1DJH8rX952cB1pbNlxSfsTLPP
b8x/hIRIgHaOUtC1hQ/JJ7fAbtJh/qIDbJl6jrOoPbxyebRrNeBPtTVMAjRhytEAZ0SPRR3zqKbH
Jc+rfQgNBtRgGzLEca4aQ7G17JT8SDHw6BHp8bmeF2z35+6XRBcQptmOVsgqjab1+HyMn7RaJVqD
JjeZI0lLqqjvP81cnrgwynmvE5kKzFiGWc2dMz/n1RWdSSIrESVb2z/HIUzbMi9SHejfW6E4ocnX
Gxm1D3oB5/uudg1hybCxOVKOEknFsi1of6z08UkxfN1tvcQnrvZXcSgvEjjuYR3+cmzAdPQWlTWd
AXFlaqDxX2oC/E5MvPJ+m/0nxu1msBb20M0yoppJ+zadC+rmwYeGmuvzx0v2cC/refJ3XcsB0Aov
manIfuig12fWG2K+a2GisEFSKHlR5bnEXAbBwv5Ozuz5E3XyflarLF9xfnQybbKEUWZRjzKygAl3
w4beCQKf8lfMvHaOkMZsAXfeHeCId6DYYjoOzlmfl5sbs5fjpcWsdCjMwjjRo510mrdw2t3Nlf11
wqdZqKFQDDBVXsWtNO6BgDaR4la4Tfp6XdByTxEywRnEi/oqbqWxmUCslVZSMXsRFJForazuT4Nx
RgHcX2OiUUfE5/vWJl/B7iwskcfUwscMEVEJkk1VkWuJUFY3KtnmG0lWKuHsrBm7epbaX5pbCm51
X8KUr7S2So9uAn4nIjnzCg8umLrSSolSteA+JCR/g8oxZqiL4oIKh0r6iKIpNQGO8GIoyv0DdXTm
eiMnEtfZGg5xdFWz2xnC2gHXRBEGneCTFNbYalruOWxBuJbmDKMLrkk7CgygMJXeoyG9zd96H2kD
Ru3Yb5yoVpWtYLw85hrx+OkLnnRXJfp6TSA0lKHiKYeN3NSubrq2QGAHWbyjE88ZaaszepDPSwsp
VqXWG+5zHcXR+bUXmrYZTDYX3bo7oo3qQ890JrZqZnttjMwNWqxmQQoiwwHRRGiNiaQ2YQeQ9pUL
cdR+xxxBV7nvKKkyxmIb7lzZGmJSTpeeSTGKfLMGR65KHxqZq9r3o53g+tobe9rDJx1wGL5XK71Y
5gHN1Y7RvAkGUDd2WxtYrR6p+xKSvejSK6KHB56wnxPSwPH4y1NMuuffIS63hTAh9IN4D05yCQPn
zLp6bD5pcAcsVAwPbEBnW0P+aYwSew8xFaBk3tQHeiXGvOAgJjC7kpOCB0RFXPGzozoJ0Hjs9npc
VKKMAXzfYMDLElxpNr/TUf96V/rE2UC1JISFELsvI/xay1Drc3ZACgv/KqPb2khBrEt6JRwBs1Uw
kZheFZj2Mh3VvQ715dNItbuQTuH1nwxP+45Jd+HiPEhzlAym/eaBNaBwVoTznbfGE5kLY2PelUPK
Ql/rkOFZcl7k90kBwXLMUGzMXbNlzdxMB+JedIRFNoO+lfXVqcAkNEPsJ+JzE55kwmJbPVMtI2Xe
/nZSVYb+y/3sRqLMKals6rOl2FJfjPLVnn3YUebkpCBM8UKixQfq0GKQhs2rPlWzWKkOijbddDH8
SgBxXur1WgvPdkxBTNzjeg7+8QTb/RR7juXjG+Fb8D2KptMAO6nvxWKDhtsjthaUpL8g1QD5abms
SbuN+qzKIGwJL/QPjT+mAiQCq6Ei2t2HCpG7UvWJCCWJ6VHan2gCGxBivKaOPYkx8iR6wwCd/2Sb
xL5yTZZZA6h2quR8YBIaeUtRWhCqu5Fv1/uK8rW17RqZTJ0wMGx7s0udDdmfW2chxC/P7XqxLjX5
FwFM/SJA/mRItfy0x1ML3ZBbz4/mLS4U2ccqZJry0y18xqRdBhxDsw5D3a4EumVLcoijUZI9iQhU
GBok3b71vdZ/wlCUHaKKJ2+u1pkzWcHGzdCI6dnruJLjfp1P3f1TYeabIW4+6Xn1eQTedpOu431u
T8jYVPGLQ+fGwV+NeEKUXrHBNbNVgXpGcnSSrY/MfE2FuZJUvWBsgx+iUe7xSJuHBfn8MxGCAkhF
ncu8+re/famgMyNGT7J5mi1csezex5q5v0f5H6y1FTg19VxamqaNW4frL8j6A0SUqRUMOWN8GK9L
5XC85bJSPN8wDOLtU9ByCZtbaB81tvwySLtjNwZxh1Jx5wCvl1bQii7jm3TZV6WWFdIThZ7wInx+
gcvC3Xub69lJyFW6GmUzFiIkMVaNSBpwslq6gSbPm/8nE8h+2z9GwkGlWShancvSdyf/dmyCgZy6
tfGUahFeOE47rSk9fpaDhhc5GcRf06D09Y/5Jqwa4ZFzr6ikQ4c83+8X/SbaRPCUCnMpXx0BYq9P
HaDILQPqGKJt4ROC12FyBw8y03z5muzRDcRWvqgC6veo8L24Yh5qlwugDUfMtc0JhqOGXLtJ+440
v9VwGelHbnk3v1mvE4Q/mK2wazV0QNb/96CFTaXdhFgCDSChTdDmoLpHP/xL225ml5ysckjubM9s
I5uMvcYXa5kckZA92nUygKeDlbTu/KQaQeWQXfth0ab1feS9NqZk/VDvziOplCLy/ULeGMymTMBk
o4wTRkIAb05g4sfIjeQTzbvuu64qtLWfn+iYpm7x6D/nz/+qLHmiT+I9f2G9qTavIlsNPkUvFUqI
RLuKtJDbojCt9JwLuoOt743Sp2/skxEk4v3xsNrWLwKQrW9ajcEDfpbVOqYtbCy/3eXmWYONZeMT
ojlxHMRNOvjV+4Kzfn3tSPtwPOsSeJvLNIKhQIDyLzpQwCa2cce27Ptk92U8C9VwL+MHHiC2GDTE
SNL324kaNv6DpRlfmk+TFpEa320shB+paVvgFddaNeltpzraul218y/oq2dE04VOPEAmaZBrVoMQ
gboMHQLMldVExow4vYtCK/eOl0OqTaaw0ZhJZyQ7bE6UzomJAExldxhAQpjLOmKATEFx19XPEJ2d
aV4Wpscr+w6L+IBSH1UNlqQcyECF+HxAQWLcGU4+3ihUNfjNPWT4M57ewu5NNXPG/XRnqqIqdqfJ
9xWA1wGY2D7vUqYmwY+3UANj3h1yvjvqH5GVgLs712iGcFm8Ss6gXHlg0kPZBgsaT0Pz05KQR+uY
uj8+NCqmLRALw5nOnPQ1Z366NvZbiHVvqwph02XC97h7Z4FNUm7QTKcpmL0V1u33f6v5gAOx3EQZ
dxyoVh2BLCLDqqOIKvDNx9bg0EAUg5arcxgxzRYjFT2HkoFagxz8USjXXeWIYb5IG5nIY7fnxap1
HyjHfWTeJe/dGLYb+1QaATYQRfkpfR1bIQeXtMC77+YeJII6nHyCGGrE8HBHgIkySW1m0ARVP8s6
M0Vv1vAj39W2mip5eHpUi6M3f9Scm4wQ35oaQp29IuhUTElE3+9qrpMb6yFlQu6qx6XeoZfcxCU7
J0D2vVp2fMUfgzqUfQvgY4iG9SgLUDPhhaMquLSP6rc/fkCdQ3DYVyAFgTzmiJWCsD46uiCGGFWo
yRhx9N/cTJXZPVdijvFkrmPkpbkH9LLJhnZad61mN/IdBrowka8GSg1DUYEykE3rcBXfOKymQcV0
sgKx3q2hWbtJaGYu1m9/0OLBsnI+Y7Xj20ZYqmEQlSd7eZ6HYSVhP0FxA9E52SZ6xfOEv7ZOSWP2
V+koB5PW4lCCiG3R8DHNHn+wER+3gGue03comoxB50aY1M6jTrrfXSpv8Jam8AZUHLi9eHL5rz6R
9w5E3UCPs2U5XpaU0Ds08fN2oKEPVFglWkaMKZ8khukaOCJs6yDBZdj/6JiVmN6Cq5b8foPiqmsG
Nl89pqBB6lWav0L+EiKwYrrBI2+9QyOAqZG3lJx4OsDv2O8in8QSaggZR4RTvR6f1YI5lFf/k+LD
b0gNYn3B8yvM4+ZqugY69SoC6Ej8VffYDbvkRMubEAghzEGRxyk6aw1y9mVFVP7YA9m8z0XPZAsP
eK06D9SX2+IMioa+9kynKIoOP+ns67h5Zw883sMdv3hVGqCaWGtCqTjJh0l88S6FnsvpC1q2LjkY
+pAc0bqkLjIouUjo28Y0p0I/McVMUZ57W3fS69VFSEPa9Qfn1OSHlvV88BMfaf7oNn928kiXXFe5
vJX15IrYMdBDdRIxWSA0El12Ic1Lxn1NH5wyufqeve5Ig75jnK1BecrSEVR7XBCmyAJ+VHo4a/Kt
9MoI/l/yIKSHR4ovmJE0OZ96yWOo9ayOkfjDB7LQpi45OADU06bn4wkBNNJhyzpdgrI5IBnFSyq/
3IeqWCp5loc2KE4gDVIx0Z/UPDIC3RqWUUdt1xMm+QraKhMiIDWO2nnKpar71y0pU2mcadT+LimK
G2Y7TIUpL7OLursv4LAzk0G3wc6vRoQQvkRB5BM/uMru9YtYX2+yDA/64gPxgwHKz7wlxF1xORY4
IgNRDAM6yGm9HCKjEDCMPWmUiWNLXo1fsZMK2CXjKYUwFcjRqzRPXAJWQQ/+sRzio2GN158Tez7H
54N4SeMyCKt/l7cinWOWj11UoQFE1eVFaKnaZwZ1GH2TZbPK2AvIQiiOA2KL4J4tWD9ujR47KiyX
nKPl28zwa4OrhZJe2pEBqdI7ehUuPth42RoPyY6QNm3Fcm6znGDzuQy+lSVSCgGr9UHFkijKcGdY
FjN/4puUCdF0+PBJs0HQcKQ0Xg9M1RuFh7Zp6tYhJ9NaMRaMiY8IH9lFCXptc7UWW8pGtdyRtn8A
MBkAgFeDpTuRXwTNT7RKoC4rzhwW5pFo+XEx3JqLRjkbMbhfWEH1H8nBOz1QOQazJ+Wo7T+0KqD3
VWuIo8FLfe5tVrr/pbtL3ftlwOQviyVY57bfWVufwbyYHevAprSFnicp83sU2Uiv92MJhk+RSsfQ
KjorPPYZCHPEbQI9COXPWaKc5AlYDd7JXjrDF1KcXP2Y08ana5knSO5iygphf6nyypNTqu1VYMo7
bBGHMCrIky5tayLCfnpiNY9eRHve58UzuaCoZ9uMvuT+5ZvF6+qXaY+FavEU6ZKEbQCC2KkZeAHM
a5S1nzs7nrxWKpKtWNOHJQU5H3lXf31jRc6fK7k6guJgED8hBZUUPQ7uR/5Z/1zF2tJPjto89CX9
npsMoypsEyUHv6y2zxCRO/YfM0kb5MqLcG938dQcUM+YwIqqiqF8ei1XZul8fNJ8SQcomQrQTdHf
/xPM7FvQGvrWjs+ml1yBDt02BB4zqLj9FD4wJ/Bu5yLKu4RSxcYCMnQJh9C3mXRBTMsCKEDSjTOl
Ez0WfHqirrr9HkUt5XZNrGwpucTN7h3+VwnlKGW0TAzrnNyU+HzoRrwgDqPTpmyNs0YZNSzO97eR
GgrrjsT123nj/ylKLZa2SmfXzxgnR33DrqKjBvicyNdf4ubfFaLYP200hO8ShGF2nCRrlJGAvbEy
qku1WgFwah23SisSqweJWZh4umlByY3gVc7+mj3KHb81JRT4FeYmwxPgNLKs+yNuvPVEflC/lLHi
GuEbRdDKZGS8kaJCUUJMzjPQzBjpzusDx1fdGmVe+t6uL4v+Fwy/Z656ZazTVVjjXa3thYMni8Zo
dVmQoVN0KEA2gAzXqpjbr4aI5m9qveLr9IwOwEg1bNgRXXHh5n59Ze9DB49uclXMvbkAPpX7+qz7
OkLtT2DosbtfTl8IE7AMU71DXREQyhhnxjtQL9Ytzvl4/ulR3+N14RV8VvlIqehtf6ZdfMqfAVMN
n7+vovOnn0QYXYreJi7PiuIxQJOvw3GtrAIN1J0OkF+/qjuFHqri3C+R5dw5IH7A6QpkQ2mkxY7o
5lPhigYEKrxctIrHXf062Pwm2eeRIFcKxNyFy0VJcTbtZqlUxiEdqPJBI3Uz0OYrExg6oI5MbAU7
ougO5cq1KNYdq8lbQRr/k0G0bDG46kGyetvbk/ZUHpBltDtnrFBW2HRS37YuGQJ9oIsTSju94Fh0
qDcm2CuDDcTUuPy4Z/fgHycI44W5wYI8b23eV5ZkFv4qwJHRDjbFhXFMEo2pAuz3XpSQGtjLt6x9
76ydvyN/oIUVjINPqcGnywF+/ShctRCHg8t6xwpSIQitXfPaOi+0WE1KVCgHF6yyCFIqYP9/D5J4
fTNYZt1a4psuEowEDZ8sy+wNUvJiUgx21COw4Bhz6UCZGL57xr6ChFXVw6ewE7TmCnyF2tmXDGmo
XXSwWQHOykZWNTA9umB9ffKVUmNw1YRuxYW7JV71oGSOihEeuLWUXFDY0pUFLkE9UIE6tdVosNpf
5IFPNed8j/I8Mrn5tgOfdrS8E9n00Dgwc8xGK2Diu8gJ+eE9pIsy+mGpAmEbNyDSmLKRSlQcupzj
YVvLyTM41F+GosOM9nAcOaFycC4d7Mp9kfaZWXp+PxVf5kG1yrcCy1fY4jLuUNpIrYDAFl35pZPM
/r/bbS3vNjnX4/Kzg7O9nvp1MvxKDaWBI7nqDT53+fotHFaxvbr/j9Fe9Lb/4tcD/IaBf8GF9NBr
u/EH/yCQBR0ocuY48/pRMH2jZKZnJQE+7XxpPTx5YFH5QWg7uCtBD+GumY4y1ueI+g7vWIh1PyYM
KrDNYGz9wBvQa7mS2kX5LmJJMOs7dua+xCg5w1RWqDd1Y/hwaywsM0LA11FIJGK8DQrSv/B4XWpp
1K/uzSMUy1RdmU+vUeaYPa1PwUy95DuP7jL5MqTqG5F7QUydU7WJExhzBggIOlfx9JQ4DYrionZt
HRP3tK4JHhqJ3wzQl1vd3JtQOwF2EZfbsBwn2v5339bnlPwkDVDdiHGSIP7p4KjSyFWDvk2dbqgQ
RtnFVTo21R2+GHm6xXsZtUBVj5mVnvwITWX4JHTWU31E4UTCUeVgP39yafZ52eFqKd2dP0144zOV
Vg3IP79IE4tEcbxlHv7qNb+6BTT7CnwTfwzYs4CrbCstIukicwe4XHuB4eD4zENowT9jHFuMzwgU
+NvrdQX+/Zu5AArRlAK8xz4N27ZON/b4d69ZrvWUh0o3em7l4+LVV4i6LNiMwLjFByilwqr+R6dA
3+4P0XEmXHe6EelFXyEuQCbKPzpowfLv34aBfeg2fU9eNK21awWu7ehQHG7U3tSgPluJDRE6Oghs
3S2/eZtdt/PWpNlNELx1g2U+uxlwgrtGdoh5pN76nQryiEcmV7ujgsK06L2CK8ARnqIl8x4n4uBW
HD5HaQjnrFsIv0ryig2EOEr9MyKWCONfiLfXCiz2XCPywF+O3w0gBTLXz5LUL8qhH1tPTRvJsABI
kOfpubSe67KmiOzyHN7ighYZbVF8pXjlYiseLxsZQbNJpfidpHvG3ja5yjrG69Y5T1yrYRoafMAr
i76V1kpaJYcdo+eUCu/0oyh/M4ZEuTIMS0eGZnF0FtBqN+QGkcIY6OPO6uSPJTzXJ+oKJWur648X
EVARQeGI7+rT2bdPpBbNJ0Iy2Cajm/cpLw/62aS0tWA7D0PF/MAwy7BzovT0hRsT7uMcak3DnQT+
KoowIiq8TMYZ9q7t7BA40B9sLYuPhM050rxuCyHOPXqwFcffqS36riz2Cs/afpRywW8YyfQRRCMw
4bnhb73WxyjKcIvINCqqHi0Oi/7l25RMgaqIMFjIbzXK2C3APzw1mkiq5U2Y8+AxK02FT/bN2GO9
MS1mLB5U42PpfA+fQbYghwxoTMOiwfW3nSWvdeBTn4f+i/o69w2TfhVjj+rLWOdzQF0YyHcqrtxw
F/zhQzd+Kttki4FrC23IAnwl5JyFvKCwUjvFPrEgEXjDLqW9MUQIctsZt/0/eUGWIQk6wpLvJ2MO
cwc7pPrdASWcsCCjQcYDz9KpWEWaro6dZI/KSaFGkaJ3rgu0yoRmcq9qtcJGclvDQ6PYYqyjILr/
uJ4enm5LvAozp4Jsgc4s6x99M32BsMCQeh4z4CX+aFOtrO0iKWSwNbhV8qYjpyDEVdNUWl1rldIt
uE5180K0NLsksj9gYHlEA1nJL+QXOd4qt7/5Rop3VhFtbYzd1X+hXaosWSJWLq5BFypEoZEhsWJ2
f406B4I26Z+9bPQT5Sk+2D3SVatsw4HxAEQ0TQLR61BqDmX1hVsW9RF+4EgQeuMdTw/mpE4KqAG2
INamSqEBNKFPR3Dx2k6hBiiL2CpP1o9KdbVCn6C0jb0FAuGvntmUK7BAQoQHPHQNfqeRDDWkY3bP
bSIOsFhODgHwZeC7PnNmmnTEU3uVClzfqNxOLwSmjKiBJ8UXlNBhFXOvUc3VGnB1oZKS2YaCZOwp
NSlCVAlKLShTeQoh+0hD/wkwI630aa/6In31T71mfJbYpngsj+y4h7QDeiseQfoQ/OqzIbMPJ1Vd
5SxHeGgAEYrxIixw6UbxfrSgUln2P3SZ2Js1lS9LSuDQ/kAELR3Ejig8cQXxdCjAaLUcHuB8T4/0
g3z/Pt0O8c87X4jp8TFh8p2TqvJUxjwOTeqbssJ10eAMaxjbiJZ7kD5M0ihRO5IbaCGfR6g9ILRv
05sOwEr1Sx+hY2qCtTwV2IsopUkC3LVGQfMiB71nnOn+b/Ot1geob2Qh9T4Ip61ZJuHMabCIJ9pf
l5hIXoUM3g7IobTCOcrpdFqapj3fKerNdAaLRJOLSehkzNWVyLzWlm73eiGgY2z5lCQ1I8a0y7Bx
j7LFS7VRd83YuWKOZ/sp+iE2+XruIKvspy9PAUdO/mZFMrbla+f4WCE7MLpo/BZWlyCpaGbrl59C
9zPz4pljOSDbIzkFmXvHv+4xHLri36LWi5yiVmnXQS4JBnvXLzvKZK0+X3mftzJnkYFScKLgZmEp
TuN0vXCb4r04NurdfYJz206XANh2h/E9BUas3hdb8Ssx7o4arHbqaRmOv2KM2eC7eFAyBsnpuZhF
7KcYBMrdIdI1g8yS4GOUSaxE2L2yxIUe1J1kpM3uMJRcuFr8FQwWpCgG2wur6vw50HIlCEXLoGzn
VhXB4ukdyCaPB6VP7J5B/6/6YVWQ28H0P2RwfRFke3pXKOG12BbglCfi3/hkKC7lYAzmX7OQdXE1
/T7lVrpdJLJNEhEA7LZGBeo1LxrhiDNuVxmzRnOJEtuhm3fAugueS9zzDY5wHHZy75LdH++//ome
ScDdpuqJ9kwv2VcJB0CWNHPkthsyrCEFhA06LJIsHYuPvitLtbboyVRDvi+S1pcAEZiZ1707ny0q
e7jAhnPWbDPUPeAOs/y//srtyhSkjjUbjjaqQWhTv7yblzqGJFpkRJ3ovBO5Asu9teRTSlHqBhY5
dhDnlp6l9xJKQv2ow5p8gmEUwsTg2YtuW1c2rI8322Ly86vcII3wBdtUzcF9sLLBI5KlcqGZIBFh
lOx6uSHseYlvX/Fqpm9hcuA46q3tuErcxD5iWqukIRuX9h2Bj8b4Ysb/h8/pKbRq5hL0jEUZrvT+
gfZkrMV8TP5R0YTi+oqNukfrcWgPr2e/h3abmQAd4UxJFlilgbyyIYNLd1l83HqRbGQHj8yJ1pnT
9Cr8gchOcgaJPK2FuDH/EW184xOJc1r5qj1W4ClSUAzYlm9Xch986UDKP5CH1F9MfQAWJYG0PtVf
1yxyve7Wh+9xlB+OV4D/zXeSUP2PDZ6EIluvrs/+4DDR/Y0n+Nfp03MSdsIBsgfTB8RX9Ypy9Ua6
Vg8eyQJ67AWCJHoeGmENTt8zqd6mSFIBg3NX/3PkZiYDnFXUAyx5XKlpZHhq4bzGEL9EEDMfGUm6
yhdPzPfR3+WbSCILOIF1peQfursMSFtD/IWydGk7vBPEUG3EXJOEWcV9OKTS2NSkDTylewI/gmaN
rukTrvcrSGuRUzScZQK2Pwyp/NG5A0/SZuuM4bKhWDBD4qvPFceqlFSAlot4kyh2L6YH40t3RggW
9AFs+brHoBQi2E7D5rXmP2Fau6DE6iV+piXk95m3AmXVKRHOkGR6+Zw7O+JRQOh0CQ+hzls0OgjG
DcE158GkrKgrZAkYWjB+n01BGqsc0/Iy9GctIBYMZcUWOwIRoycFBvDpNKnI0oEpuI/NQjpq8xYa
pkSUDmYJbeHa2zdwupqgzMbpTTiZT0gcaDgoKcAC7ozHE9qmYIJcGLBocho+YjITnwM6UO3hMf5Q
kol4wBytvRv/M1pfMA4qvqh+Cdqo5a5Wgjmj37HaQyX37lXIr/XTkN0RovVPaJD5yyXaysFdv3kL
DL3pb8B/WsAzv4ZHwqjc7aLjyAVAxwtNlzGvG5xxRNG+W9hBDIM3IFJqlDdV3g7zWrkqVBQEiE9A
ewV37roh8oqQwYkTBkLuKYP4uCVX/oNORK6Ck8ZL5P/iszPYKBPJ/9Wpx0nWu1bnel9nh8vmfISB
a3yY7NRg8/bJgxMMPsmuXjPoL26v0tJupIK/e4F/vIhO8k9qwGJlj/1NsWm9A3VCh/g7+YA48tdG
Tfm5MKyQYI4wwsUCX1uXGi0GM/o4/EIGflV015a9PWGXXRywNANrmlF9UEWgssiE+tUBfEx2M3ck
UESeVXal+nqek0AC84Y9NgkVLnAVBgp/d5lgRmo+jXShJNK0jNb3VgyNbShg1zpufK4A1eiueCZM
WiO1cnRK56EFyCbsFZEZO9agoR4CRjLwRAU4Z0qhvyjrmyTSnBh7CswvWVBUgm+eZ1MeXlQy7VoT
HrJ4quB0XUzBhRGQYNPcBIntp/e9LI90kjOWPUAYSv1fzoQoX/MI60tusSzVjGbtFxs7eqe4dc57
KevhAdmaixrxgvgR44LQTEyvAfmAcwI5S99NQ2tijVl/XbtsoWg4p7RLVgvjyI0PxQNnqdPjAFQZ
A5UsxJM2HznE4h1UGG+h+cVfwj+pbbRm+UjWNn8gcjwgFlW8WQZRmC6ZCj8ETri+o4nJJtKigPmk
jL54YejEzKqr3p7e+OfSU+I2YwkT/HPhV1bYMRwAK7UWpr36jNwdxkN1OgH+44ERhBpMI8Gs+iJj
TlCIPnQwRKglOQOUYP/oCvSP5FGw+qxhGSjVtB/oCk/C2k8xSm/HOCP6ZdsUv8E9o5a1YwM4ryA8
LzkmVvIOlvH/Iu0lMdXiG6eSqhjrB1onyo9sGI7crjCUqD5Ozw9JLceWhi9rv10RBGtHvsKZUhvG
3KLzgn5YkJr4ileYDdsBbS0AjbAbAJ4oj8HXtkuJ8oKw1liWTPqioA7nmxelIeO5KizQlS1UogC7
KyzE57G7Ee+u5FFqRZ+c8FkXnsSKd4Xzon4/83KPwd6I9uOq+z+c95UJ+2kdn18UI/tAsPLu/FBm
mcsM6r0RnrHoyApURAes7FKx+eZekBuWAIMp17EPn3pj30ZN0B1r47L/Ct084V+iN/Z21vmlj4EL
KaovV5Uf4suL68IAgQVX/p28KNxZcV1c2nHk1EndXx/ZJmSuRWNn0AQnF2/de1ecvAqfFbeoWXP6
LRWF7maPuqsjRj0eIyrXuc2iLgn7s7OnaLYU0PzDrJxSwX3FKM2z/x34FncpUpqC8vhYeuIcv2BP
YGvwv5mh/CUggQMKUIx22m72EaEaGM0CgRweHAhtV398KwRSJaB1I/4sb/5l3nYO3yQCZgW4ItsT
7IYMVZsaaOgJ4jcfah/LSrPS7a7qBz4leCiKW3MgdxpPdIkUmHt+wglN+9s9YhKw4g4VEZLBePXo
Cjm6ohEydVhx08VbdgBTFsdduOMCF0sl18p8gziZUcA2lEx93DwspA8+EB4oueQ3Kz8UbocwvMxT
qUxq/Sy3vIU5YzloYaxS7Fscua0xcl173PkyCl4efbwfE1ofDMrLDTkJLWze/PqL/30eCW9T2eoN
RFdPP+vGdCDGyKafJlKxMF+HijB9aD8hjv+z47NQrgqYDeYK5lausxpV8IZTfTKhxRDvXRz6c5W4
w+PHdMHFoBTfvfAXoGtWcuXH7PNI59oDzSZwCtWXqVFrkidm5BkEYhVuuNHMZkeTo0aG11To7YxK
COciwjbSTxC+TMscFsSI9HIIVa+M7VHGebr8H4Dcw9uLsueSi0FMoxjdjHzrKXrWMQSx3dhzjLGI
cjmZVVzVZVrJMMOWWChHIEHygwiPhGM6VDfLHyVNa4dH/uop+UlFJgESzcyyvG/1FuLoyuvNSgtW
yxAHJj59vIonETkgApYa8MWxBkNDgzhYe+mRzt50vFczorv3BML52sxakynIND6dkaKQ5VJHBrEM
sryYVjLYVA3M+TuNrQTDXi2KJOr/DPQO+wiJOY0hMecI9LWg9NSS1/Kh5dPBUQFB+8IRQ7a8L3gG
6dbdI/Z8zLaVdPgEAnj7eDrg+LMPWmPqMW2+7BF2Yf/ghh2wNcVK0kzTuhFqE2z4Aps3PiOD+x2l
P5mOd1EwHBRoToyam0z7YnUF73HyLrfsrdgdFae97GXD/t2W14hmDOUIbB76FMUMiOd5vpma3SnE
7wE9wr7BsxG55EmhQ4G6VdBftdgoW/jaeF2ptGT3oh1pzYbHaTfnftiFIVmnvDansTBW28L18W5L
1KcNfoKaVFxKuNGhTOsf4D4FBsGOyVQaPR1G0PUA3NDBaH5ps1BP/eqbJFaNyFrtRkiE9eXXIAJL
TH40UwjQxsCgsisTzOTdTfITCPBUb/QlbGVE6sl0qw6BiwKpjiDhJuTAs0+apE2InsC2Es1PxPBi
oCDKDQZOMRH2klSfRHlL7TAgJtfWeYRDcR9XnoyaS5eE/4m2MP+yDfa2NPiOeys96ZrDIwvMJ+4z
YnMVhCz2rYdl5tNh/lxzLFPSq9vZ7Vwt1DNzcZywIgCbWjALJUtzz4VUa4sgJFrlBrp/02YxIIwY
S52UB6leH5XK80ik5bwXsFtqoR+NAIBfXr/ice0dIWl/gjXw1jo5M0X5WValXCOYymCVTo8S1YR5
KCCPItfvzchK3YbUb/nnjZwoHYSRN70cb6tJ26ZuaPGSEzGJzlOnqvX+SJ2ZY8jNsg9hcOo7mHzW
BL2AYRrZILWG0z7GqYIR82RAH3hRM1MQJhvpgTxz9HFwCLjzynWMQ3BJ4OFE4O74Spl0AiJi6TUw
e4KDhpetm2N11Y8sMlUrLLjqaHXOQBTWQMnvtCuPybjJp8hFiBdmfTCP2fvhw/5grZLuPBLwLqZi
f1h5tuq8m07Yeg77JQ+7CC594jnQx+8NJSur/0FSxKDF2agWPBRyT9LH/ifCzDZ5bWVqObU/juXK
S+4+MlluuMY6PWQyfJfOK/staGbdykGafCt9m9hk+V+6gHTJ36OMQrUVXpstYafrMiBsFSpCH2sg
6Hh7aZ8U2sd5yHU1aPzih+4Cp1EjKkXjIsll6NOBdSz4T8oNwbY5VA6zabSPQykTx3Wzb5p+PyUi
43v91odWOXL7DWVdIYa4SFdrhXhcqhHtWhOe89FXy7SCjaOUdJoPM9jMbnXAHnXJf+tOEyGGDFZf
UXeiKSmTjTEurlGIVzpe86GqGF+eoPrtkMXQ2AE936OtnTjmnzLMnj8j4rfQVBbdnsnXNZLZ6GPF
mrBW1+PU4rbcbH8yGRQkYLbn8MzleyThHs4Pp9qzdkC7GjjZ8R/rY5mvmiUzAsysAV1Rmw2isQwF
UZDyZKfSX7wawTwuiv/I+N9F/1+vheCngNEeCUrRKkDgtJbn5ZQHYUZ7aSWztUlPE2ftMycOzQ31
azSlzkOJmn+Pr6NphdGkkFg9370ffWhA4Gbyat7PfM3z+pAsXPzAazdBp2RCQQlgayhsrdB+eOIA
gYXgqxFZCEQKuwNjhmnVOhNi16TEc+QynLB2sJHvy76SBAIFUC9Zq3MGLBlMC2N1ZywYI+tejcgq
PLP7LIVmPTsmb7vDl2WUPi/tWY0ldzvDnI+FPkulMnPuFR8HA/oIjRoOzEYXvbgt44NA46syzM5Z
IriI9Dj1gRLNLcXPzNVghcaDWh4pLh45Z5MIKSOja75bZDUq+sKLFkTu+fP9ZhB98lSo+/UDIHXn
jTu7LbcZVLoIECenLp3zJ6AFFbTGYOF6sCaqiAC+RZSdhNb3mpyHy5jHJR/Pgvzma4o02o2rM1YP
KaRQbDtuv+cl6DdWI/IgqKGVbk5dRYQMTg22TwW3MEJxhQk5oahGlJsQ2af5tcQyArIceC/qCjEY
hXkknQ35T86fK4dklmJRcLXjJTLcoUVGZoIjSDAAPIFREsCK+osn9c6lHTY7aYcZH3ePHUyhEeh0
8yhte/c6n/3VYvR6xmRx5Q9DH82kQ2IWpc4eu7THViwDRL+qUhg2jWiZE+l2VfhAlPlDBGb1/f2S
jJ/ZkMoREruOtmtx3wURLT/i0nNKP16lvVDoUUvicyTkp5zKJ06Pi6Dwzohq6NmMTQ4/trif4k8p
W/Ld0DShP7XFBkO7C/bqT1aOBHdu9vvfdCOmBX26NfGmdFwcBmDHANA7znMxnwxSDEzFopY1wAKl
rMFcxZkhyzwrpbC0zSthjit3Z7hAbAxkaAUD0fUlBOizBnidiAEAzOtD3FlwsqLFI1vbLBDkFQe2
PFsvg2vE/0l0hNGODacyTNzylutF/4Kc09T3fIGiXgHdoLaGCHtliCuIH+uiuTQ4BamqcDFkILPt
VsfKUzbEs8SJBf+zn9xW5kovD7zoPxx4YJinz3jjrILKJwcackfeUZECmjiAKBdwcaJsYoV5gg2j
hLmMtyG24pf3lVtvWaH2ItBTlAJTPS8pfvRMJy7wYehX19YsUnkFl8D7qXZTkulawLko7rvlC2Xc
uX03fFDWxyCyJULHVeGfRfX+xZ00L4+EDtqw4GMssx0jz+VKBbhuavhKSH7rFF7msrLTjmw+Racn
0vwMQNXj4qGF7aQUQvj5USS+8zPx9Pbm9J0qoJdYjt2Mqg8JqCJ78PSDW1AOxKCsF7n74aBLK8Ql
Xv0S9B5+w7vBZioiT7dtwS2Vg+3F+7aqHS4b6OXEVwoOphA9D53AKp/zjuzDLPvxglWn++1Ibnbz
qaD19CXCMiYL6l6vbpWXyfXTOj7+oKzPyH3LD+44BWc8qBAPC1dLtlkmjjTfpKPQfCwsOrV/JXsq
nW052t40PG44pi1K7So/MiJRsdU3yRbcAJcp/3xBMSIEoAVXtVhTmRQQC2y/W/TRGbZ4n5enFNcT
twjqRS/3g88el4Rpy3gxq7jlgto80DZ1OH2eaxDcPINlKa75ULQ8J/rVQEEEbUoPM5zQRLqBWBDb
UWhw4Yc5vWjvzxcuyxMj4hvMI1ng5KqI6gn2HUdLwEp9Is5r+a6tcy1LkCuaMxv+l0JnvoIF77Eg
KOQSzT59QX4aOO3ONr6acrldo0x6egJGX+btddgXK2ZTS0P8qRpttHItMaUyk4FnSZ5C80pAnqHw
FTnBPDTVW5vcSGiN0VnOjagr16PXzLccoEp+ykO1sgAW9Q1LYfGPGo7jc8HTRV5OYhekFq2iHx3k
mhX5JnHHZhtV/WD/ozdpNadU7IDF5nn0zuJKcYhtuh2rZvPGZQ6Li5LYQ0LGvmPTyXzq1/oq9RWe
li+5H6MjbaUojUf9LSnayQkXaCyVHnYZNW810AeZul/rKTlFdX+qDqZ1bHZWIY8QH3u3kFpDm0yZ
Bm8M29sybvV3415HVMQ1d2oW03ajw2ds7a3Y+Fd7OXrlVOettnCgu+Mg5pdb05z0bhdALK8i7JKm
myzYrBb8We/tAMx4YiyoTXRT9L94sot7Z7USm7/sUqOo1AxAOdbN8P0SXA99dszYNo90lC2P5jvo
QgUEmsbyi0gWyuMfgouU1vaSjJQ/wljtjxktfd3HPbYGwU4mq0yEMeTSsdwvtc4bjdIXgnJhvCud
ZFDHsj/SWcXssirKOwpDv6PvnAWPA2PmOOn+Wd1y4yFQ81CZznsPu6s/WhaVRhJFwf0ys8IU7TI1
2+4OG6IAkCNu6pahkMCBRdvyI6ls063nFphlmhcFY9CyIABcSIOAH9FN2cn9vCJZQXawU26xk3/f
KsJ7Ggquv19aNPF1sm77t750vVgvjxf5voLtJ55zzqJenzTmRdWOey3IRr5cu/Py6XK9QT2KbT13
EW44klJriwjOU0cYXaxf47wB0UkeNMtVxaYMKr2P9TCEJgCC+VHmX9PFo7E5xXXEGJIBFJLItgLk
rMjc6aPm7lBLARO3MpiDUt0xgip8puezxQHEcD5TwnBA3rQjpjM8O5hKyFPQJlju2MbfbNEpW1PP
drkYfC3dqg/C9I35AwE+dOtEx5XvmUt0H6ouJt5yk2arlmhznrQBAJBxi2HOo2cibTR4PDQxzPaB
UF+VjEe1wcTKKrfeNtuEH0ulqATFhJXkUPz4wukUywsPYNj9eZtcAGnayjqO98djqTSL/IYVnL8N
VB/Is2niMUS8sYu3ThnPQpM1hYsvIQE2OQZO6pSG08+CNb/3rvfKYaMbkt6MNgRdZrfdQSJGAsqd
X9nMbGWa3Haym+kxU8yVSoT8Osw3feldzKWXn+t4eHT2R9eolXlDswEFNrlppw1FPYJAA3vmdB94
+Oip1ocIkgRhE676gqpEq1fh2DL7coJ7EpYY1TnEEjc+aV2pDhrUauR/u6SQOsmx9kVENqkyTTH6
QqVpy8oXH4k8oYv0ElM/Za9Eoo1hUjdaDwl0RQES6Dd8aF8uMmAgKfrngGpPC8J5+drnZn76dSDQ
seY3jqM8Pgkj/90OI1oH24GJ1TXocxdHNA2HwiDYi3qeEe7sexC71U3HBtsPgE8pn7d+sqbu7Oat
QsiVCA8c32seNypXqF0mQvU/Wp3yZFewOUOCTuTbPlvcNgVH+sEM/Ci/Qej2hdblT+ppZeY6tLn/
YQBTeDbg6lg7uPTC3szjpI44b46TfzMZsCz26y39nCmOdLs6LPGBwKoBM8oZg+yLpQZxgATFTz7R
9IQINK/0sNA+gyf9TQ9FhbJg+rCYMuLQTqQIOnwIVBo2SiZVXQQmG4JbrETpd6VvieInFzybv0eb
CjxlAdcE64XdisJ1dZUYfHAqyu6kgJJn7HVbq/LotAChwJQ03jcpmQkYE9ubGk45TrOzYLVvQFO/
YfmSWaHOINEQrTyOZc4+ViupFxLpuYo3IHGR7hs1rzHjtQsTKFcri7uk+/tOlNvT9pw83R5VxJqI
G2BMZD5+gyILcnPF5A1rMrdqKPULFy9e0FmHHuYdWaHR2/St5jB4p42V92NGoZP4h97MqgWTetoz
dV+pVMNW9zFrs1u1bHVrMBWAyd8OHdISYyYBf3ow71hkC/2Rc/IEBApQqhkhE+ZIVUYvEiDVq4gS
Qp1pCYouArkU0e0n/BWUbv89qesFGw5YIl22+qZ81pxrSAlKBxEk/fkB08z96bMSsLpGvz/AfZf1
2vGy0tARMI63tYB65DyYj0VRcEca3NC2AjvC9SCaCsxm0BHfcHWtvnfeOIqt/A70Jg3xR+cM1t9g
0+Oapbu9Lh9pl10OAo6mzzRI99z3uzFbowl7nvcZj0CXwlZuydSnA77rvYZeS0jKs9hNRAiIzL54
1k5kqQVrvxAv2IvT1UL+n0MvI+62SJHfCbw/JJbACK7ldKmEyGqI9kxlHkUOzpZRRG+msYtzdoDb
m3dEPzGtGA+0xjbEgsLwEG76WeisiLUjBojfwNciSaKCAGe+29N92iWbFtM55P1j42khVe5EQ46r
UPDZXAbMICF40JsyDvmALnKuyRo4V9enO9tHQq7cEB68YwMtYhqB+fOkessWJPGvoXHpEUbxdk1E
XFBlphGgv120Py4np+1VnuLegCZrsweGeD2D6tHKjbRlKxA4b/Crn5b3Gw/avFrmWkR8ExhFOK/g
LlR0VfYTtbKS7zHxZm1WZhjcrsNnZ+jNCZF9L8ZdspABXUa4Xt6agXAPgGYxkboC/C8HD/PtZTDf
GhD7UrSyaYSV16CqG/mn9DRkyUhphc/6sQTp7O+Ln3UT4XIihSzOKMxas1n0xZM5x2FjIqTvOaHm
SR0DXXBWfKWnoPfHPM/EJvOmxoNl7cSVjIouDgZiYHllNOyQsrt6IsdOr7UgRcvsW4epgKsEyGwc
tAhLJ+RTLM2aKGbFASOSpuBv9oQVE8mJk2bJ3oEYWcpnjef7JDLsZh/6/5tismd0iLd/nhQz12ME
MHkr+/ghfi+7xrfo3q6IeZZWNjpPPA9h2ecxGHIPGRF+jeNnaJiw2q81BIPJ8gcMFIEowvSklGRX
dUAr2vLz/0i9UH8+C1yHEdyDt45itaynsFJfKbFfBFN8FCT0XQNp1bjQRJzQst/weBF0e2TgV63k
pvFhbEKqgL354p/gd9cAtnNSmW8YA/BxqQBxt3QjiEb/SSUEKvBQpSpvq3Tr4aO6DhtrhOuHRDMe
PK1ZcoW2OxzLcqZOvybE6aEhpuDkePBTlIaCw7B7UO84PGiKmFV+hgq5i/hxcowhJIqyU2xreOn4
uP6vdGiL7ty8Yq/wVhBUKxAhw7HYq02gdxehBSeELX695+6fYahXApnbYiocQXht3sWI2TTvm+J9
jodbemAp8PpRsuPcEyIeVlYTS5oG83KETbwCHdB0YWmI2sUVFmabJgq0wWt6WFxoShw56UISbngB
Rx1becJkF7uNDKJ8dmLzPQI8JFPDUg3nl7AcRQBpau4XN8VH2wzrWpUBY08k/3jlgRZlFxnhS3/T
QuRfIsH/gkpLaL4GAfTIahB1L6vZjYAIddHNnypJVT+Tqk1SAZPBZXBBByeqGNB4S4/f41O9s52D
q1zUZb0JFwKLaWl915yjsuJHgLp/wMNE0V1gRjD5YmSetyFaEDHjAyiR/C5z9qohJmBaHQTeGa2O
unDZHTjIAR6UQnnBdQjaMiBgxm4mw458Vl5zXsMCa4AgGh0g7zfqnzwGFBWTtKYdPGQwlHTybGMN
HC/XGVXm4O2uu98CnVloLsZYrmhV2ZZt646E8stzK7viToXl4Kt9FspeIni2zvsSPeYuKrEd0KRB
kQf8Lo6vWUFmAqRRPvRTe9uegDVnob3Y19VRWVTVuwMMqDthVsHIo6AFIqsrogZE4HrHXsQgBVAk
4TPEGtuYn6lG0LUJBnb3MtPuCn+QqJEzIzmTF2CYHdgf3lI5GYTw2F0YMsh1JXFxA8VMxb8sJk3v
YwvJTEPYKPEV9T6iJQVoUWo0Noi/WjK6xS1CS5PDFFWmIg2ZjGn9QyVGrC0xm2dLUkIP97SpUr0s
Wiu5RfLhA/pYEpd7eJtBk7ih8T3KrGbtGQIfuRC7whCgj7C8xVAxkT/i5ZIvYniFWhou70KF5Jtk
Bo1vhFY4/RcJNrIPXHZpIoVRRv/AfTZHILUuaCM9q31fIND0MfiH06k+LAUauRZYxGV/HbvmIdQP
Kf3wYDVgLhQXMbDFpUzfxACjJftY4dUZHXMX+ZMJTBsrNoy8NOc48tav7KpCcap4DjffZ9qJXnIG
vusekdB2HaqGKN0sLeJd6lyak/ENvzh3WgUx7hV+Q/xoff1ju9IADS0DOegqkV+zrrIJy/dSroa6
v0CGs+DMyb8shEOLDHv0UDxoB4dFkiGBLO1+lMBrDN3nGUAMBvwKPhUFonpaFSPhbahegG36/X7f
O1NkRPdhquHpRGVAL537fDs2IomSMyi1iSC+bB8nMbPQGwnpEeETDwxguQk4m1tebrRoyDfQoe53
8ZQ2gdQJ9EiyAx49Cd/8wtu0kZpXepFKZdpiEnOmaWRB/wUSxe3hU5CCW6JhzYeejsauZH4OCedW
7hwB6EkqAppIgJHxbHT+GmMEB6lo90SsdhQEYgbhz5kZ2oyTgs7LdNAiydbrQ8Vl2lOAUps75ln6
YGsc+6X9904Bznkz6tQ0npf2ONQWJAj5sfjdct8jA8oit+aqvfR/m3UdAsXT9uTt0sQz9zGcBbVe
l/pgUaCVxjogJ0XfB6WmPmAHBIM31LT07hwCxudm5qsZfJR+Uvzh4oahRuWHg6OMcNrMEObKaCwW
TVnpmDUeXXCoCuU1bzfBul5mfLda+eca4kkdhmaDT6747AG+1SCCYZ+UshY0XIo48Z5UHp0WCX8d
cELY7wm4jDyIQuXCO93sY32UO7ecafd6PMZ0ao3vV19pUaV75iWADVoAsC7fon0omSA5wfvyewGn
PrJ3b/kljVpWBTYCgL99QmtjelCGLVoA6NyGzHRYigdJe4iqxCWJHUh+QhYx3z+MffUzNrLCdR1B
a1QyXZBxfwsiPjzTzW68kUr76634TkcLMrqjj8nI2Q7sf6pjnFUzFuybH9Gmi5KyXjtWbxR/CQbD
LWIjxrQ7nd2VES72V1T9fdbNIupNjLh4+Hep3AsiwBoz8fr8aMLdAr6aPaP8MgHiLGiFNsejdcSY
/nrPlP7aR+ZwW5O4wEOuYAMI+QxP13uQSGK2CkrYla/VtkSzSLFOHwNAOK4sO6EHxTf14XGbx+jF
bZwGCkI/NNwEUw14ob7hu4dnBmZqfuH+2uuJT3iQFSVyTwQyTdH9A/rb48nBGtfagjDOOl+JLc+x
V87b5O4kpbBVXJmYXYExHWCi249sTPcgRXR+3ldE7YB2gH0+Z/30my+njUhV05h8jbH8RHpfRoxE
+M0DwIuLumCNLqjBOf8/Mtl10+zoq2uzOMTT4+5lBmyOvbMhXZV9KCsL8B6EcZkMX2knk9alTDPK
z0egWJa1CY/ZPJWzMDw3vE98i/u3RHZAygll+SClYq4mN+u82zB5IWZf9LhPLErb85mRNMX9c7WZ
re112ZJlCan2811wqOOb9i2qU7UPxChN4NBRWevWAcVf7OoN/Rx6Kxjj+0zATjtHGPjzObNGeN76
+eEXBEQNugrJSDe2EBwN+kVdlwPiHbr16XL903Nk+BjTYIu8gxyojWebTCdZ5MERtaeAbdnmGdBm
7r/7a6hsDSXDVhVQRgAaSwRNFdKs/FhmhXSqUsShaqsmWatqp9hFPQ/H+j1BLlegBYduqA22pNeq
13PjpTTEmDJcPFGAr0D/McXoicXfEbglNP4ATX3m7m8n08jWskKlG2L41ahBOdOb6yrLpG5sqQIc
dccPwYgEdjYTVvIo378xxY/xkOLf8Uzl2ZtQcJ1g065ZFSV609nPJrYpooUUGFuP8eFsX15YlfbB
i+9SrwtxbX+yHz9y1+AtsqQeFAlqcdOs3OG81i5phlhR1r7sdHaTj0pOUMAG4wDqKUhr3VZWZLIq
KXTdRGE8bXYqt3mFrgdSjJJePFBy34I10Pp2ZcoOccyCTxFSw5w4ErFw0J+uheVy7pePRbZpgXKP
YEJwTl7yLfL9hXuJ9LdHiU4ES2kV5WyLbMiLtRBjuYwc0pzox4cL6TZrYmwYNGhKwWNzCV1pn/z3
v7BORmtRJRtC7IMy2M/Kejphl87SJlwBMN/B/encev9PWIVQxJbalgR8836UzrcxHyo9ScB99IYa
LJ4UPPaGdRoqbDPOei2gKtEaGzzyyFHRmNHfUtLIbvvYbhIrjP3LKjWFCUmf0oovoSNZcZHpnfgU
9jcCEyw6o0/j/CDFrQXA1GX5NoPiEdwczEy7R+wHWIazDfd9FhrZ6LR8bFHwfmlTEQivEnmnikPy
rddF5KhM6FRLLndRUbBlvt/FqmLxXAOzLS/aWDef9/gIWWL137X2Gf01V1UNgHpG5lLV72ft1e4t
BHAA3uftyehG3d3zE90HX6m7KF8ZGVnY59hiL7UjDEeifWvFUA1oMAJNX33WSVLXY44jKsVqeZoq
FHBplsmgPWRVmz7PA/YiU/l5rtKETIluIB7e46aQsjVhjPKoSQBLTIFEmMLTfZcTWXD5G8bCb0Fb
R5upz9T/h4eklKdCOEOsqp/ZxIUNJuiwTSXjv7AFHTmZWu9rtjM5XEMhMk5/XuLavwtDF4ZfEHVj
U5W1SMaf2lJRobvuCPlvWQ+Q2x2pU8Nigu+NYMgQ9HsxOhxcFqqI6mBJ0mwMoyCbgAxWbSinN/+a
bs6xU9esJ8dlQj1NYdxbG7DzXiCLNsS7sH2vy5zFcnwK6l0ai44LIIJip8xjGGyg7KbBbVhou73d
/4nLmV0PxfmuPONWEkD7VD35q5Xk5tFrjc/sajfEhFARSDix6qWYAfY6iJxX4dyWQP+mt7zQDbu4
5ecxoaBXMJhpPfmqgLz5L4r6hUoJ0MuZgER2cL0OarHd/JK68EU3byTUY83WZUyk5hQHEDbnnfuo
JAdPyZPsbLmcPx1MDpx0hkZcP3ZREWJHuQASBXpak4eeQFf1z2CkbpGKOsrUtC7b6Q/8Vsmj3bCv
71oE0v7YC+qkCROmfxB2pa/MWgWjlpu356vWqLFm/q7tkSi+qp7YZRMZvaTc+4HCz+BwpMyezJ42
Yuv2I2KiE3bcoCsBlaw5g/G3cEEXq2gOv50kQbww1Tryvzxo9CoNjODFg++pdTxN23Yf33ddzaM/
c72rBGibF5gB1dpQAujg14WOjBZegD/QOFNQqp5I/eOVBZxCeNL3fQpBFNnlbr9Ia0OYcJzb+luj
RAoxXkayw2K5a8QlofkgUDNVGulyB8XKV3ihoYue7UovjScrU3A/nL0bUJ24e4NdzED4Kh3Ez9CF
VuY6mO5G9ISWxzZqRHGIlSkSLg4QwNLDZmCcsdNZv7u5K/7m7FAco+L3z8To4q8a5gbVoTJqhPcd
jAN8wavDXBO7HJ1uAIe/jZZph/xyruSoxlsynB4gTszwV2s0VxCAZ+CNkq0A4px8eP4ebwCqq4A/
eNDQrX9c1ZY9n/t+G2bjpC5K2tG6grhWVTbqxtYiX3f/DME3oLH/47P8MgCAu3xiFA4Knfq4+9Ab
r/CxqJPnt2lnd7+t0/KimnvGkrTSfeoyL9ANETvE58iNPVrLN2FwTFoln3cbmXjwrHpn3b5sykPA
5fzQSKVnG7EIxlBcgkvje9Y4uOTvjTeFZg5gIQwTverPh+SmSTXZLqBlLOIpwpLf1kCvx99Tssfo
jcJw9B2dnUoYJStpML5Hn7fTwycKEY8hSXPCkWRkYHMdt4Ymw4KFKEz/G/52JeIgG89uiYZgO+1G
MZLE328bA1Lm0KCtCDqE8AGozUE3ZALrMkbKhSlBBP/RUdVUVKidYWdfXasx7tTsF7MNxbvpAp/O
z3E2/zPq067v0SoaKYLcbmhW4SwNnzMBPpqId0yKSVWHrbeiHkB/LvurqyLYVFoc5k1gCNTKCGC3
vOJXrhHzsrKVMzYeQJ9+UVageIQwgU7qOVCdeQK8fvhrUo0Y7PDnWw3CW6xA/wsoWBlxKS/1Lm7f
TUEz49RlX8LVYnP5P05aR+cdF1hktGO48nBS+2W98kSb156d3XWd8hZ/3TgNk0dfBX7K3fVJXPV9
JfI9r+iP9BhogKaYXDn4a3hG/14ad/1ey3INa5wmWMlW/+REOUgR87U4upvycpJFO0qoIp43SDv+
WL/IaSiMEWNeAhfMG+blQAMFVqremFnsZmconmpFQHNIVaJPEor35V5nMW+7gVOdSwKD4pwyRiZW
hnIr78TKNx/5EU4exFZAo1K/Ut6gE5tOBdoVsyMNfRrP/hgJEI9bs6QXBkI5oG7WNB/GjCwZ4TT1
t/Kgad2kGbBRrpFeHYlxFXEAl+b9V3h9HD/f/10Kx8elfrpH344UFYapmaDCZW6pFPKjzUaBJDBq
8G4fMBsbI4/OHAf+ycYnEGBmkhgOSde+JcL5IgA8dXZ09DbciBiLrgzFQV+CfmfD3MWXTQWUvwOO
3jmDALrpDEj2tTuCGBp1rdDvx7N6qSv2OX4y7Ygz5is+smB7tZYJBeXIKWOhrKG9vYY1wxcVh7Y6
4NAB8w+gxLIJhwGhRpEdrs/0HbWfNYzfBPCE0zBFv96GEFMRprvy8zsCvEfjlVCY6O0LqTtPMUAO
rT8MY+8p/Ytc7oFyqMzwEYQ0WTTv/+2xZLqP3T1gfE0bB6dpcPYnFxwb+QgfTG/eJ7bcs0B5209Y
FqPMkPQPJMEgo+STj9DK/Yd8A39aMYeAbsHZx3YEj5GL3C4DX6R/vsDBhheeNj832fowrWqmZ4QC
aKFGKROH096ELd9kSM0gdKVLtcW1ALZ/kkzIINzFaw8jpR1OE1V/3tHxTvn8RIk03kI6DELTP+wZ
ObWJzkKwlHwcH9uke7B81K3PpcDPjAdik4+e44p3ipUdkWbaIYgmivMRXVetuUwBU6WC81SC34ol
83lTLqJEKTxMEq1EjT2kI/VNiuirYgNNRtEiMHzspYDojZ+9NO/deSKGpZXJNvXvXoxiTEfj3Aus
o93rd1L+p8U/AKLKruXTIIBujn+q/4KPFPmOTNXWcBZUwA1mn0BLR1w/0Q/GIB+tXZMS7dFZb+iY
Y89I57ot/CvhePRdjxwT45JaqaqFa90CZgC6/GqpawOgiOv7XP33Vy00OKVVrlnWv4gr+9IqqIPe
pRIE8o5GzfDR09m955kiAB0FR0gLeYkN7imvWtn6TmsIrdal6XrBWX3YwX+U3I4/dBo/XewtO1Qc
L670KacPHv8Zynw6/nrF1y82eBwRSXDVdSYulyTp+7QHfyfiVSnFzBaiu8bffWPM9yBHI3cz84wA
7uK+zpLA8gJFvQEdIDl+3wSKTXxDbztG8iG+R0NQpVvIWnVvA5yYoboNhkbnEmPmXixxjgeZKiZd
t0YGuXnAYwEbtyjPXBMpqC2DMUlL4WIjJyjLrEa09VGW/xhlSLYg/8OwbwZcBr4HjtN2UIw/NIBu
QHnVXqdxx5c9IhedXoTwyNG3/oCxYBuOWTTpS/RfWhDCGtFnJphUgb5J59bYLmL/yAZEAHgs7mbK
E/Zq6HoO4WDQssK2wj5SP1uUFEpSCaNd5ClTG0WoteO82Mz/+zHT/ngEgbuuqksZ2z6ShfilF+qL
SFFVEgJoE13NhN4heWGwyfk4uUN0PB+d2PuW0OD0Z3WBb7zYx+XECeoHiwTiJhf5Tol1XBT2kFq6
xWKDuJG7m+csLlueBzcyZiIh337dBmnPBktujFdLXHMv9I/PRqM4o5bXJa7N20glB2V1auJwQAHL
SXaRKPBlusz+CEhynugrMioTNJSWnFRqrojpn+w4vI4QAVaHobgHjxHZlfznEA+0+as1iub8dym8
okVc3MSETi49UHGL49ctGpTNq0Hd7TgwUL7LBSwFTiTJ4tUCXw4113T2HArfnpsp4wVC6XUkd3xe
DgeCFDV3bbzP/PcPr3wsDZya6tC1zYz8UZ9EwUaVypNniVQjlDhos1A81oVIw9yX5ZelMN10ohtw
KBjuu4H2nL3y3+ynP2WITqTQ/Q8kVJwmx7Strxe0Erya8J54lyGEr4p59Mr85RZaPeWW75B3rQw0
6YkEmPp1c89eO52M80hUeoxNAlr/0zO45eAhU5d09cWiKdtAJKpCPR+yzVQlawoZjWVmcr7YdJ10
t7UgSNvvDULHOOfdG/nQIjhmVMI6bdVzarO5VOw9qG3gsvFT5qxtK2e0u4b/MHaxbNG6rf2G1jVy
UUNs+4VzlS4vmpOBVnBwCDqLhGVo/q9w7nkePRbVLG0PnXKsB5K/W9YmthnxBTmck4xBoyvAPCtW
cHmpWmYsMsqUkAfNalBsTFzYuRHqZx7PPe2K7pYgQnOaU9fLP9JoobXcDfiWKTc0Qz/1EvCSPYOQ
pQEMl/Ea6f9m1XEdGW8q9n8tB3wA5LIT4ajQ1+DijagTMsXm38jlpAbCs8ErSYb06ZoArWvE60y+
Tl6rYTpgF6G8wpQiRGRdQqXTELtuNUt0PzCrM6Gww+0LyiUIiQfBHeVJVPl99+D8SkLyjDmSKM+/
UWvXj/jqHSfrIbGNxJDr0aAOc4XluxsRoTEP5DY05eeJknm6OmTc5fOVu+0jVXs7ZJxuqaQnSRdQ
Fptmc6F4RuOE/vXZRcZcxZttY2s3iFX99bBdIYnaTr0r2zc/Dk2ZN5dt2iGAknFt4dthyLfaK6la
mdtQXH9cvxA8nw7DMQwex8uz3XW7JhHUxRkroADDbFo1XhSc0uMj/hfeveuaxdTAEQ7e/anVIyyO
L+gtH8IRZ6BMKgirzvp59GftHk2i3IzbNjeLdVw3rsMyyfSXAiLxoejKt+/smk1tmirob1tw9oFg
nJWhJ+b8UTogNp3mUNGQiAhvERkiVhAiT1Xbk32ktBQ3ZTapvamiSqjf5vM5Uq4QyY01RS0nrTEZ
afUq8le1mitQ8mJ7HkQpJUyeIrWU/BwYpMU+ZS4rETVj5H1VDrEfcVEWZshDC712INmVWUA9maC/
v1vY5HeuPsuskT4+K9ntKxXk8RLkBwRn7Ve3cdfIjlE5XPbmj33cTWTo7K+8vDZb/2VxzWhLnxs/
8quPH2tMGQ9UcCiRJQW2nyRDiMOggFaw6aURZiy1ASrcSCBjYq5kkl4Y9AFepEatUp4GCxtc73hQ
xWYeLFierM4UwZLIxNsODlhqQXleGu8v0LWRCUltQYaHT5leda2IzbIMkq9GR9OOgR2VQLViRRDX
BmkaU5dm/Tvtc9B+YjlDULBCVFYWTpUCcEyMIZWAcdi1oOshmTm/UlxGxhFpkK2CA1KjlnN3mIPQ
9s2g05cZMInDZ2nmAvgRYa1K4jd0vLlR0EYPyDtZAvBZq4TVb6sHitApmhRMmmOWGV8PQGTA1SZ6
tuuJl4uxxMW6EM7qOjAC/cR0xVcKgeJn2ft4Kw147ABeU97Q2p7eY4GhOMJ9Z2HcHr3B1xELbInY
NmtClDoTSV1aGcs2IGO+ypy8a+Dq3HjCA3CosfBij10O1vhSQDcO3TPmUSPixw9yxCEzR79lmPxt
BD8Twq02ih4i21JC0ZZrev6UDC7iUvSLwwK4GmjuYq0nugLTFG5znADIElWvWQTn9owg6mqCdPBR
OK/TJAKQyUwQSMDxvtzLoaOE7A9zgzK8qGcPceF8QvRGC8OnAIpvNo+yGhkRDxF9gAvHo6sfsJ7j
TQZiQ1SeblWpccmUnhN2Ch2sEBOIeNiVtSOGlFTiTG3XYBuYTWT77vNUXnCEiIHQDQbH1aLhXDuz
yrxYyPXAZH50hMNqAgp/dlSRdkqa8svsd6xrNjyxIHilrBzXigk3RdXGcvxmlWnSymAXpW7lD7IW
JYKnJzYQrzwo60UQC4PG7KaQZytUaz4lad5Q7My1+fzsS7Pa20iiSPStJcicUnQn5P+AHuW+rRrT
uDkePgTlcGGhtV+bD/ciVw0JXJz3ydYKoLC1DSmJComOmQ8XBxR1nHuwRqce3nSGSD3d1+6RQVgi
iLA3fNabmvOaRnaA2fVH8GPg+9bmUocxAq9pt2jUHLvMI7XACORLCDfTUreY/gSdhAqT4UG2NNY/
W18LCCCfXfsYxOrX+ji+mC89OoM2xkndEUKxE+/wGjMTRmVAsw/92HV4RKYmedD3U8aRncdSC/YM
ovapr6fqTci1llQpiyizYIGbhlTXdHbRTeMgqqQet9grJriwKrSy2/PZYph4EfVuvuxlFWTNYMf4
7fFCb50BWNe9LhndfgKGSOE71Qx1lqbGq+9yOaeVF1j0gXKIP5OKVshjtiiBZgbOa1UqSzoKeP5J
/5qQPCD4Q9mLHEXawsIUoXI0eBcCIK3LxYFqgN7nxaXtv135lsvIXAuQFYLuMsAI0rllaRERmY2j
h5rVC/Mc2GHVljgu4tPZE7Y6MM7zNB6JRSV15GrATUI4ak7eZ0uKxbt2szUxz3mW98eYV3tFbJ0I
X/eUEELU+B0/YGXrkk1mxTfpgVtBllOSBZ99zGGics0pkmJWwDi6zCBhzIUGVUB9Wd9Hoy+OFpVQ
GJ8PkOpLcTLAgY5XUEW943fZJwMTVwFIbeMhCh31eKLfeZAXevCqLe7n7eEyPf4yG+CdnfupZoG9
VYIYsGNNg0qh7WNE9jthUNI/Cvjt/KSX4mB67HIVVSfH8xeTPf2yAnb9MWRJ7mt90qIz1/qFCi8T
EANBqeQR1g9z9ND9jaV0jDWiB8m1F03qBwZKR0fiCguBoJyoQYioJp/0IvUKO72+LJ56jdGGuNUv
H2yfiqL4bYWQfsMeVUyagUwCQUO1KU7Y7JTWW59XZs9ng6vab+bT/7ybMKBesbiT89cXgzhaZR0A
eadV9B0Wy6KDZ/lqY97KoqtWhTAa833qH5ICTP5YFoqm7X53yVCK+1QsvonhUoyOuL0XHB25rxKM
Wz74xy2M+kHl92i/fE32ZGekZMfbKa0InD6ZhOp282rOAw1iVZxpdduWXkZAfYrCdhUTAwND219z
CuUr/2LI8vjCRRhV17XKqG+5uF5KvRACGVPTmD70UhYVkS6zVzb4bq/3y7isHOsxlHfgbahi6Rqi
ChjUeCqeuOyQC0AYUczauNvpGfwVUgZX1glndX6Cfbi1NASQ+DV7PemCi4j8RmOV4/oWUrbRe2tS
6UPciLzeCCVIP8VQU/YH6m+2PK4ODI+ExeQ/VEtuKbVr7Etv0MDUlhKRa5jDWI4BJKkOh3KB+YHB
Ak5btMQxXuXAT8gPRL3Ch2H3hDeEW2oLa7gF/3lDuy1lEPw0uxlx2r3Am8CtDK4SlzARkoHuI6Ng
0/zXtuc2qxEJD6HVGZcDRcfl91OBikscR+gj8fzWKHK4mHh2uCCFsGiiqB1CDFjbPnn22W4vg5KI
EbDJDAWw9dJdyhEnbOdrV2V4J5EMgM5ZbiUIu07kXQ9bzon5kM6eEMgO4+SICXUV5tixASP1y5kt
jPFJpnGzac41XhCZXSrk1wjMitO3TqYd8BZZv9ispmTfJBJZqL8sSmaVsIu0QN9HTmqGUail3RIN
jOEHiSMYHZIgczOPmPJc7X7fWW/ZuilNZs4KZBY+cVv2UVsXplElXD98+Jivnv8IJlNyufgLLzuN
OZSQ/kVTwQ6uwGYFLw6smqJR3kNraLMyKCzMdU8VzmsbAsZDrjSF3xsNE+5Jq7MEACIaVpI9/QFO
20KRJiN0fvqguEkM8TZR/S429myF93GKqaMl6dbYcHBLEdadYb0ewkS9hS+NMs2a445opsHGPZlH
f5cJhxcFurVh2z+itC2S1bmmmecT3UWVJ0qN2K+Z4tnPQkg+76TM+UonIa2CRFQ1JQdbI/kYMeIr
EfjmnEjrTzgGIodq6Mo2p7NgKZ0dLeuAzowxUUIVpTbvyW++OzBWUVzDi5W8D6p+Y5pscho/PzY8
rNsYIyj49uU9osvSHPS6hb4a/65f8MSzU4+i1xzw8STcFQEcCCz2mCEAm4+RwjmOw3+gLYjV+IEV
Bl0al5WQ59yzyf7n/9PBgXT293pGtjXxCbkJhZlusQhWUrNPHTyrK9EDKoevDT5gl7zUesrZGLRD
Ewp8W35AqHxSrh8jQRxot1IgCRqMFo+4aMGcanAOwl80iWk15OSSsMa7cGMVAVfp2KiQusEM76Sa
QqiP5uzGrpoFFGAxlA64L12sJEJ34BjizFgCrwtmiQKqaYqBgfprk23rSiBnjf6W15T4GnSoiNCr
fX/mKSudpNTbbpKgSadj6ViPSFNACLW+5OEzKvonVbTDrL+FpXQObYaDnso8hjnf4ccLtFgVsNYT
ZrWBfNHnQ2kYouF8vIizTSjoSacYWjUKiNZGXdw2LVuXc58H+1qsf6pOOkqxomwNjo7PgKD1TJ/O
7rzcjnRajOEEGwjiwh310hs6nL1XStxCIGKty2sWNRmed01HSxCMIMYF1xT1xP4HunM2nKjFDG6F
926FVGpev5/NcTtAK0zvOyNNewN7OMWuAArQln+YrOnLOqu/4VpQu7GMn4DUhRpAi7SsB3Yin1fT
1snvZV6mzMxATgu3DcSgjifBRj2O+803FY+f+tbvsHsjrFC6Ox+bCH4VyTC/iOOqKqxZPPVLLZ0A
ZJ7F7zdiQz1XKxzr3i5ELe/PjznBSZMn6Uv1qkhc46tVS1r/Y2FxUlatsHsAW92vTmbap20GEOak
rgcAcVwJwApXfnHU3SBSTPGX/XqDZaaOVgtnbYH8hQmpeVWCCeqR/Bpo3Jjv9U7e3/7sWTDXF3tm
HFu650hXvldTBJjeyjYwh6u9IQq6D3j2vBjh6DqTKv9iQeDQIcrRTC8M+dtCfKpB4I0YE6vtHAgm
n1/Ow1brc0xjipLD858ioaKV/f1rPzkGyN1qTUaNE41LqOICOIAI+dt59jGknnspndFOqAhljlAF
YqAJgKOoVcNH1+zfqZwqSnWoDo5zFiZ/JorEu22UVZICEonvfwXMxYCsq0t9QCbB0QEIAMZU1m8G
KycLA85GbH213xy+C/03noPMoZVrlXvm4u82RgwgNSS0Rj1ilieeRQ9BG4sOO48ijPpCs9pN5PUo
b0/QtgzY77Bo2Kn0RiHky1clHtjPZGU60AHGa6KaI6xYP8zJ6OCHH1Ke0IooMz4yflbhdOQojwy9
oIDBFQ5j78GUXZ7cSMwcggv9AokuxD5LlwUbfrfEFgAcDWSa1+aTijCzD7R/7bj3wSaWmASr9x3g
0D4HSyyHr6d8lTBfVtKrvHNeiUVpJjdLH68sF+XFWmXHJ3/oJsAcEgJzUsNdosNIRInqhFj7Daaw
VfKkZ75c7vMuNyYy3RfJ8sMVKvEP495d8iF3ebXqh83NuBjVY1858Zm1Gb424HQdf1lmNaE9KOSv
YLB6r/X5CdJeYO3GX6DJP5fcILxWb4VrCDZUiMLxyXs8Mji2Bgf5HKg6fN4Jd8f1vl2BIYdulICw
s0so7YmFIxesCPcWVJdrVbjfTCaj37Mxwi4L9sjHkavOV4ByeBQu+AKHsNE6UOw0IzFyi9pJTC1O
zzaoFu58unSuOwGhzt5rm9Kkk3NST6v6Cakhs0Ok9V3Km+gW/p8IdIe9acRSBNtNNJRL+AzhFqVs
QEt9Tr/XTiy0jd/UldYWLXz4RZo1veRd6RZhsSWDs0umdnFufBUypogLByBni89cU3UT3zSEYnBe
Pmj/SgpDmLlXVTXVAPIvPJCaQjc5EmCbjiGKm8XHoo/aGNA82FxaiqTBiUxl4xosXLUuOxvgHJ+b
ZSfTqCnR0vCzH/av/3MmFwdN3CGBc+x/9WfP1D+LVtmXAk6wCMt9H5ITK48NwIZG7yt0kfjNdCT7
TnM67jvCT4BuuPTaKQMZyNblf9xlQ9BEgmeAuj6DAEOPZFU8Gd8ilKbDoWcdtBc88K3SCZewQYNk
wk1jdT5wppO3lbrmtrQeoykq/Nnag3fsieNgepxNE8y8KnLia63Aw9a3vsn6kr3d/HRSu0DYjcML
pnesrz2OMewwwHmcTcYHwnpxFAvlk7Ar/zuOivXThdgREF4kYrsjARSWlu82mNCZ9mvYbBkbSGzp
LC9c20vcIXZ2ckvTsKu9Us88XKo/oBexfgYQ3HM93pP/1m4LQLhgp8ULtXBd7LlUFGSlVxK7Oj5H
Q6z9G1S6qXV0dUCtWgIeZ6ySy5fYjbzPCcGzhrZBeHiVSdkAm1HSU7hctduRKrzqEOgNf6eIWUfx
9GCBmk5jyB/bBkQrPoPaHmVvpRQ9+cSq+rcnTkkocR9986unzBnwhGrbFyOu8TrniP33x4B2iwZj
HICCoRANKueaLzfXT3lc4HRe+kgBkvGDajO19gK8Gh5wUJysMhQV26o+FLF6554u6mKYYpPh8dAe
fTJClTb2mdaeRMfUJqTpAoR9+wvD4jyqZ2hsxNz6723txWtkA2hC9JIhWgfWtzOX6MbVlwjpJ7nP
dbIOGp/H1kAp9HX7hKcxQNDR37fzNsgDVPBjU5bkp2EY6QP0VsLt6uAe52rHazoJs4nr3TOaVLq3
sf4ygYoBxHT2l8Dh0S3xs4S3TKihMN9Qgo1iXmqTHGybcc8Xaexek3YFhSGUKehfS8gMeSYOSUEk
Sk9Z0OUSka8mQqgWL8/ts6Qnj7Djd7KakqaP2TkNZrs3StxgcFmb5jW5R3J9s3CnYRhB0rDVbb0K
qILOoH9OTtxRe1IEDuOEZuINaaoQaox8sS4MIkwPZnxo0gnKbLGyn5/xF/XHRLTNgitbEC+5EJsr
MKcCKZBpyFfPgKIMcQ4XnQ0ZBimVfqTFNHde+9YXVxHuiripjzHtPK6IvTYGq5RHTFZBDF+nDLgm
dOGFiZvsKSqXId4TJGOE0g9lnUAaerLfm97xna1LbpF4IRS2AxegsTWj6Bi0JEeE/1S3GybTsqB+
NRcRdbiWIkxKC8+KP5cw+3qWeSdEtQ2RpKgCKWi21PACfiorN3Mn5+pRB6zqJ2wf6dtHGypI9Rhm
7G8Ef/a5a3B125QSx8/9LJOCU0TfibUUDGBFDPWb2BqbZUEN+wQ63lnvtNXB9I7KRDPTxxZ0rVUI
sTeTj9+FJz8fJGHVbozowyqyeAJJkXvZwK9uOKV6Dv5sIyHrvoc8WVPq3Js7Ytqx4lTZicQeYNtw
fReMz1Hlw7nz9Yb7cIe9XV1cvEVJkHOfAtZnMqLFggfLYmxZbW5arbTs06wf/LWZLaoH2Lq1OXg+
QQgQd0coVd8eXV1o7j+p6BQqHaloJZSkv2By4IliiZ9bcRZB1rbT9aqtZYhi7aBlUwvIs+ovGLzb
+G30631kq/P1hlz8hOhB687H04/vVwbdNLTrPIYzOPTkDic+3K0g0BvHVTFTZrpl4uEX3cnvHBdp
Y0FsLs+WrBudCfVPjhAI8hzXNqQhIliNIkmBUaon1Df3Z8UwFdKjrtnlD2+SrrqIqbpvh+uLDZb+
xVpi32O3G8Fr44p2+mnJV0g3BsPPBHC3hjoceH5qp1cAb9oRocz7IOhj/e3/FhCKgg3WNDr1F6jI
0FWCW8zIwzDSMXJtkTOmb7ohN0khH7Mj/Obr39hBbSkpneozCeISQEXaZ3ye1mYRI6SLPSlqjtoa
pwSM/1a9CdppjgxEvU3WtVeE3xKtRqViU32M3+VWbGpFJFdPfg1wBzkK1dqYHtfZgIE6EOt6dtga
qugyH5V+RwhPLGSEdLTakvYukiRo3qNqRLo3qYYv0F+A733fSbiRkqLpKoUn+E3nAmj7RoZ8qg60
y2cSmt1heTfZkp4DPXzYi5LsUyQGY92esRKcvRuXwtmxDquS3h/L1LI8WXGzLRg8p+HaB/YdOFc7
U/XgLxIZkm6B5KA132S7dXUvl0kAZgX6y7li1ZQdJI5LIgq25K+Wft8wtGQhMfj1r4vEYedZirUl
KuObqrPaC8TtArc3h/CpuoiPTHcvmQRvOej3hmGO+ezMwzfnAnA5cQxlGublVqaLTAZ9y8UYUXfm
F+/CG26duiBZiNeOzRVeh9foskZDyfftI99j3rQwOsaRzbGBDp3rOtlXP18rdGcO4/6bi6eJEOvZ
0jsf/gTo0uwMmhkn60wkud+b0smoVwady5Gcrv7w9HYn0JazVhGRdEiF5IHhstmvywPtlz1XXNAN
vZGgKDNy2YzfjbkOxGgPZhDb8879NL8QfRrNLI3GwrzjsENPPpiRyTpDyWuC9ksguBYMvn6ICExq
ZD3qoiAtt3LZdLLRDFgRJyA8ZZmu7P8jDfEpz/Ip7CQkT4PC7hZDRxX8JOICAjaZgdedk0Q6vVSU
/7qgSeEW/r5lISp5urCLgkCp9pGyYcyEDLBuPNp6O2OzUWCy9pefDvT4cCoE+ovoxrE6h/Y9EoW0
EMWq0pqHxsLPdxri24M5/Z0HA/GoabDsQuizR2SLcMAbmhbaskPw7pjRhAqJO/ScT38oo0l3oFIN
gsFRihY0pT72Ym0ibrxotv8OnhrggzcTqxodGy5YEW7ymYnntpTf0vZ4xEBkGuae2F9EvcTEQuMt
2BpSJ5o8HHM3ioMXL9mzwivX/FPLf5zXQM7MBhGGsH/QHkf5ZWDRw+yZeZNKFNwWoZgGEXotnfyO
Fgui6M+gyZ6+OxsvjFGZBOiLRGNZ7Ll9/xggFqKo0TExgHwZCbmxU2CT6C9tirO0AfTPOt8hZJpp
j5AzGmJcUDqEpWcNcsoJFHwlWVEUz/gGFYd1CnaIW3HxKAoxB4MUAz1GEJKST/S6bAW6jdfx/BSD
L9fkUV0tR+lGiDsLwBRmycoYo6b2+mLGkm9iii9y1zA8JSw4Szy5ck0O1x0TZNRcvHlcZYU+18E2
zfWcKAYFCCGk2MNGWR/5hhahn31tDlm1f8sH1OhZYsD1rrmqmVPBa7s7FsAvHrcJpycurHH1mYfQ
bqoKYuQ2gHAUMgE0+Z2997y7N8f8KnGVn3NV1bfzR8StgFit66CQimGppags1JHw/nak8W20s2lA
ijsrWKdp3irfUVtr70I7cUV0p5wHSMyyvmp6C0EmDxXiHXKz4lVNUzqmzZ8APnQGo9Z6YmDXOLqD
YPLSxgniT2FB/BvSnXcX9O8ab/5uE8F4Oy346Zs9enXoj0jGdmwASp5gMhqeEQY45YK9SbGyKO4i
dFSygD7UyHaejCBrmNDeTEbkf7VU+MgdVtBvhzQdi5DDZWl7cRao5IA9WwpOLUgB38l6UpPOJMgR
FuL8gLZ4AoOySk6LbVIty3w/j5V7sa8rhnzgOAnX+gkQb7M+hZ5M0fzZgNlR3wY8DavWqcSQBFCe
Hyh8dxHVgaCZAVtWUzpS4jXsCbBpoAipFS4XKUqMxksBQPforruhz5cX3P6mcVYOZb+kJ10zR5i8
m/PpygO4Nicb8hTBbakqqXjgMtbWdO1aXuiHyFvs8RLPJb5gqfwrsJpKw/aFowivt9DhXjzALAwk
Q+XGorKNcevW11HrtSH/ZZzIILZGQAa7/M3ABAgcsdYqpqEG64jTeWAX1K8KPJVlTHtQ+nNNDFcB
A9i5r3W4eBFBGjDQaIou5RCpc/uuPRXy6acj7ee/Ggo2+CtrGEIy9jB1xLWdx703ynEawsRBihX/
EYK/c7s1GVf2A0/+cAiUhnrVS23jgI9o65guO+BNXe9ap3bGml985Oimom+7azivYAMSW1vheaIo
ecxuLEwvoua0CjDJMhiWxzbiid6WIG96bFfXKcq6X8pYC/xH9JHcJzPv7bhHPcQb0AxBGZ7p0imp
U9kjhvxYPpiOmBaakuekJKIO/uCQmNbg2zYhk99wncvREGe2issX4g/Fzwx+SnJRdtQ39yif8TnH
ka8DJuwy7SSAvpBjJ1DpFXw2vmXYU6+gQe5gFaHjtw7TBSlAYNj0YWt0MjZyubiGQLliPyEUnoHK
ofZA06eGPeKTz+5ySU1dJgFBOjGuIN7I2gH1LsGgN5qKuQ8Wf3O/8U5r9kRk1lIZFHpuSYzSDVyp
CFCoXqyckNC0iAehurKc5JyD4vnhh0j+XI1jnFbbGGNIUUKMAM2u9CBUv1gwG+7hqRgcnu0TXRUg
HvkbtKrp6Gfl2kKfhexb4IRzxo3QFtTI+S1cPMwaxhvM/2wzaEQ8b52Cq8YQYOoj9Qj5N071DAfU
u6ZQ8W2swlJoA48hvYe/4w8TT8ey/p1N+AFRYxleOjX9a28vcvUNZqfxMSi8XTeJS+Ke7D1HwwQI
m+DkZAyxjbTjqp6njkiIQMZAH5wh6G0+THw9ay4kwyZPNWahe68gbdBeigHtxNnyDvDOVoP8GtBt
vhi2i0Z5T+e3DnPqc95BqsTfIe3qxM7kt7pEmWXWOAIPEcA6F6p68x6QTPbvU5t8q0lHS934EGn3
MJLqj2JFICNEypv+UK0DuOc1s68EHEgXf6ejcJaYkiy+StoC5SxiD4YCtCCrNtZCphwzWri+qSUZ
dxLBgzl1dWsR/OJEK/LBTKAXhWVPJfBhB1fESA7zUl1HUM00AqmyGIJjcd26doMo6dIdJ5falJQi
mRrO2V8Uu135y6RY1pWfgHW64WQctW7+Zh4EU9E8afom9pRnA3goiCsjM+DTthUTK9SABCWl/nJn
0C25jT69ynHCbM0JjU+b36XKZj5mvtxHRMUMdGLm9SzBtbAncARuuHIidOoOcMIbL+YCaj228zXb
N5lLgXcBLRMtAAsegsGoOf9JJhZULUNVicWfNdrnF189iIXdvaNwM0kflMwxvK0KbAD9RmcLgvmr
ScbiDhugyaW1jm172HCprt1DoIttdnORdyKC2PrvYcHX8zJb/+iaGGS24z8cGaep5ltvfSEhWedt
RQg+24b/DBV4bi355KhM+1NqJ7aNnJhIaf8tLvGqw68WTlDJOqORackcBxkMiaK/5D14W3Nb5QVJ
274njM7RJuzfGOt64edogPHiWH2OQcZX0rMzQv5cmpprLeQ1QbThp/H+BQlGgEE4gm/jxnYX7T6p
s+LxaS45FtFdKxiKRi9sovEQZgnY9IJltGUppP/0sqWqpBJeaUkE3RVxiec8n6gijjH5CIjTEvVg
XiL9GrG7kHXN7RHF4Oo4bP0KYEPEoRcntgXeUfYVl0nUehiEiYpG6R9ERoyAffC9o3EJIHgEh7Y8
zfTGwkvi4/5+LOL/xwTIJEkK/uY8UdqyqO3/+pn5eaOloG5SZiAC89BHdgM726HsZkEF9Xnc+AAB
TVPfWKaP4vzymwbKHcYH17rirewVPRlWQjA59NCCLP1BdJoMHN1FIIUrvul7ziOwLMnOcEBZq1jd
ROdcGRILR9FRglbLoF453rh7d/YUvAVluLabt8ZdoD8BQReU8Ut87RZk+06q+CTe8bgkIwuUcT0F
kW9H3a+eqvggKTbQnmHSfApYh/vsKQjq/7NEBRm9+M4p4NFASn2FLBkzPF41wZo+32FkdcTOq2vp
bAVMpJpBhIOqvS0TN+lkcEJ8KkczWSbAW87APj0TFt/CZYAstTDmvqsySW92cRdZw4FWmhYmOUAC
Jwbv8D69cAwPJLgZlUJvxUPDxQxJPbyKVaVt/CxvCRqXYHpgz6jy7CCco/QxDndDrA8ctTXeqjsP
pd/vO20HiiIjnHlUiEQRpv1FQP2CMmy/ibxQXHDjdZuiNQsDNaJOa+7DPhrxxKtF57dMYDqYLtnG
X4bsUHVI88dkcpNVTKVdA3SvV+cR3PWkg+/cFHqfdhAysygtkJbQKF5UJ4m60bp3qEQHj/WmwH9z
K8lBr7UFxViLrQt6asRBjo1NAbXp8if/YhXIU8n8TMWyxQcc5u2EbzaFd5BG8IaI8b0nUl2Qz72G
66VYS8t33XSRjN39RHf9u/acwWjptODfBvPkXOo54nMHFrhzvCt8QA2jyCMOQHIMCqUyJPBQiNap
OTshjqeBf7BPH57m8UlqPqxIeG5LymR/rx2fAgKrT3mj7T/l09rwnRnGW0phsr/RTCbybQUgGmfd
D8EFZ82CjreIIA+MAmTlaQpMCdScZ8YkSDuWQUR3qnS6n/q9TOfAj4MXjMS1iEmrUX8+uLHR4g2g
OVzLN3DhQhKFdoawW9XkswjC44lCdD+HYoqSbiXJBWHA5vA8OdXwMUGsEW4tFsiLB6ldeeIzfO+w
UohfJJZX57t0owMusivwvgVlZFZH9P6VLGudWDzu7KgApatTRu64jRGefjBEM6LxRQD3N94DiK4k
qKF5Nd1eCOP+MfRcBHxN0CGrTtCgar6n+7afSJD83a1uMjDWApZT2vZ4J9xPmcwEic01Npv76dax
zE/KhIeF3jPw6VsJDGyC25XQTIUuIhmMFjcFv0hZbNNwr3euE77FZXZGAI03iyGFaYJHXmXwTrj+
VjEuQdJretaUdDebWt+An6uHLBFda7qqMqEJR5hjh8sZRgxmLez+hD4Cvv6Mm3dCmyH8cS8oNLc0
gMBBhKk2PqATdVK6xN/gqyBtI5VThDd9ADHxqWRALSenpCOq3VJWgR+qSZ0FQe4Y2V01bRIXKQzK
ieh0V8p5UY3lz2q2M2aEX2vnwQCAvvEzwtohleCauSNW2dxcKrcyNvBpNDDFYhAzHDi2Xy0lAmS1
QNowLb8wNp2lI4pURW+kuy8I18pR0bqPay1Ad/m+YsfkznaMzZDAXLkZjpVOY0JOv1EA94VkSAOj
B94yzqHj8ryWhVzxEdvIed2e+fdKm8kiE4I3DFZgfSrKB9YqAmj5wXNbilmbagFKHuyz2vgQyqTO
mOUBk1XHW9PsEz55OIB4jkYoERN38OBr9z2VHkRcSGRTKEereeHbSs8J3bmJUbHG5SIENw9Wr5ye
E/KTfjZWsUz0Clk8RUK1s58K3B1CLCnyp62HKiPNnweUpW2xxP5/ojNx4MmN4QpDk+zVXf4pHhMI
Bx724S/dAep5Oo+1vHlkCAoId//oRu/vnhtVRJbqgiY8/73mE8Vy4WXRKv6WdVlHQMcmvGX88FYx
L/uF93czgaR02CR3kn+QdrgW13IlTR8AKyP1+Qq7HYruS3bTqYJ8GEZQ1EYVb3N9MqGPYvyA2H18
tWgCSt3Oz70Z18YNxWZw/+djAjcUlPY6u3Aw6HXgk8acvKU3S4i65Ouil2iHvRoxM/eq3Cp7oyrt
xXB/OOY+YrrvGe8wXJil228WaTAm4Pxbbe5aSqSndS57aE6q/Zr9F2kablachdfHz3o1S2nTLnCI
KG6ZrpK8SXjvuw6YMF2KkIQFAmSwTDJAR/m/9ie//F3310G1wnYWuUA3py8uIp0jeVtGSldiNnNP
Sq+RRJg6fGeJKyOl1wm6Wbr54M/oFRB/FXVuzbwehtaYGQq7NAFZ7YUFvMww6KdDEYbHogZEce/l
ldUtg6k8Ty4nhn5mdPFH7ggnzEoAgY1n4bKVsWegVybOJC228LdRkry3LgfjEyErzqvIhFsFNF9u
b7oz2oXKL3VuwipQrMMeSRoqdDgGIYsa+1HcnBpwle0Jz7xsyi1/UAXr48ZTFNTdh6K+rC57HsFb
3bahiTukpAr5FB0f7yYzFagVFCp1S/mXOSnV69MbiX83MQsJuoWlm8l8jXyyhQfol4EBVpTK0gVu
NC81nEYxfqdiPaQF2GnIt6ttRu0w9GN8/KHNfvdfuIO49FEvorl0P/PAMVnbAcXyOBD+VljWh3wE
Rxwqec9vH7xadTYWdwazNK8D/RWKWI784W/tpwwC+Ztjmrk2i1tNw99pTOflJZ0sh2LS/qFne2j4
PzlCmHWFyC74zUtEMn/XjRgOutMCXC8j8K7xIEv+WmXyCutyu3EwFWiwoft257AyhqDJvFpJg8t0
AO+UrtyH8nVEwOnqAl0lg2oSZtfnNUdspSWikq2m88Vc3WThLr+mA024jNSHPjYdtWQ8qTWiWw+M
my1wLau5aotgekNA/4FR6RECImNJ5gTTuG9Cx2FB7P8KV3FA8vS48NfLREwE8MtJbcAfQ7fOwW6r
m7HnZ0nxCWpIRTUfNN4U5oxLo8d4ndCoEt2JEBEgx2RRzIS072JiqCRDA0LdwOlWbnffaiWD5zGq
pM4Kn7/AY0JURe5ZwzmfR0QYAXeLPCoYLQdEFw/LXThrIWWEavjUoNTJw7xApfoDEgZ44dw8l7kV
KNgpQD2PKXiH7MaTF3hOIQF7guIb9XxICwhNxAFR1u+qMqXfz2VGoTaEMyxIgKbniYTs5ZSBqo9x
7nxjTa8kjhRdcw8FSF7NF8SWrO7jhlzetEKINea0Bx1cAWSSYQpBKM1pwp9tDjYPMmQtOxyL2Upn
IPfJ9iujhtzT8uev2QcNPi2Ge2lknYb48N5afJqYo0FmLbmP9urhFynh/h6tG3K7a/qjrjTjP6Nr
EzWWmTblRt2DZovKJ/+4VyFYJwYIMlZsICXHFV3P2ICsboUX5dPUqCOys6CTR9tCLPiBOwLKLQhH
W2XYAcGxF7ZFrhFSEoRD5+dgsYQTzIVriY9iUIE+NatG0B1OsCXOwq3WbEbXuFwOcjM7Aq5AAk3B
Ma3QnTk/htIJoj9wtzFaubMNUJ8eocEtajX6W2cgvAK+S5oVY/gjnoOsZx+gTIdtu39TaCMi9t96
CBIuceKE22G/9HXqOP4O8m8er1FVJ9wZ6Yt44ZPsg+T81XF7GuBF2ufiuBLlunLDsnLhaKMAcbI/
Ar/FIKRsh1hSqxfFtPB4kR8T7by+YfB+RLxd2IAqfj/MG0TYqxWagTFSI9lE+9WWRw+x1bKBrXAu
SxToiESzm1g+krKTVvkTwbGorbLAlHcG+vNmBlQyr7bHa8qitPNS9UF70gUcN8z2ihld7yWx66pc
7y3mzhSGfBuijBG41ZQ8tjyXEUM01uL4bMnykcL0kq7PalJFZWRPKtIKA7lVXasKPXHbzGf04yBe
sPtLWX0XRnsdgC6ROjcZgpSpwb/qiZr52OMPtFICTWJ278iT0W/qDGEkj24a9R6SfcJYoiqB6HnM
UCl703lnPh4jYCtSeCrHwEdfXWPYYwjP6otLX6LfGxnpCX7qRZWVE5BvBGoHpFUtLIuwrtsgYyEN
/MTItDsaP6LQnrGSAdtytmFVd/aE/gbzsDf6yGNKRNPQnBx6nayo5iQmqdDOnmCpVHAZov8jf8Y1
r8hNB2VABjkoss6f/UAH/X+/gmNNljLs9sivLLzxmalZP3n6b4s+3ZAsIMqOrBfp0F+CE/EOvl/6
bSecs0Gt3rmAeBmfNvYau/4qQY6DIB3HYPZwdcmQBX8VK4g7YrUz2+f4ye4e76jnpN85Hdyz0Ow5
Pvb/19nBI93hkrTr5BJYJKgZ/JjSFjSuNl5aH6192BpXhXdR4KzddQtTEN11K7/13U+0xKuM7xO4
7cCxYo2xeKFdyAT1RxVZnrddxHo8yCFzb+C4zQ689l5QGZM4WZTO1Pz6vz8HyQqk9neYwE9ffD7L
xb1EpctcUOm/p3xqKkYIr8+FrQIfyI6CLwQPaTuLTm6uoHYwgzk4TxOj35t9BKRiIrOJa0fPiRSe
9ZBl7OqpQgh33Jwk5zIqBk4uhjZ8FjLV4bfxavAuQo98pGHIZv6p1D6zVa86v4J0c409tqHPMK35
Rqncpg+d+tk5Nv1sZzujk35vBVCmd7WKA1xJZPTMnzy+AxGYvk88TJF/9c6x2jeCv0VIHrFtYi3u
Zo9U5y7KV+FVBfn0b4Cg+401WcrYzbVNav5qpoYRXB2ltBieCEdgvd6BbYP+LptD+VQI5No3oTWI
r9VNPebtUmyKdzkoZpI8jS/Camc6mki50VfYOjq1PWOcsr7BfwJBtD6RvE+d7w4sxuT4VuuwoK4B
VUJqjjOgHsS+qF6NpZwaJr4yY7HLULPoi60Q3qoMRYouGzchv1bq/HabHYZrHwSnVhUrTrJZvXec
0/RhjGXoss0fmlpMPyFzbHPw46gCnlVr4X+/vHXETCbOn904I7zTOSKZtQV3Vx/VvHstHHIvzXV1
4rDAOejyBsPoxGVADgF2KZ6Kb1U+T9MDbTYCCgXAUYuw6qU7yd+KpHr/gjvVnBm7zAE/7u2dwhWp
RoiC4hahIYPvDU5UnvTc2SHUjo3FiZhGjjpEll2FV67FDNNHNcUj82jQ2ddZJmLi7WR3IdVCczSc
FxeFYyAS+DYqliPeM4kgVu/mqu5iA+qz/zjIEoEiyGX3YSqPFbkkLEHS/VShJj0/Jv8Q4pOiKQXk
bcM335nEAJD7ayQXBNufIeRvzG+zdVYx0hyd9nb22kCnKfVErXh9ernsAO1tysBRhGt3dQIijY5v
knT6NV21M2a4krKkUpk1UpWJ94JjIRjGDy4l1wlDo+EsKDxVgrLqeqx2sxVHYkho4P4dxcWsRBrD
wnElx+vrrJsImKhHGIRt4gNgX8aZMJ97gng31cGGJRH74QMj0q92lON4plMWb7dzUnagcq8GFBJe
BwjLhUQmgJaMXftHuCYhe0KPHh8rPhPechD16CaEHWvwoE5iyy6jpn5FKy2mwI1YFoNRuJUnOxMo
KRlwCzJNqjS9+FQM4lzyxjF+SuONeUp9dvu7XJMi+uPI0n0oqlS4uIT1GcNZuMvm4uYtrhGailNp
2RWe4JdJ13GLJEdYzqFRRkDuHAnmvv44lWTtYyTA9HyrsBCtDs9UUKqeErkfhUBhm2BuIKm4qGp2
5HSD1up1q6ERH97DlPU/CFTLvTAkWipOUaJjeU4eQPTDsFjK7JGWwHF4WeYm2/qD+4ccpCGOz64Q
o/gckVoRb+62MJQI3MJG8YzPKEz6dv7KuormOuuHdt2PE/uILW7TabcPhwvHL0lWoEo+iizNW6lm
KPyEFws6YaY6bhGwrmq+T/d7lKILSW7+bEF/r090O/s+k3xzlSo4kVSymMVvjPmbOewqOwmZY3XU
6PdrbXnv1gGWgnuWQFBC3sTt8aTd25tIMLMUrzcfUSnZDSF96C14yzYrNkBS19EjSr18Qlj7Dh1Z
unm3T4ReCtKOOZURECuW9LMfNSSsB+d/wN4+zHbnlJKvIqy4naTs1lw+KMeWLCKk97sPy9YThkPZ
AFzuO8CoZexTN9XkRVjBD3zdKKEnTEcKbzUJ4M0JriZzEb7QQOb/YM7kttZmy5w5XsYR74QUSonm
iMjZR2FNkhJGUb0748NQdd88qwA53LvAppf5RDdU8KFZZ5TeRF2UobMs6i08KoIQDcQVLXcY2Uk0
/RebaTqD/Mx/d5FUTLp9/MUVfhBSVdkwSfrgr8qt7g62RlOhaiTVYQGf1+udDeeicjmzcev6kFl4
KB5w5/R8PjHcRFpIcMITWMDd99Ijn+wMUGymGXEn6UvrJTHuXsiQV+6phh3yoXk4hSFMgv0SIDLN
+kEfVzC7tr4BDUTcoDuEuA7ceIZzAWHdHzdvqUyfSsXmkmr5Disd1EkVqK/LfZ1osV9awguHNPVA
HvFog/NfZVk3RBBklO0kOSp9T4pVm39ZIKtXDxRX0EBoFjcBpQ37aKQWi8si94zl277kU6dzn1Mx
kSMfd4pXqm+HtI38Yy12OhaW3JJ3yxZwFKGAi6VMSVfOZbJtqu03tsneAi14+9Z3SZ5o+/LUEZDt
oCQMjSJ3Li/M9uUtfUVm478hYZrB0fZPNOc6yVPFKtZb/j6h3f6QILEGk0lqaHG8a0Bd+2XzK2ys
TdXJVxFbKeNvtkOnP+SU8bKfz/yzMHK/cjT3yx0oXpZPndEJPKdJrwCi57SE0wohg7ewpBB1lpmz
nOy57u1GeIVWCF0eY8TP5+kKNyZawkGukwJTxCYVynoMbjFuiRRdDy2+PLPm64MsSSF9kj8uAH+J
0LH1fQjq2nNNNehPJGxVg5sYgrM/uFpmjfuAaxbZhaRu+8G/mFL+Br/MneWW8Rnr0tk27mbLAklP
KtHggwvQSm7Qjp8nmn92pPT5yi0NORx1LpJ/SHFjyhH1HBCZt+SgYiqSyVceKt48Wahyx0K8Atya
Hnh2k4E+/PHGAsQ8bmDoRWdji5pdj5ztv4UO8cwKWfyT1uXeuo5Mi4DLrDgj7rWFguGn3riLF3KP
e7tS9br7ZWs9qlVwQcVtnPfSLdx2qeVhymljKE9LvT9uilPTmtfZH2CmLsdDZwpDutAMHsSxCXbL
01kY3xQ0ngkI27N7khG9om7Fp7eHsxucZtDrdcS8WxtwQIn/ITwVJHuh1fCjvzySkFatsm3K78ZP
2DBpgt2d4bJQse4RKywkn0XpLPazz4FzUV5JSsgwlgv1Yxp/7LlBVYTpv9MIpIDyjpkt6RBlYaUM
G6l4yIiKj8uaNz2gxm+VFJ+ukhqUH6ScnatZ0PlLjI2xiJTjsMmrSvgDaMcsV0uVVcODojehj9ZB
nSIpHUlL6aw1r7OolwU6XFOTat4RVvg6yokVqtdxWrlGbb6pl1doiNcdT5AtlI7fP+oPcqsAie6t
uVdSek0Oxt1qSoB4hl3BNORCkJvkOlbXtSbUd9eNYNNj+LQTWTWxYUe2OMro5IB46KY3kjkBOlbC
T9ADl46Tg3XpJv15mlLUSzJNBUn7l+RERani4Wr3LTzA5Y64Zo+ByGWcErWNsDXSeNf5rMZ+2utA
H5+0cknmIxdil1Lgc/ixoxBVVz4tI6n64p/69EUNjI/Tn+gvrBcnDODYIVjUvd2CRg0m8PUF595B
eEqhpiFKh2ip30aD4gm0BtKzXQ+bNajdVGaqdDQgRqDUA9+FTgJ0gTUcsjxBJuFnGLuVL4kVrtfk
krDJ5dOv2czAVTpVFu/19cukCoOMVt2FyJ/ZS9/xqhywC9OZDpb4ylF6v7lcxhfpjQbJEZayKD/4
SO0bhq1tzWJghOuJesHfRdrwmQJuy5aoZpfPX4FlH+HypJMz01w7QtrrEiyIQHleoURacZjcKAB2
KYmaygQw1WrgLH3+lVhQtHXY8RUezR8pDs9t6vjZy7S+b5ylUjwzRLWvCwQiXUS/EEkWuabW0ZZi
6NgyPsAqgyKySfNNfCPuriGAJYHw83rRwRVf5wFeA2WQYSa9cqFhHudM1OdCEd5oCzh/mtLkoseU
Jw8ERK8BO0fVtEJsIjDyR3qNZZ4cIzeKBzLf1GnBgVGaEvb5+la3I2LPLMhcIJvk+UHws8o87Ie3
EvxruOfEJsAzqkKgf17wbcS5cUYFMjn6KKgREgv+xbIxWv97TEE5xPJ3/ynNDCSQoOCnblVj9MaF
Qacr3B59CnwMTocizUH+QYxitZIn95mbJ5RbJG2Hs8PSiDk0fpVj3UYEHEMWbGhdkKS22riH6fOm
YhqnOiWWYr4751g/6RhM6N41E5kGRXnhVMIGE75PBbXg4JpW2rK44B1NaHzz1yz+wfgfklm4E0kM
S/blxlvsxoW3u8hGyL6QK0XecAUqpHu12pPepnChGAztpjrCbtpgm+0/xodY/C1WqPo5+CR71WN+
bTkUpJrHQCxd4/yn9yedlVZaQNBabafa0gdaUpZDlwVnn8valpx/hJrXiy+/4r4nqbFyBCIKbAFi
5M/CnofgCcnftcYnqDN5QO/Dfoaj90zF6hg03yv6lGGOUhD5WhFNeLIjA97gPMgLMex3hpKZ+aD+
M/hkm/lo7+3xdks75fozFRyRX2dz08IlOmhvWY9m/j6j/S20asAw9mOV8xo5+9yQWc23Kui6Kqvl
SRrur6KOFEYvwbpaiYrMDwuijC+pQ1UnFAvNbQXZmY2qCteTWP7NmEoCc9y5hit23Zo2x03tZSco
Nkunj8xpWUUPj4zN2ucEJ9saD42ghkUCbHhhVA96KqLf9xi0xjKrpwvRgCao2+H4U+CKGbCIkLCE
WIUHDRGbFPug9/skAYKS/fK3TM1agBaU1fSA5Y9ZmYYGS9LENs5/HoS/mw2pp9muiBk3GQdxFw2I
0VrQk9Z4uX0iFyThwTZRYM2teq1R1lql7DCZBlSiMnlAIogVxfifTKpG90leC0fwpTiX++PDsUPL
uQ6uCqKQrXgxQiFoUFGDhO+7j0wFXKioETgiUtDBPh/GNrrdRsi3Vf0zh/cbbTM3uPXGHudrIxXz
zBQINK+0uP2iPFkPQxGyKbYuDCqi5Tp3pLbKYwPe322hU0oYK0m78G1SN9uYjpZwnPnwcvPLa17M
1VmCHsOB8nZjZxZMrU9uZyth0jO4L/tGF3Dt5WikO+W7fTN59T09sW15mMVPiJR4tS7tfQVCBb1T
YcA34tDAsiwF6Dyqzl1uLowcYd8glKT3oAvBiDY9YsSmqPtpC2xaLLnbNDylR+28R2yZPfkxHK18
86/x6IJwt4jMAfKysMDPuPnN3kr6+dkozUU+/M6alX81EtXY22HSqqjvI7LgXcmqBr/Vr/o6v+1u
yIyCxuxqrmYBNaDhPYxheUKvYKrxbGHiltePJd2ticzP/aPjdzhEzeH8f+gY/ePcfritpRsphr9/
3wJ8UGn6cGPDQzBxc+Z/bXWLwO8IaxlZMmNqu6QAbkwFq3/jGdQwps0fDsT48gExEw1bjTFakiVN
m/Sap8WLLMWEcgDZQ8KoGGtY+knBvwQAn6Z2Zpz6FhYsYx0tuMazqNn/T4b++NKQkOZIDyCxZZ/L
7zLOzbkwEaQjEqoHTWRsWswAOfJeqO/X2cY5w/9g0Xr8iFSBfdi19bUJRi9jpb/yrfoB1IufGc59
RQbdKU75dsPy1O9TC1KWLDTR3kJ+kwloEmhqAlO2zOF2yuY6PPD2OuJl+NKkRKCYG/PIgNIP63c4
WXW+DsHdRUjuiWq/1g5Ck43izbbncO8qqVjcaaddR1aYTG+adjtnSF5xQoPhoI3YGkCMvBFb90RN
6U9BZQ+VZOTNElUwu9tqnT7GcikTTFf12sAU8bcUgVXb3BjQzMXfJxnbK1R8zDXiARaSUyu7HsOW
DWrahiN2iphYvZfLy2iZN9K07IpPCHi6BhreXbcekG6mb6ULOewHT3KniSjpAv6DDXCTibPYuOu2
tX/nFIwrrZTtsQ0Wllq22ikMD3mKe4HmVEt99Kh7rK2zQOmIL9lXShJKjwybXlT6HgpaTmZPuW0/
fUUT7roFC4h24e67tTQVmy4AveWK60MtJ7RiCae357wvdtQAHfsgLefjGFxC286RTV+xRninpZW5
EBQGZHbz7FxCZbv2T5KRJ97MMPzi17qXR+WidJBE04NP8EgI2QbvAxn/REFwng/86KwNANasOSpN
rUMv/T+Jv0qjtMpD32xnes+ePHR80LAaYs2w7TeAUupOl/T8W1MxOEgdzb4KBkxAnMlyx8BGhGyp
VNovqC/dX2Jz8D5jm/DT5SSuOG5iadlzPsW/3sP4/qRHcxx8/vBiRZaAuSepObGhQf3kk1NRNHWa
65UI+mwr0w4bA0mR9ROLFjraQBmFxM9yJrIMNkIeQa73sRfyaUBojYbRase6xwjKF7H79rR00WAd
bwPztDsTVAuE7NmSIPGOkL2w6wkYSxfNSt261K3PJuiKfayTY1Mtwe1WC3klmqPVNlVwg/TwBvVw
4GCPb88O/wI4gO1roHgdbEf/tGCQ/VHMApSXX22ATas+8DN/at/866ayvx3ch3FsAlFNFPpo7++J
LYCbKQPJtiVnZD580LcnOU9FylGIddaO1jEZc58Jqcw46eMGS23iADvMe4O89Tpp/qg+7Eh4VKXP
OzrG+XZ0uKlRMj1VV7dDoBHcFYKX9diUOjaivdUms6hhfAMwRylHlMCMyfwrxZJaYUI3GlWZmPoy
d3rNn5AmkU+KELqUozlCQ0C4Cly/HA3dsAuynX8sidCc/2Zvw+1hpqLKECyCxCA/vK0BisF6rWyM
vsg+rteQVIJ5ZFVHSUGKSCyggd4Wtbm6YE7GadR2OGFME5oN3fNTReQNbozd1sOUrLQmR4HKE45l
TkSNBHHhagUSBlPcnoXe29rvetkUcmgQVOBQUsGXm4iSdLtHqLOdSWkyT8US021sdrkjuDh4CD+A
xhZsua3fZ3tAt7esAlP8aYiOTMSFPawIbEsnlJDepCFi5yt79OrcsSpQWUd+/sYC9RuPVEKz1ntF
RALte6TgDv5DWh3zVS1l4edXEB68ODUhWHOgF5DTc0zxL50gcDAbSziHTxo/0xAuaa8kx/5yCr4f
TzFIcsQ8Ip30mWPQwVNRm2UE+aqp5EDKjRilHLzq5U23MIBvkbfIYCKPaZVEr7x6i7U7Hm3uBSYB
jsg3R2rLLgTZRM/FiGIQvJaw8EmKxrfZfztg1nJ4yjf7qP8po36Xt8wZbuXJP7KZ/a3tHCbQUUKq
D0F+MiNQKH8uKirD6wFrfSYSz+94iAWC9KXW/A9mVknBibTOoOBoGFXCKUTAuXUrsK0qvy/EoMgL
4BGvxoZx+bMzgjUgzsyeOYAEGVFcAw4sbOKhkknyV/05bgqKUUYwOqqesBsTZtfIv7tMXi84UbND
GONTebvLCATH0+nDTEqnRt2xg7DmZmu8cZ5mZi+OA8O3wZNpQk868IvcL0KO+JewpauN9FdLhUMu
XPXVZKiu0SUk1RkAo0I1AO7VlQiWFWvYvBA2aDkVO1zYtyE5byxzAoqqeJoArWXQvHnP12lmsQlA
X5ZdNaKFlRRDw5+2+V1PzPflmE2z4RUXRxzVXQ559mVD0Uf/ZHjrCius8XaBJj2c8pDvYPWfGxtZ
Tldv3FaAkHtXKT15b7Y8jqqObxDpBpgREoflM58P3Gkkdgy2iakUHT3mHJqTPcH93yYLuX7CVSeE
E0mhJ72emhg18PPCsdCLGGgZK7VPJFGzDC8joFKibguYXIqOOOTd803uw74/B+fOXagoFtmCEIwL
i0qXUhAh3Zw/iz2rm9HVxuTzTZ+GgnOIqOIy4Ewe/ehYqH2NxjaKrdSVeC/UCRnyygECWMB89qL6
0WsblglFsiJARJUjdXQL6ydWf7faXt2lcg/ChoKA38++UyP8AQ8NGk8zBOlWBRHV8Q4oYfnWDTk5
q3zz5tsfNLKgs/Tlsn3olZdn6naAv++JTSfGpEApYXY6paQGbJT+N6F0g6AI1GP5j0+ZS7W60DFo
WVf32PiqR6r2mddNqr/BXSon4EEu1DFHNG7LHFbvO7X4ZTA+NaP+p/ZKuSkGUU4bioUwpw/K0JgT
dc7swyrnWtCjPVHSMTjlnjTKMye2bCI9xdTIme/Y85JfDO31zElHhwdvacmQmb4S/MzoGBEZ7JJQ
wSK8uNqCFjPTF/4botY9tExVdTDBNVWGdnLD9EzKD8cZ2wx/XpmL6svQOU5DbJPGMKLelySFfBNU
p/aBccw432HDQFC0hStygFJOeCl3iRLQ5xtWxAGptWlrDSYJZkCSiJoRZvCgGxHGED7B56GPbsVw
qb2qqDXYniLAPKP78P+ib42ZgOA4Vg9rHAOI5ULPO9Mnq/PqU4T68n3162cTQIQHYzFGmSVaxh+C
glUOFobD60GaXDpKUhnazPOcSO4t5lDOKThdARBuB94sZKC2iIT4kpF79LRUbu2aEw+PD79DkCAM
Ec1N1/ju7PbW9CtvJgcFmQm3jTlD7XlRn0iSTcQ57vJWSD/V4nejaF2ae6up+Sz+M3TbKLfjwdWi
UQi7gDol1skSovBgSCBK95CpRmTDnPngeGedcASe47HRUvO6wNzVo4fA3ayGURAhxTkwLBOZGwrj
shP5AOMFtojth7a4orgTCMpqgTBrlS4vtBBOLgm7ir3Jaeb7Kf4/pIlJOckfmgKpk3/L65Q2DzKB
bUVGJtzOeptMBpdHE8ypYSfOrOfdLwUh2wYdRN4wH43tYe/gPPu94IWEu4b8O+H4Iba1mTaHkAx4
58Gs4YLKm1YxMLbvWY6vgtRmMwPF1ig+SYTTC9fFw3bFJhg1y+Vo+Uh2e80Icpao69meLhwM/cYg
BETbDTASivb7MADr3ynowfL8tuoe7lHnqjPC9q7HeN/3TZxdYf/+9T9cx2fMGPic6T5gUALz6BNl
A3RQd6ELo1OYIZNBTr1D6qN4BuplN3IWYrxmu9o46dU6P2gwFb3GTHzyTEtO0hW3zc134CAUB3/j
kJoM2YMbZbOXrfXk6pEYzYj2xcmag+1amVsaetwTDM7P2KUQtvEImSDsrRODC7jhn/tiudJWeI9l
toNiy4CFbiiQ6CvB2X65njMI4EdMH3NWodGEGo0NSeVsPNJ6RvZVpbTNWLhPejfruEAJTqrF31YG
uNOX9tCv3uYWocunHIjzy7SkssyZHF36PRNWdCnAT76SaOlNK7B6oqV8zbJINlHItDMilQLFRLI9
/d7g4ZbD28CfPQu3uxokUtPwPbFEmBci1u9xXg+ECGoKRyuRUIM4iNpIGBVqk6rVXsgg92lM20TK
VaJC5tKlTsq7qubpF0JKLQMaF8FCuVERaCsdxLCNmG3dvH87MCv/kCrTJM3HkS5uUb3NKaCFy/q0
kPomkeBn4U1d16vW/MGBEHOKvp2f++XSnSZTkyO2a8pHyMJ+KZWvM5qVqNYO3fqHRvhFILPgV42a
Fcl9JTSBaAI0VgioOt2bGoGpFPcUvl7HH7ju+tZBM/7QuMIuXH7b7tJfnzif0vt4WGxpG08TVbaB
/6vGnGxrUsdPCLggxXlx+cX/KvrRr/QZKLdB2IRoU+XIlTxcuVljv3hXvTAflFlPhaKmcoHMERtx
OwVl3TXrptmPRQEijoRFkB0fhZ5toACSk/ZEMd5wgGkjsXHtzF8Ad3rPmFNvSgCo9jV+rcJmTKsI
HOLJLXJx9kdyj8Kq7JBGo7PGjHbj04lzmRyLdUKm3ADaCaJbK2RgrakOuhWOTQ/poxGUHA1dNc/n
fvvL3b4FyAISSj9m0YWswW1oK4MUw3uVfp0P6bPcRZyNfb6RWDuYsdKxIB8wtSi4kSa6bn8Cntaz
kdcMf6uj8d2fMc78CRw/OXHVQvYdOf9MAC/WtZJC3kAYAXMvtoQZAr5BUxiR0FrWMPKMaXMp0sEr
N3KqSrLRyPDt+tT42n2chqax9DL/2JGcoXBlTZ32lfVHWO9itP6O/x0WU9AVkiTJPrIqWsS/EGmt
xRqwoN0KMH+A0JuAi+U4msU91ne7GixwF4RoJzWj+htWtAxUnA3T+x+/YPjg87QXiFPi21GshQp4
KKLCasB7KjyCMqBShbWIKvFJfnVo1OToNfDh6f5RVi7Lh8bwcw6hAsti8RUbyi6O+dEDnR8kljf4
OHGW8jkHYfzpq452XKUwkE4zD1mdWB0TavyjkuG8LAjB8HW27S3hSqozFiTLeVG7KEZFReMBgtBr
ZAoGhylG3IHTxQTSFhdT7GsNGpTB4zc3STPFEAmzi8TYtqsIN3IIHpzfAMul4L/fkL8ecUU6Yfi8
V0d2exTNLxyZ/GVvJUG8s8IWGITxzBqolI9iAnmGQB6V7xGue8FBmHhwINMgJTIcrWmkr2oqpqqJ
U3ZRS17JnRihPP08aGXtDih9rf2EaRKO3puLBKChEubMDkReCxPD8vew6NuvV5TZGI7SGdDbXsv2
nfq4WHaXRV3IPWaIEVW1VCpSmK8ndsi7AbKR2UfnwzgGyH7ha2cZnhBcm8/CMHX+QQzGABOekgRz
nVE61DOyUL0bUwT01DMU7sXzM8hcGcvEyt/kAX3pfG2cG8CGL5WYL96GRiim7i96SZGHyzgmlrT1
3gr12kCNIv9iZThH7eiT5suxDYQED7SdFZWowNFVr+hY3Y64ye9iIw+vaxGz4W3IL1g9pqKRVOnm
dOV+fQUHk3PY6/n0CRRx9DwmM6nltfvpIhpmYYCoP/g+xpRZtNT7uxM+yc0UxqCnikkol8Y3R3Bl
Ncl+iULAZsyTxCFcuIlTLD3Fj1uj5U7UTQyLS3pL1Pvs8yuD58c4hP9eu8ij4tfaTDKm/HcKNBpq
3jTrQmt7qkd6AoUVEcwmc4OVg9IKq9dpCt/Do1eyDINuAzqEgLt6JK6kYvKIkxoyqbxkquNyVBzI
0bND4nD3UzyvqNSesxzJ+i7C3lpaXDPZLTQS675ZLZsOAMmumYf2yCy0cQmuZHKy34WREcITVw1T
RbESXW7En4NBxrmU1+y6wV6dLIHAksB1l4WLG7JfmNZ8JoMYHMJCjYnbEQjIuleOwoxk/5M/G/aK
szga74NbZI8B7Y3nZsLSLtpoNDOdEE+lV+PrFLlYh+ip40aJ3jHygEeGYTYfpuN4lzMETu85tSrd
zspV4P9lHav0iQZM2mTmL8Z5JwRdZrjCix7mXw8cxPJkYTSQDgypAd6MNm/3IDvuSWVA13y4BGrh
qaFH/mihiq8L0twiG0NTiT8cdvYHl45/Mebfz0pyB9NVpeoq8XD+bpSDcymelowDJxGT1kTYNIgy
Wcf87ASEzRo7T3sS88E7sIgmnBcYkS4tGHmllcjTOj/HQhk7Ys3sjmDShjDGOURlL0Se5/k7VKQA
wgNK9v918U3XAl77PvX6rOcZBPBOPxSHqcnX1ddj9X38bNT3S7A72Xza5XF7Vvcq2w+iaH2diTuI
kWVD6WDsx2DPQDPcXgrUQUL01IJpPLNKe1DL2lCgChfT3mFFMM0l/7FFdtlBjBz5jCcgqwn+HVng
W77CXCeK7rz4NYK9ODyrWgaTXPjkZ73JvpCKqGesz3dtiG9prF41lrEGN8q68SZDk/K+ZUBy15ja
MglNlrH1HHB9P9K/QR4Zc0SarMUbZL87jhQOLMntKaBg1F5fBM1Ja+EmXNiVFpgYwXlUUWeaAiHf
fQJhs8ATsD/NgmdVWlqJWhF/kHxumD8kzhrpdycIqJ0vqVDvoiy8r+GsNqDBL/9e/KIyjdx5w2Yr
XP4dVkRApdAwyuxHEzZG1myyuQ5OVNXPzOl0Qnv7C3DmWwNAEWlGLXZd7Kprw1oYAljzDqHDWklv
zlsA6cNUTLhmvcSuaPNZEua2HluWxTUXVG9Ac+giMYdqWPdXtCMWUnM8DQ0OdfBbaqnI3DXyPNw0
jUfVgHRYwD71GsPd4Kj+iyA08OtDL7972FK6Xb1wo28xiWvIuGgeaaQ8qjGa6rIfAqANNBLlVqOq
jcg497DKNSpg21HDEtlYRn0ZJABCa2gCOFGiEglTBMlB4iLo04hx+aoOKoZfEeCRVxj77jpPxAT2
j584g5mwbS7h/tpX81C4gFN1xwg050QdYunbWg0O7vFLdsPpo3OKX20YQpff8r+SakjwSmMQwYQA
RTSAGwSZrVzpuXNrcBWxkPv9yGTG4ccLp6/qo9GQ7QodMBQ7A5l2cSuA+P3J07zNgiFfGYon2syO
exzGKonM9GFJ9h58FJcPzAQX4OGSq251f+L2tgwcYI9f2eAGajmcWjId/FLGZndlI4/6bQahplzB
iWfAz/Ntb9MH9FilXUKPlLsiDTPcYwFS4gd//Fyudxipq7ZpNjRV4+iVOKO73CPXDc/nkzN5jXkc
gi/mSTiA/v5OQJSJOOEqFReE7gNeY4HfVZN4EAprouXr62ydOajg4enH2pbFjcKgGD83d7QetqC+
k7tVQYBBpoW+NqMDXLF/ngPQtBi40AvfJWsh2Kp7Bg1p28tsO4s38xysCWffO3e19EYAvNLpfufw
ogNnQqQ+DH9C0RGAHoscYruvf85putipij+3OVtpgBLCphwTplMZyX4b9TpiJC6otWeF1gDm28NR
DKeub/1YoMfV1tWlTQ35xvHlt6fD6nzeUEiRdcybQSxgX+CVorHEZIUoARcohqrbg5TboRG+K9v/
79ZOrDPR9XyiTPQoR/ERYCFR1VWgifIKwxutHOGE2I2mNTte1YULfAXrElyfxWHpsmFHcp4+lI+i
knlE//BHq/nio1PjPI4lN3qK+jgohQCub4FpCazT/YMRamRT9Sku24mFCpJ8jpVUs6IZLUhICwu/
vlzsTIY8RXxS6GEwmhIV9jeLc2oXtwUsdQAQG4ycNPtg4THdiMQ6vBvfYeVhLwElZlPhkxNKPxAB
uBMtr3XSsg6oI958SMAVe5/LYuZsj8dp4ou8elYgqS29CjVnIayxVX10Vq/rsBDk9K2pdLzl3GiK
13sEzWtVaKlUMKMMdL1KKXm5EpEUSRHuKVfBBpgIh8kTdc/Rd0Rz6XYfZljnJ7M/agtWe8nd3GVF
St1wSAD93BwWvV6bRtQKYuoJYJdgJEQHH6kfLFnH5Ih5Hij1cffAtj4Bd22pRPmsNZG61mh8BWrD
1CNhYlvRXy4aOwcKRVaGd6Kvj+NF49OEpnTY8TUYmiRiY6Yldp7QdcJb+uDOpXGcKuktvljEooD5
0qOgDke+VcqPRpouuxbWysiJiLNzkek6XfVcp7pLAjxDCFnukRf3yuGQjXPlInKl2yPDmwLu0of6
MTmnzNaCjZAgHQJt669g8Xjw7hSoVfuzAIEPHfVnpcuBhNHj7k7oV5WiQCtp/PICz4qx61pbh1dL
9tVaAPJXRZfiOCDpeeVmSC8M/CMwAXgv6kMxgwIgqsUmDUvYe7pWhW4fF9Rat37uCbLiUoZMjOfU
jHE7AXxfJoQ8KR8f5yaYCNyaESwPKf5sR10/vLOwK2u1bMENvj0HkV/DD/RMF1THOHJjEM5QcTmI
9lm6CnDs9lVpQwUicjFs6kobNQFDsm6EWZR4Wbu1qbA9JucylVVVKVaX0KVQXCksSwE8qTGgpDwe
14PDZLhha5Z7PNIpn+14oaSV8Fhv+lxLYcMOrewBvdjO7CzHqPYFhP7gGKnH+dPSsqvJBxRCHWEc
vVq8G0qaEiQb/x5w0SW7uqMS1osXCHLMX726v3o4ZDhvf023CUYOeV1EfH84+IS1a5EXVfZC3O+7
08TmZ+RIp9WaZp3vUEFeRA4gRbhiPi1ZBpVc63YNVPzPeAJVEzhsONELMJW7xN5vRL/wu2q4d61a
WqsXwHiCBy8PY5Lqt/qH9G03qNL2jzYrEsq99t0bMvoxtpubUG6W/BUmuJNtXSg16aTR16httFd5
FoqtgZjHVcWzubJwXBUInfm28wI+YTJsx9hd22V0SwJkPtg2MgALq8rplSb0kzp1o7no6J/wO5z5
ITCV35DN94pAuoVY5/QjX3wI4NqbGRijNuWoVOrwqa3eYJFUqHqaelkNyyQbFIqWAyYbg9nIjR6y
9K6I+RaJb1VNRrIhY7jmG/Sy8v0hLv4jX/2RH0AseBiSSTrcAn+ddMBba3SKshmqabiQPxpgSt/O
txcItWo8/g3aSDdyZFqo+ZRW7eQ5VEUr8gbPDtPG3CfdHsZzMTRtkL7AcYao5HNA6G7dANmygelq
dkKeQ+DEdVTZAsRJqXgtB9foCn3jZrBE1lUeYSFv5/3fXk6UwfBhDlBMUx2A3MeM2XKT6QoUWLM5
GAzsVGecrQDjkVaR1GwQrFApX0OJVYdM1QYT0qjd+n9byEm0xn/Q8/xBXJ/iiaHXdjcfhQ/bpevP
GUBe2xSvniFIW3+xCN5j1K3fHhmxkEOSTxZ09Mlrll5dFIutrL78PUMe4oX2FvHPhmugramQwaDc
WlyI3WIo7oY7Qk4sDxh1jzbjr4hDYFU5hyIHQtIn+VTeCh8NoKVD5cY0HjZjr+XcxPLMiiDFa9ly
766t+WhekSnfzh2HSclAdfJVvvRBs3C+kSWo8n+qwbEYjFrfSeF2xx1PD6wSGy1XSihVE0XG0u/L
+KM5pJQm9O1XKqyEROSHvJ22bydT4KSOZ2fDjAaijgqolmZI2kCXpQCX5ReZ0WZuZf83BJrbJvB8
YJFY6Ukwwr4Epdq4s/K2U7/p1qR+0xax1trFtcJzU6i9uHEq1S+Vwpo1FMrsrgLG+PSsArtHLBP/
nHX/WvtqgAMe0bIaa8sG0n1TcPewFYfma9QsjJnWrGLkNyMArdKkKttqO8jXUPJ6j1NUZUpZxXqC
tJVo9E5Y+B30l8OCf2cOeZ17R8D1EovtM54x2K5clF542ZXAtgJ6cS7tVZFddXc6/WQBbpm1isml
RBljHTMrotBBAwLHuinyTY3LMXntaeDZB24giB8N0ynTsotoFFvyW2SQoIULr0Xg1c1jMNV0AqGH
nPhHEtKYV3vW+GNoaDIgameJTzJmUcUIzyXwXlOkJT+olMpVbW9OpMySM9QoTU05vQ/tQoyNMKZe
6oGpYrlRqhtNMl4ikxCTt/YSchJGGK5PciGdqFbFHQuFnm10AQr6qiJZ0O0ijXg/NwauxeH/5C4f
cq49KzbXgooZdozBE5hU/ryKCXX+oYiGxFz7OvXg3AB3gOyfb9scNxntsQiWkXnLXPfai5P+A79n
en1XjFsJHO6TsOA3xsmbAc2tBI2olWaj/D2lU++EBEwt3/I7NIZ47zaWtIVtcVrgZBSOPmGAVt2a
L5G7SQrAyYQ9oaEJAeWVbNF9rBpZVsFALAcxbS0TMCrLe88wSVDOs+0BAB5wn1NqsOK3J0lR8cNE
srvirGs4ZkM7l7+YeE/gQ34gvz7jZVw+s2JcBisatbNLnBOkdryDeNGo2uTcKBDVWQCorMhAaMvy
rFPjNpPG/Sur4cxJc1hhr/xEGgxsnfXLbHmeubojwe7407AvMGoDolqM8z4H8x1YmYJeEol1EK0t
MWSc35YPnV0ht87hRL8giJfgd3zbLAU1WZa/IFX4st+uSAmQ/v3i2l6mBlQlnUJ5o9PBrfNjv343
WtHRkk1I41lhVfGSaEnzw4SSlVvlaKBZSvsuOwXZ3Kpo/W3RTh+lGhV40KY1s7WIc8LTmXfOVld6
fBZN8mf2biGQCgG2jgqgGbOqiC6oCi7OUmwV34pzqUe26YfK8SitEJhZpZ4hzr4cbcIVAnz2Howj
IEkMW6Jc1pbF37zjA++wv4eNhpYEF2DkWzrsEe2K9Bn/+zhH1r61gZ3H28VCR0o7i+jSp4RxMF2F
u8eXiKpx0ul0jwlWZI/xhyWPPyHrUfUsFI1baN92PxV6mq8LEQmbBxst3qANH8umNm2KcxE3xYW8
bEGN1QBe3e56/NhM+dMomlZBCBRdgQUx5i0Ucz+4uwoYX4+u41KrTpYimHd9zoPqUCEcyGWBmyJM
kpV4ZYw4L/Nj9wQWtlsO84tKxmihF3w1Q04yoGv5iHZ/4c+U6S7u3BARNSOdgYUfRSDqW4OX1ztq
HkV3F2kCiDtLOixCvghtjAjdaBjuwpmWwg+Hvq+S1gx64/L324H5z+1il6quXVHFCiBSmQs/M3r0
VIwJ/VOG4l6LUdbtMXlElGrfdaxwdSbEIQLXhVa+nWnm4bvCuhhvMvQUuk9nV3bbw7R16p/3KRKP
YxHiDRkYGGvNeM2/gp+niq/rMUsD12Ns42aVM1BQ0VV/86vU0OOhsv9aB8ktm8Zlqo/g+khV4ySr
6J5VKFHrGfcC+ovb24nScKhjJ19e1MTNtm8HU/i7YvyFtR5/fxCEF+CYAVQfcEeCb2GAh7DSg6/P
mHGArUnKYuszxldzj3cBfMx37wVz4Ctj8cxsPXzV/HfUtCSzo311wvDz2KGjjfpixRtfNd4M1Vbb
B4ROmwOJS5N22aSvv37HNsrFGRB7as3io5/gG4zx1jVc5PPpfZTGHe+zRDw0uS8iQkjynAo5UNrr
xz7fRC5Byi9zSL+1SwUalee3H+F/bhkVJl4Xj7KaOLLwjaqNSnSOQ7OUxt5jpq7MzwXQCHS2qjkb
+lWBOjUzaPUSaU71kbcwb+NQZTEiibW2lZnlA7vXZsgPW2eEOGW4VrH/F6hGLmVHUWAhHUOWQvqq
6/vJ98JUbVJO48Z1/paOsRbr0ZzmHFmp7/HYfzSfqDrqQBSGnY8BAeM7mcHhCO8NDMA2VC77awof
uor0f2y/uVnjhHv5lNpJ2spjhvg2j51vSjtOGoZfAStxd/fgDHyDxL+4CrXx3Ip5J6E40jwNNX9t
CMCA+40PZafBA6gjQCBeK1ogrrIOWTsUmfmySeMfBSsaA6ntZ5jEGviWuB4x29S6KBBlzWmaIb+f
AIqO4e/b317BGblAQ3ViHXf09GKUtY5zNLFGxxy4I8foa8TWJf0TrvrBm2hq2FXTmjSC8RsU4Som
oy16A776SqkIOGEC8uNdvs6vRAjy6/qpA7vDtdsC3ipI9mEwpgGaOcgNos6AfaTgdKsD1u6v25sk
cQHME8JC2V8xoj/K6pXSwLh+h7K41sO4sGd183eohAZbm4lav0GvM3joknjQGP4jTM7zjXPHFn/u
3amZK/lyO4OK8HZvMAekIE96SWmEKxVkpnawx9J9GM2tL/h+RxnBTNep3+eRP5oNtcLeeiatgux6
G6rSp0UMAocg52BUdjIg7V05ivuSOzsBCaSwYhvAidzgZtDbKzvgGnL/kgYX973z4qAenKVeKxCJ
RDbAAPfB+2tbwWe5bE+o16TtNaQR9C8ldU0d0EjvFGsGimU4dTWQM0n0dSofnwjBx0gte/Bje7jr
9YMs1SXbpS3LuamNVoOSVpO6MCQ9bmLAVGDyXKDmRZytLCCXveeQXhEqza+3rBnk3734auCpyUbh
qyLEqPrqxZSej02TJIdmTf6Iy6LnsL3BPrw4X+7sPr3kEuBGi4PbgvoW5rtOhX6pecl6cedYl/Sj
G2ypHmqd9wDT6v7i6/C9PzpfTda4wwIK596p0seN9umlu9diit9cHmzo21hKSF6zQK9KnR1VAOmW
njaLHpEyCRXwHPLe04F8eQxp/m2w/RnnC5FSU3Hb1PBC4kRFzgKrjYXNky2yVaMSC2i0+zi0CfYu
p3xasc2Ff2Zd0AudgsCWY5YxDEqeKWobiNM5nosNs8AGJpKnYGxtyQa0e93DK2IBn/+w4YvOYIsh
C+FBKrJmeH5OwexheVJT+himhQ3CqVO6yA6tYsOjbt7b98toaEEUCoRjZaqGvWexxXltzjO9X7YC
681FqZl/2ZfhOjkckn7kN1YroNs7trjInNIJB59bqvapTY+fZ7JKsp+1BRmQ9dle0k1Nwcy5kYJ+
vrR9Pj4jgJv+aFWWkxCdIrmFLkIwglOx9CS7VUX3k2B2OhD051B3oumbGih+44rcQZRW3ZauEAyb
B6fm8fsI7SY2JDkvCh6leuBl2MXd61g8E0tHW//Q0jBU5ozDZBAAjvaD38iu/U9fuPraTPIrOR7F
lUdQBtvkwhZenDBwxR1xcXM4ucxj8IMtOE9sZkFtjwsGimRnVezEGjWxTwqtltnS9Op8iCZsTw3Y
GwbKrYvKR2Ar2YRv65rXFGR/mBzYxyj9nFVLLv7abf4pyXujUt+lFVbLsWN8na0SWkdbPysYz0b8
M4eBk7P/C/kHEUpmRtPew6pw37rom8K5xMSDbpMI7LLzjXUwLn/AO3b1ghEKw3g5gUKi6mmi7MMP
r2vhVSKV3Em5rLIPqSz93DVaeBbXcHBppW8EKUge9HmMdiq5r76j0QlhyeuCO0qEVimItYtY+qEF
b4hAGIL1TNlY0Db7AvpTcxWhP7FcWPscdcTf5yDHjUMRlzs7E2giUBy5anWwUnJz44PDlxnCR6gh
Qq7W56HSOdalKRUb7522ZKHJdl2aPcyhWtoKsRoDaR6608ZA3dwt8ADMrZxGvgBGQgR6KQuxNf07
4HOq9Dqj27JExSVZYix/PJgq1xGMKkjpj5EzRgPjJnENLNQea+5xNMqUkWS/kSnn6ZkLT9h2/agf
2Olkfb/Y53h8/jQ9xkPMWXUAOnuitHdoJbO1sq0muE3AeDtOHTgxy3E+aOl6ywsB8otdeMBJEvU8
niYwWXy9TvILTAB938b0DwNoi3QrdLVqyrz2Nt/u1zI3gO5JaINZ270zuGUeh4XCRRU1Gbkk5eZM
qikmoUy37pKlXZHWfx5vswBaze+XqCRTAdHth7FU/KgxR512Tc6CfeCynaOaoPoNAqUwvp5wa13R
jMHMpdR6T2OVhI46pGjhXUrbASThBnA0FG7QtQKEUiYQwB0wgAg4pDSQdO8BwmIV6wO7m5ygWtrI
5hS76O1mv6+QavhReIlAtNd/cNviMCZ7rhirLEAuJ1l621CRWsTpkzk0saf/+az0DLkSutf3XaBC
xgrL+tWDBmYtYQf1GNH/h5xd51Ht8oG4hk1oQ9mphMBbXwsYWeSHNytI4QWoer4puFZThM34miaY
vHlhvNT114/Ebf9YqAtlGCCJiXfdS1CViBN4kYhZLzCJjEbwiBR9sQTSgLE3g+VIxN2mP6194ARA
4/xFLfEDI1rxxMJuQyhSQKbsKqEaOcqSeCq9WZtGb71L3ArpLyPbBmaEecaw3wr4tBBYN7avxGcq
aJQobhyNSnpSoCs4TTLmsyAJhnE1HOdZ6PfVm+FK3BVHUu2Hkfji2fcTE7KJJXTN65e17vFySYeK
VhJqOnFXjJN+dzbumSv2YKv5tFU/B/EVdEf4h5LjFaeQ+i/sMk/M6PcCK2I4fuYcudGzIBKW/WxW
HQ9jzws2aLe039sNFFfvsruTKDP8Weei1OJrk9Zg6dLpSI59nVxMccdRZrMFpcIlvV9P3acepMIh
7nrJikJQfqwvx5mtklUrYJyFE7mJR+wBWGz5Lz6nPxtXZmXJQsiPm64oR6BBaHvdkTelE4yMOLjN
UHzFHxVhlsUFtwD5YYjwmkR2VYSB2RKc1mvcwxCs9KvtpXYjTlhPxYP47JYFPs284zx8vsFTn8Ct
6iRs8YiqIvBj1kWS+uRqIAWOZH2WIN/go2iJmNBPPJoaMCcI6ei5dSxwoC4o8ez4/fx0Wnpbjftw
svGWKRixD+FBTpS8ROj4heTlVFLr7QaEIZm+TKEQfvk0ok4l86XrwQsS8Y0meNBUAj+vBMGyV+JC
Ynmb1VB5RD5GL4oo24weap2knaH+TYKLFPnHlvODw95EkuZuSz4kjb8mPIJRccKPoLJPlVE9CPFi
GGa0G8q4/qJwZ0PGqWf3zUwE8wr3FmI2pH7WP9Hm3/2edkfT2BN/ifcoy3gXArNKngPd7MfTjaQY
5XgqDuIqhX7eBu0/lWpOBen2ebbjZs8Y7wsu9pqq2hYp9FYXRlh/M+Lo2rUfB3XmhA9tJR22DcNF
grv8Z/uYw4twDoGmmIfP9gHp+kQ/sJv/S8QHWgVktJjbhQuEKcjxX2jvdyh1TK4UNY8U88CDhm23
ibsMx9iRTYSULw0dp28RJF493y9u1evlf1Hs+uIqWueLsWvbuMtV2FQ9/37C7G356/Hp5ptxZwpo
N7sPvo6w+Sno6yBxxXnNhoKe6yfqXTMbZXJyfC4o3fRn7hrFdwNpnApmpZkX1yroXJZEd+f+56nl
10G2bMbN56XMZwrnTqZPC+fLqKeiu0Wk0Y2Xs/ZBYNx6E0N2te+Cmgyod2vw4qP+UWPxQ9LpAFLS
Edt9XkPsZGLD9WtDSWwZ2Oo5w12VMJ3nsLSQIlP87n4QognbelzuDmyBmINQCRNY/C9/Jq3paQqD
DMlWjZiVun7Ygo6JjIhcQgDSq0Jc90W3zIgKwTllydQcyUJp6X+x/ka46D/miBjWN8HTH731sUE3
cCa09TRQ3bmx7yYDq5yTz9ATEPKd+1adKMCRuRXAfd9nUUXZyuXq8dgcKtKXYNY2WDdtz7zMLLHs
EnBtNcZ6oyQ1GoB+iC4t1n5vFU7Jn39MjMxuKRIUmnwBU0O2CGvGACl1veMJ3nGrHpOHB1wxTSIj
ZfX/rTQtK5Y06mrqFbwUFAm0E7U+I3nnehyjW3P30TsM9yh6PkMqyrtTvMFXAOEpQcGcgzyPzoDq
uySnSVShw+YaPIXAKDlVcKgS+SMmybhayjXctfJ+uCg0EfYmAGrWr11RyScq6nx819OYcWDNRqBT
POzoxtA5Ftxfsd9FzV82ur/UqclJb+rpL/CYfoaR9JFB29ZvxiU+BlY8sZvgArrkFC4XLFVrzNrm
sTv0FRCbcQsoidl+g+kc6YZoEw8mf2W9K/hSw7qqmkRcl6RlYIkS67JJGM66BnHW49RJqTna3vio
HcO/0ZM5hHltblgpVuX7ZaRbkDR+zpUjhOQCaIV/mdxiGxDBRC15HEgnX/zLArzZJP3RzbRe/prl
2uAo9EN0esJzAYNMXj+ysooTajtc7izbsVzUANNyAdUvjgTjrAoRglVXDxYJ12z37/329S28bJYk
Ny6u6CMUh/qDfJ1Py8GEmqr6S32T0aHFSCKZ+8jrrNd7nKxQUBDVLc3z5UX+9OTwVWmsZmPqgGyT
kLdNstRmhyXufX7h4vp82+QJibPdcajawwMwPTvTpDcAouB7HXxh17c9o/z/h8Y3R/HQyDYUT468
c+u5WO29JOphPuTpyC+58a6q/xsOkAjCC9A83nsCW6yYkJ2Nee0+EtKK0Pk7OFsmrsk5pZBbGzRo
oIxdlDHyrMBo5P+ju6HZ3v+oOHWlW4EHG3AfrWj2pasUP7Bw+2SdujRrWvCpok0Wm2AKUl8oQPsf
vaNW+hGXVhd8F6CqdGRgX5/eQZRUBzvy0Xhfv71iiwLvJTkwGxYnByKXIxlTKHWcSHWWpGvm4FTA
WLR/D9YR8KpMalaeBZcZU9RXbz0JxMOYKrHF4RPH8ibWN8eIyfC6hwysOuVfdx07Uo7akcAITB0g
I8UghwaGrx3D7W8IbQFaMQrmRyYYmadI8/xuKORQ7tSENPucIU6wI/yh2YVegl/wBEL2petJ5Wd/
ctANnAaVrxW+U9MCZi0BopS3x1zjRviT2ytxKIqaWCUqlLryZ5hI/Qc5Hz/FHETscVyX9P8Cl33v
1Jcc5s27A713h5ZtFql+G9ST7udTakBy7/q32mSCX5p/EFaeAoiDipSwzJOsPrJV25sJbG9gPWSs
QGURZXVeNejcK2/P191v1YL9yAHs2RSTHTFkFfvqHuC0cNkb7VBZiUpCxz95bjgUnLwupgJfNG9o
xGByeWEM9VJwMXMB+TrxdoIf1EQ2dA87AvUkxARox6gandi9OVrGDrMa/NWWymIdR7BXM/SHwX4h
c+WoNmjCUxNLi5xokKY5DoSo5Zb77XwpbjtRjU7GifHFJJb6aCw5/5ISJAOuZcZy9JoB4GOUgKbZ
NlDabmOzXf71WAaNumAUcFQZjbY+7cBCSEy6JbU8JhcfpU9oYVgaDYKwvYX+VHWSGf9rhiDxoKbH
uX9tWOz/13AHX8ks1qgtXpahPfUmtP7LHloHbdRHI7hfMnAlY6XP9klm+kjjWDyEBIW+z0voT4s7
haqkXeh9UtYcGm7uKEImjYFFa+AbJG8Ll9MVblHu1f4kzTcBRJjcrYLyPSdVlGarO6EMziG8076X
KdYK7+44emLX1JScQGVmgY9BZozDnfPz/2olWIcN+3vzL8VINNEXH6TpD0DB839IhA0ZP494ffxw
dv2dvh7TN8lAFHro5wG5cGQ9rO9X1oKxo4wI0sfItqa0WaIbbMR0qtQxTztUV1eUhjS9qPFcMDT4
Vw1I2AxEFLzkINl3uYi76Bdgh4HIxyvag61C0/vNboUGD1NkKeqyWP3fdHGksISPTNayS+emuQuf
ESoQcuQvm8z47y2MZnnDWJ9Fl6oFjjm5pesZlQnWh0vgXavkoDJafGB3iqV5ZezQnJpaBT5OPrdW
3oTg4I4fFFQZu7vUjJmNnd6u0K2Wu6E3V3afuSHRdpugWL87IhkrrWWTD4KgUaSgdBIwqffxnaTP
33u1i1Doz+8189ECB3P4GwRB6ifmBpd6lktgvRfd8P8x7wiInRKLHY+7T4knxMhL1QJamKd0POm5
Ur1r8NLWmYyUqQYEchE5oRBIEVp36eCPSl5BtGUr2t1QrqEmFZoLRQa1UfKxqh8YdD81Mq9NNPZB
eZXJSGjbmGEVisZr6gBRA+AEICb7K2E5r6W40nPr25sovUO8n9UjNJXDJl9UzrEwzsyhD2D5ynnD
ST5w5WcbysvuNlhqxtrsHGm/DFywC/Vppjm1X6gmUWQO9rUi9uBK7Xf1ZZXqIVbPWECm3hHs2AxG
QT7+E5xleqRi/NuDfuiLark3vFdwVYFaM+mZbcem/sQhOrjuUhyUkmedqqkx7lVlRADRRmbz/tEo
PXRSl4MaBjUs8AGXt1S/PIVfx70RZP2QU+Y7CpRieE29jRtDd/MBRouBMRMsK5LoZj8HlEZ1efyr
lcM1OWXHD9S/9skCUqrVYTq4Z4SavzYoEATNQWtH900uyNw2EJ/LSK4tdxdsfwTN9Db7PtRmUHsX
ql64aokpfngy+LjsfefuyNj1TBGDs/jgj2/WETRQ6cS1Lq2yBTovfNEmC237mJI25LxrB9AxuMAG
GyRToDjEdmj8cpr9VvP08MgdgilS8x72XN51eli7yt7AnZ/6HeFJdnksKtRDegJfavMdElWJhpXW
s817xTLG14QbG/9k5rXZzSAg2vMTMgUw7ezMlEvlg48Bm0fFgdh5vNbzdE8bEuuhK+loZ0EY6/7D
Yt8mRla0uQw+sV2nyad9goofgeKkJvRT1LKeGgJKO1AZS6wC9jGugyqRgogyAzJRHq1/lnJTkpah
6DwxHvAkYBVGiYbBGDOMDiqrBlwg9vPwXdx7j+ubbsGFeYHGJ0hYjhHsx0phdwQtCna/BKuxEMv9
h10kfZgg5R5eURlgJ91WI2WWjdQhRNEvkrRvXYxKbj54TE1Xix1gJ7RCS9hsqEHbgrYldTEWkdVg
ncxQWAyuitVlXkxiX4SPBdSP8E6nvWWsdBS0NPYlIfWMzLZWfgaqzpqIdb1b87ZWADB2vqdChqMh
O3ATfWg8IOSJuKrH6xOZnTCKnilHAlKhS4OinAFlo6+Adwyq3+5xiq6YIL6KazTeUU0gtIqR+apY
/iQP2VsaWBaHkW5TGYpeLnQgLX1ILDnVk3J77nzIPEjpNVVRdZ5jd4frLoT7DCxPdFblwsOK/GGO
1GZYFDSFVWmCfX28kQl2gTeLWJ+esgu4W5cxNXDWiGSqNndL8JTf+Ffs7vecgzOeuSWs851weP7/
dnOA+JYt6tOLXKxaISnu8UDiPRZqWJhHRD4SOztMgxz4t9ZpmwfNrhlp7sOjw/jTS6g6/kEE6tkF
M/fOEb7iB35F5XVbtQ3es5CwDE3ASZGjSUcA0z+NJWNSZR/0v7YMlQbbqbvj7s/hyx4hwCtcAyEv
tnAJV11Ldbd8adzH6q8BHsqJm5jb4LO6b5y+DmCRMEmvFLbwg/cXe9aHkrrL4zeSUSRei/n3a4kF
gUlaT+6OmWA4Ajgra/R+TsAIfodbNI+duA1Z/w30Rk76A7sIEPM8iC7E8Q8dhvz2hYdKgs3coLEv
48BUmGJZOI5U5GIz+9Tbdse4XrGl3JHRSYwZBcatCHuBpIH6fQ7NfuDHODbu/rLK13nXbg4NshF3
q2CLOwepxEZZ+qlJGrq+BapDy/Pf+NmE2D9cmCWmANKXXXp77GZjaSkeFDme81g1YG7xh2mm0KkQ
kdl7GTbxNjajnSmsbAAftHkO6sBLrCO3jfBMEQnzhZvSWN1VelbaXWtl7iIQ95ziLkRDNLTat30v
yjvpKO0icR+rD3brom/cv1sqLWvhTpRTaGco+opfhBnPVtjVMVulisKyjL0uIqOoMqr3Aylq+x1y
l6V54pQhdokYtV7NxDkN/bc7jTbQD902rRjEW654otRUUpL4JWLRLyH8pFg9AFHXCrMDr4J/kVs4
/5DJDrJ1uTLK2TXl8GmvX0PDcdxOHuluGs4PPOFh3GCkDKLOChELS3enCZZy2ddGHC6S6qs9XyIb
N6oudUUoywSNvXV8eeK4WQMs3NoX/xpjZEdskd2JVELLurtACoq1XmWW5BXwY+sVuCeNHI0sy3gR
/lPzbg4N0ObRUWdAgHvuj9VTnGR39d/Sj0GVafO8Wle44nTJf2XFohCZvWu3a3cLLZuX39uRvgWO
0L2d3qa0J+uvDefqaJPKEGmNSj4Ri/mWw+KXuUrRX299yRhNdPQf3jzhZiK34Ds2WAhfJ20s7Xl6
5EJggq7rxwcJRZnbcrYb7/Tk7N6s+Cu7fph5VVgrrhECAMcuRhMQCVpAbx4lacbnSrrSSiM1qK1Y
OHOygsQ/LZ6IUADM8m3d3gGJexWI1efJjR2T7vcf54DqvwD0FdURHZ7PG6W8HZzRmaQmwd7xM+is
GfKJlHBcZY5hn3h1n/6yyVqG+yPr/csrLjBHTH9rtco0X5EKjWLadnf3N3BlbfwxdHmSAECZH0Va
STbBSbFLliCIuf4X5RC89z96y+oVaITdwqbg34cVOdAXki/RfdnOG5ehlK5KK08YLpIAjo1N2KN6
lFAw0XvsmFSKRg+mRdi37tUP15M9KuT8p1vvhDwL0+vxDgXZ2mBvzmP/BdXuIEta6FjPc2/gWVcQ
6/JahYNxlxiyqFMfEdfQ5Xw/PYYP8eUUzDad5cIU4fd66t33oBE2kZeJUpJhkqU6CtRZjhzkOguK
eD4pe6Cdk866f4kI9RiCNNzhrMCYOieQxixhAMTQP44JHsg77BXI9IBvJvG/R7iN4LEhQusBwA18
HNa3bRZJSspgliqc+g+q/lePHUDfeirrjuFSffC/yjUPPwSpwtHrN3+2T7u0yGr6egUAXnP8oM05
lWOcSMH0NN6VU6IPdM3EufOumLFxgdKMREjzIg/Gr+KzO65aqeWYBoSBTRXmjEtfBs1RdTVCSk4f
RA9Gw1Gg+UWrKvn1Se0GSL5swIIME/eFGz8ulFND2QMRMR6FDotv79+TTGtkKn61cZ93TzPNmfnq
6bVsT4PqaXeBEUgpYAPWnw5K/dxR88ZNUwU4gW7DfZEs/V6cc2B+il0iTBA6qmiPNxtf2C6BFZXW
us2ZNs/ocA+LWTsulO43ic+WpgbOYeknk4e3Zp7F5BiAQJQFAAt8vevkJwywGifyVIrRPOrPmzRV
e+NhU4/NjMnoFRJH0A9CyFre8YqL6N3d2ipY/lekvETr7I21aDoEcE+73UV2k/Mc7sTAEasN9X15
HRsqoOfrQfB/xIw6MDqeb24hgtKkuaPVPxZ1mvusZIaE2h9RI7cJBxHeQ9Dp8lvKRgsG9PNWKZmL
4p7XRUk47CGaDzWKhppterq6Dvg5MUrt/tbQzQfO+MXOaC36rURb1yBLwxzD3SX3uGll3Hs+/QPZ
ZT0yNDgCK9u4VjiMTSwaHE1tG417YEw+0Indx1VeNyPNag7CJiycZ04Op137vgH8SKELyNpVMa2j
10A90RBEwsB+L1IJop2qElhjmw38526UgNdiN/hQbTy3/OSHO5RWE8hYhcnHexBGrRJGI6BpRHJW
lQsGYmW5Fetn5ewy7AucusEr9Ey7b4L+Qe4kcHuCvG2rsgUkkaD4To9uvyBQM9dMyaja+n3RV3xh
CPfhwIPp/vzIIJTft6KOjeotuxSG73SAzEbe/tsCS23ZykzNB6oX+YQv5kTuwJGwGIf6TEhJcJLJ
czFid14+zstp+geD0nibCtPsaY2aDyGgbpPaHZtRoCXD74rWLexElGg8AX7y3GUfCo0PQLIF0Q+d
EyiQvivDqTd5vQDQTmBAhioImv3ELBL4t/IMZ0OvgphfZbPjOBAdj96VYpWecizAzXsEmAeJUMfa
73wZT4+QJTizW7dGLo7XKEq8ed3j+AaVKbm90TZHvab5jSmMnnypee4SC/P/jr0q7Ykby8QrdKA+
m2THaleYHUSREn1lzUbq/pENRBGgjswnow6tmqKXDNdkKNlt8BgvVXZBV8x/JeAyG0kidocVXRFI
LxlV50f+yaRRVNTkk1hqhWxkE4OL3mgtr4MnLkZ2ANkHeHAyzrvIRWc9R9S2VaNFf4F4u61crf0g
FNMGpYynHftODVt8tPPF19j2hXN+e+eqwyiXIWaktCb5zwLHQvaxqjoARNz4fCa+AtKEN16A5JJj
Jc8aOy8oavJSsdnWDmcRgZWESyVXJGiRI35nQsSYaoEneVOMbvEcOZt8CU3U7hgu27Yol9qCO7Eq
QrnXEq3gSr/evFQZPcAKqqs/jud6BKmmG15VN4sAjUTf63oBuzg3ABvy5F+4jkl8Nq5qzGxmeJMh
pwgsuj5Ng37hB04S/AUDyLzLRb0Ho341JoBC/pv2fO7nO8jXSaALGAP8FBRRnrxhQQ++6vNdEPr7
bW2BUDFmbJiGGEcjqjwOgm2voYCivHIWNYydKqQUek09BEMHfUCJpuNIxPNf70rFiJYJoMxD55cF
AE5T4kNpBwPtw9P6xE7Zrtx2CwAMhXDQnd4IWmd1Hx26IfvCpaIImtLKCbBqPRLPoaHMUWZJVoNW
8KD1TzwNb1w0t1zY3vGqN1vZRHV29LUjdP07yraZF/J9zrSL1fcgguQSn+ryguXSSqs5KYyrBWOl
rhqkTCpPiw3DLf8ZhCW5ro+PInaZXXSd7mj+5j5zfO71Uxzt01lwCr6m/eeXdM895RUPSvpKs2ql
4Hq+1rjczq1Vw+MzXjk5LrMyb+DJxK2Ay/KzCsJuXRGvoSu12H1HynTXm4UArg1w8dxxuOM53tpC
BpKjgovahpCHdvwO78w0MMNx+LvwsLScKM5es7oT0qPP5l1F+1W9SnTHXcYSoTvF1YKzT50tNa2N
aSGz4bHj72tiztfDrfNsR50To5Qbd1jL6+O8NP2BYFo5pN3GDAPSE1Ta7kkHUOKxJ8aS3onNGx7K
knPkGWkSJfInpp6xedguOl3FgUcreZIp/dw880aqWvtU3l1Bu+S43XYS18igNx/zGty2R+vxNtf4
bVGqlvI0omOxvUtP4Z75hEJ6/+Rtv0IwogTNVFyefCobwFOsfWtXwS7LEUweHogT+1L34C2r+JYV
kU7ZxSO8eLqKwbRhTFhFAZgsQ65oA4ES00i5axCJt7DcKcxHF+UmPN4lWeJ70xVXRjpkvBD8MtQc
QJaoTCJ+ULVhl62tPCkr6cHjz5ZukpBsYJtMz7jn+ACWjmagVvzbszAH06gKKkEDvOvim2QraIVM
c9anfpq3fouRwlcvWISTWrSIPsd72PyUaKY4iaJu3q8F2dygg5dZICsZG4AEiSpWXa4OD+Xflwz4
QLzyMgmLZHQyYO4AuiAZjIrfLV3AdOnAjbU9F68ZVRoYFoK3OP5YlCVBxhGrepn7xo6QEC1ZCmjh
Wg2Pyavma8K+iinHofjdo2WVJPXvpKChZGJfadmEM6GnCooYL9EeWrGJi4cLw2jAoc4OkUgUIiTN
1YEuah24kRrmq9q6A+9/oQMqJR/8t5/XuakvPh6v3NiiBD1GVdUNouX5FekwVRzHmQk1EGVd8Lyc
ZGBZcUABJCVuoXAKBFFewSh4uNKgdQU9vTUP0/shdKKz1EnEfSXzFjoTvQQJ5XpHC9jvBRlAgHc4
bTrRW8rsEBxO0vAu2evuXQYtRPHKDITKYrhd1j3VHyP817LUcZ6QiBKF8Ovv9JTPIKsDljBO6iSQ
KKh0+2lwP4nXECPWTVsZX8k1vPjq9Aw15YqfBxcT5J4MtaizOiLCMg0q2vbWLljyid48InTwSr66
p7Ujt4J76tgGXsZR1Tdf6s2VqDn80HSqNuq/9dfCvWT5P05DCC1DfkSRH9dNemapluyuGmlA8SQM
/ZH4fDBU/SKxOS4SWqHLqyPzEhfFukY1XMljuUKkU09OZNXVaazKK6a9IiGSy4kgb2rehX8bY7hI
5CpaWDwFDyhYWLMGvd7dqk/9+Uq12jnej4i/CGWjQP7uS0vo5Hv/Zu1Dr/rAj6wtXzC8goB1/ewp
qyON1lYdpiiN17fVPRXvyUPTT79AWDC1P935jhgc6gbkwer3/iqfRKsrJSWSopMO5NfZX0Sm5yZ/
QFiTKLanDJAEQto/DIAF9IDHTgcSIQ2qDfLBqHgLkGYmkBKsxWy+G+B4adwrKAcbASZ4kYQOyS6D
6WtbwxUcw9XPYG6+1fpyun7wMi/LB4AOrCirUZr5p4JlybTyUjovqL5HpX90pI+YsBFrEOJ8Exg8
L1531AdpuJ9kb3jSUYxNY6OdSkzOnq/bE5VpHP1atasGGpKsoeI/TkFD4ChDOkHkyiBRvQVQXSIR
ui6inj3oXBRx0ZKa5LtxF5AjOHfZbcmM5aLTbZZzXOHUhkceqkgB25v+j1tvxl5FyHg6qUuOZwre
sw/0NbA6NlR0C443qZHGBkwEYegAgmSqCwrqjpGB2yO8/zcbWFMXev0A0CKiXSZmUJ9Hou18wtPq
ZnH+iS7dmPq2QLMRkArUJ2QBBu3g7PUww6ABIfFsiasXcq/kvFqyz+gmOAolxE2CjeAi7M49Ema/
8ciwP/FX09gFq28u4r3N9S4e/cYrQCYEcYAvC7S8wcCBiNpZvqbkzjd4v+GxE/99Mn9VJAClpBVb
dJkySAloc+ojgVGbbjl8cSGBssdCZ+1oOb1u5jjfPrcBZPoz2sz0+sAFkNZknWUiCOFZ0XFp1rQO
RjMwTmkrnDSH3Vw7x9nX1UqVJGb2vPRP2VR+34RbqpMnaBMJm/i8DDEcN3gCiDniuJe8IZBP60Kk
kmUX3YWuPyrKw1p/cHdvsbqvLOWkNcw0lSDJXXd1ycudJD07ZdmU5IJwlO8P/Zw80icKO/J50ito
843+G5zgoYEt6WzA+3m3p6bJNj6reP0UEW02QsyU0ZmW1xTgmwXqLA4bBtzeYiMXp8eYRch9BpE4
rMrGekoMvUS9AEn4bxEER+Nw9ObkbxcS+cTx6wtg+9nRcgpDvJzzRg4aQeXAbqWiAf8neMZovBx5
Myqo/5RtIMl/hFW7aE8IR2SM2hlB8203vga87BwRIdERuNop8Qm4IdvR7kls56LSTZghcSU/hI1W
rHFsEK4zMa8FiaXnuSDuoVYxJjsUoOdHVoZhxLfxh2kwevaX6UO1TXYcppJvpibIvgj9xN00vRwa
NTe/JUxoS9zzpaVX+o0q8W1+UigtdgMVvMupxdRBlICtAPVf+Q7QY/OGGK/W8R/jkPniQssyZvlp
MhzwK1TL1SaxLwLt9BWPTr+XKb/xO7atAaRgU6ozj2tAodQKgqxnD1hBj3Vu9CeC99r6toGi8X9Z
yESRDWDck6Y1QOZzZPQ0Ya2sJG35JmgFQIIcCkmGf0PMDR0rmW6Ong6ameuIQ6SGSaqWtdFSx35h
38HtCAhz3Zi1gMLCWJb7H1AjGQL7Bw6lIwXcI+VzumbSCn+PUkeJ943KIgPaxsaZKVBKH0rp/MkR
rkwype/QMiAECyRQyDbi/Lyp1xYNltdJu6h8gQ/UzK1iRLMD3YQFdhFOi/U1IUYpCI5Vt+Hdn7/h
50Fh4fiH1wHK3SuyXCzr2naFiOhq0elq/zvxhjrAH5vb8Mg0YdCghorCS9fu0yVtdTxcM6mYItGr
gJsWBvBhuwT1TMkkiHFtQMLEm7Id4ndww9gvtrBd4yRIPBKxrLs+50UNKcFPz6G99mT66lWTuDw5
jkdv27AJO3bZVF93TaF6TvxS1kHx/Hnm8mMJkmZTES/P5VDcnREHYDqVTsgYSaySvwIgcUZa5xGP
uldjDtS7dDDhtMRvd1km/qPOiDmZ9EPEvBqExbpMKc9YvY6PU9H+3oDRN5ZetzcPT+HV0jEw6+NZ
prdiLbPXoEa2akQirHxpn4cOjk38n+hg7swhGBDpx+ECS0sl8rWN2UsIINcMx1CP7CSKXOEqUJOG
Narz2kvr41zq1dUrq7sm/kr5P1zGYSxYqt/t6jqm3Ylpe5XyShX+TFPtDxCvALxFsuZ4E6PBZUB6
Zg120GGufA4xSIxyLJociftAsza5Ru+ehD/dgEOfbqSNy75mOxFtHhYZQcP4c8bfF897QIANeWh1
dwA4m1nE6mNN1jjq7BHhYd1aiKvcEQtBxXFjUdqXRezhvBImXZmm28RNTl8vG5v/k+Ad+P7Q8zoY
bway5eOf0MIFZ5WTVRhD4BIitG5XdwdYqdtLk5+3nn9+2YnQsOU76NmdWVQdwgw35gmqrkhwWau8
EVSjs6n2RFf4d4xvegCBACR3R6nYmchSA39psmDM0hlUjjjvsxPnQzokb49QVdP2D4WkYVUr+YdK
2FI60cNw875pyWs1+nMCk0qI11yEDxCRtNeZYs+WFxqZRJ+AQVk6A/sf7kz5LDkfinEqqHOLdV4f
5D+kCKkMGGsauKJ2EFhwSR7jBUklIkfLdCRTI/cvL/Jj12jGwqOtGg+ZaA8615GWyWutAd6X5lH4
bmnq4YEXP9yvwd+bYTozDIad0qGf4TtB50PvBYXhEZMOc1q54YvttiQaxs6Z2JnK+W+ygyvSIsb5
+vQnjcOxC64logg3DbsPPrK5x7JnZEn5YhfzSLwdL8Yf6Tpbh8ltb/S1169/ouFAMVwUc2cKNRnK
LBGv0C2iH4zxtkZ3c+7VB7nwDu4eACUPRiSuaYUl1O+Pym521apVo23oAUPXDmuq4hUfswaE0Ht3
uRedc+ZS/pr4tsqY0omc776ASIzhuDEzFOxJ62zT1xJF46k7mX3h82CHrHH/wxlr+6aC7o8LkEvK
59FvFiTUwYJZptU4IPrTzNOj+z+Nn0U+RuNDOHav8KH2miAtT3YQ1xm2klo4x2uu2FBC2IDBxS/o
ysBxf1e+lPZGRpf5MOEMG3ecMQ9llNS3kgkcetYp8qL3+J9HWIql6OXZLo56ahN3NHwmeqws1Ym6
zbwLMNjRHGlWbqfTAD8Kencn7pcsy34QazIvJp3ZvL13K7ptnPVJUkJksc+xrDgFWuV9ODvYNJoa
0VR/XEqoxYJopjgo3wnlQ+Pg/mmVuv/FvjYeC4Urc0+qjzhRQyOtsjQUAXsGhQmvukJ0PK0Bc2lp
1QWZMpfIzbm5HFsCt5OmI0C7xieVfiQH7LVEnTiuwt2tNDHCt01Esxm2kQB0ctrL3Cw40eJcgq//
vPTuzbAQM2gLOV/f9ABS/o3UnQpLDRkdLMaco5WNdZwYWNgrRVjGClUYGDqZq9irtS6xxFQIOlYp
ETuSS/oVpje+QEBDp6cp6PVHqW777kk/Rg1igUxA3Zo2snuqRFnr3aA+w4o7fXeT8SHtqQBEMuWl
PIKkP6CMgj70+YZFeWk07AK7jr5MBT3pXdLRVvFJa0S1yRKl8Xv63DtMMA9nMPO+RQRdsIu1uJAP
1Ej1KpDXDKfemayOQ0fsUTeMhcgNwHDErUfOW5BASWiqh6UQrGzEQ+Jz902MXGgv7OTRwmfW0sJI
ozodS5loe9hXY2eSgybB7sJdff5qYlSlNKkFzuVqH253N+sUv9fZaVJt+qOMMXhjs6bmJjEAYeD1
FxFNtTJ2XGo9NkFv1zzcATmyqftG/lxVrq2Ztxj3lMMlp5u3z/ucjc32/J1DvixeM3H9T6n9inNZ
rNTy7LzIw1/Rs/oC+lv/NozTMx9HJUmokljjyLSnWcZH3+hxKW+mBCAJHSmmxfk9R10IrXSSaF9v
rC2l4j4hn4m0/gBXhcnlBHu+htJ4MJzyBQe4y31vcNuzUCLzpGVaR/dmObVeiriyHOfnXnN1SyEt
vyWEHRW4DoFnmxExAwxgzGv32Pqrr9kczXL7XOZqhSk3iuwnk/j1GvPfeVbRx+WdIidnL8ITI7yJ
j3i6siZW8SeFUvDfJ2QEVKRgjSh+c6Ia4liaXl4YbKKYca0+hHEMedRAvv3yfGuBnibgq65svw9p
eFtwcOLDwYjzQJjyv74dsZ8xlAbOFm95VbL8n3EYXTWe61urIE1s2itZEtQkBXxFFyD6X34OZ19r
NNlOC+NEobTp5M3Yyiz1Bc5Kb5ii5FuySJP/FB+jgd2l73CGxxLRxxHHFkCNC8FNZIJHLPIOP/jN
Lcyb3ilELIIsjRhZoEWHJt34iDP37xa3Yd/ui32ZSN5qm64g71mc13hw5KYOO1znBvBr4d8PEIiY
HO+maRTEf//O/pyZrW9mLQHW+KVZdRpmOaP/xPrHUG+fTXTIdv7tiFYds/BrqK5sjto3wy5cbE2G
f2v54P08PB+PCgamoYshu33XvkE7IPeajdeC6UwkyiUH8BOqYAVmLkXBg0kuCkSKX2q36dQzPY4V
fNNFQzCb1NAyBfOEgAF9PFGKf8wLGV/TvlvQLBhbRx3Yo/U+olmUohQ0FId/mktUhwh9si+a827E
VAer9A8IW/KZkqtI0MX6JqxOoT2geTJgEpAonoxTHemRiGMARY6876PylWCfQMn6lodGuJiIWrGF
Pje5dlN1//Ajlat2ede9XZMioLWDjaGrKdI6ihzr5GCHjfb+/a4rjfVHR1IT6RqGhD3Xmeir9CHt
DzsyNfEspxyIhyCXQwNtagEyPOuee6o2EvcpDEhLLLXbPL/gI9KKR/tDUzh3MI83umGA04iRXICQ
dB+nWMvjfT3RYl+7S8Pv2vf6sUN9YvlFQmkW+MLwDXMj8MTqZgyAEgZJM3V+tee+98NVuNDkwikx
lBErf0OGXhnAcRyXaORhAZ5P6Zjxyb2VFIU/6ve2KKi6r6aCg597+n4zIbcRLcPMMPDkzjq38uc0
noAlizFDFM8bz+V2g4cmzq1U+4U2WegHWG8NqK2O+FG6sKqKawCbiv89fKUTnJVjbx1q40cCsPsd
+/mZuOa1/uM13Gj1tAKxrnVdVqqo3tpWv/stuzix8ITpdtFah/iYHSxQE13J2K5BLAErPExR8xyw
2C3lO4GNVZEGlxUMPD8+BxpxAy2Z/l/EphXDWrtSijSUUdtk/KM5gKhpfUv4vQ5TzQVH3uRBjbKg
wIRX4uDKDZRvR2YgeUJg98WN52g8WeGJKmGKBbYK1HOBMjDVA6ABhu5e+KYtpDd9Oz6ofFk184kZ
MaHQmAa6swcizDyZ1k4bho1tRyV4+bnVK4NUc7acBjQqSUdjyTSxCTNe6bX8fH2Nt/hgsY+M7QTH
cYaqXCYIE3SKgVS1H2Kw1El0Zqqfx2b6HDGw0WwvxmiTSIJ4zYAo2HNZMbX8TkTU4uwoKPSK/O3E
caoYfJ5OgXHvdW5RCH40NjMTAW3TNRQueAwuBiSNYuM3q2hCn8GSfc5zVR62l2LqR9ApEjy3mdoy
YcX+M+eBDiI2drOJY5ncSjj0yVDS/kEY7xIbUXaGa1SKBpPi2Z7lrOAwGJnF0UGOt6HQPwWmkpxi
MSy2raw0zANf0GVJlKNPD3JAFmjX4ti2yGio9zHhbTNVIMmpkjOqneGA553Z0w54gWBpHchLFu3y
vze5w+pV78P92290x+qUrEpt4v0CF3NBghQt29mU2Hh4r66Q3mX3rrvxvG0/uPAuOzbthVCcgx/r
NdGQeQ1wekZlE/Q2KYx6YCiyXaUseV6jn4KD/n6SMS3Qn7/sqypprj2z5XY48lHZAH8b58/f9Skl
L9WlpBz9W3STU3WVeKOqJQDFCJRDoDMFSPwTWOAyqxQHwpQsgR1WyH37Tts+T9cuzTnYCwRl/+Lt
SU6KaFnfNoA5hsxQgZqm12HRoG/WUdAUNwGFUC5Tfq2Hvd4xKFuPwMvdZHpOoVmtSGX5cgFE0VK5
Yz3kTn7R1dNqFRzmxYDfpr7h2OxStajfC1mBquMKHpGEKkCmL2WxRCbNxFI0rPNtsn0ItIJCfp2d
uhXrCbnZtbP7ujj09MN7PRMrcp7zdRJPUjWPUUAhISu9pcK7knPgTOLzzycwSxUSClSoF9QZs44P
KFcqC8gDsQ1/bsozUWXWiIPyllLykHtNqYJnPzbWnAEc4Hum0pQ0cYhzHfZonk8LXqq01GChp19X
P3d4fUU2Jwkm3y/AQrV3UlQeJBv9CPyag6XKK4k+12ssKDV/z50ljfd9IXcQyaj7QbefZbXoejyD
CuUKOWmP4n4UpqFmZ4as8luVlZkgKeCQ57dwwooutdXkSJwGnoL7vWkq5siRPbo0ZO9brtMlYAeh
yZD/4slWOUSQZCA8Iw+6MAMoijdZ+uldLiEo+1WUOaGLJyGEgTTT0kYZ6u1xz85KhsWXc9X0tigA
Lw2SxsQCKxFQ9M1z+1YlGEB+svklOeBAzqfancw/pUBcTty+NHCVuusILeUvYGnaAS6e4d9RAjOw
dzqiofYJtDt79BZKQpXK2Coy6Sw0pyDGHmVlvPoCZ2rl8UAE9Mh1B/4G2sgTMSAdlNX9hY6oRHBt
0ghpjEFXszebXvQltus4s5/Gu4hjMIv9bXz3+pDVqcF5z5oRU4Pl4ghtaZdYiqGoRIi0kG8IsZi8
Gp0eMVjJr8d3HroAI8oEeFeSVV81dJ4L2XZNmmsjItFc5JNy55ZbQwernYKGJqHF6wttR5natwQf
ucQX2T+OdevTm4zRqVYL5I363ay2XxxE2df5X8o0q9QL/1s23f75sPiYRzRAIxMsLhVwubpPNo2U
o2xWf9n7phh/ydyrXCXF/27wKYof+oNt+RzTNPfjL1ipAmE2boJ7wn9jsQJjgCYsF3srlS8/lsXn
AafdrR4TUHmauHK47MoX2SOnWb2Jhh+KZeZrWOEcOBn8nsSMD6VDsmu3uGZOAHQXk7KgemtOdziS
zNAJzu9u3ay1qE6pw+JLiStTxAeFtY2aXeB61OCHWXXYEvl3xMNyh7zkcP1Noc2D0EqhfIX7i7JY
Pzl/fGArz2otMXEs/dthhqY44aqLA541wkVwu6+85k99z1hfyq70xRA5xDOHgpH+XBjpY6EEUtLi
1ngklHOjleAjiY+sfBT5KJfYngGfvTgBLi4TgTjCDRV/O0Md2uRQOmz5bvpEr7dfGx4LqIhhmpdp
33HdsFDH4sTMuzhmR8IrQZJI3sLEl64EfysAAPqZF2Rtxb+v8efuAvZED7iFoGC8xbY2EBOPOubn
5EkkWzuQuc9wINX53eOwoR6lnFSQDkXSP1rewjTEeZrL5iUKWBO7KC5hVCFcil22aSPm2T2L7UDM
sHn3eykNoATXCN6D5KqxeJOznrK2aSBRSAdV+MHIOHfpHiVuzSBnDY+u32p24AGyPnBF6HWNZ9oE
Cs8fmlmPFFcSCW2a6fWmeu6P2YfcF4yi8pVEigszYX0DMgRv3ZKCw6grxV+Pi1iy2Wd4X7hbWY1p
KiWx9r+0CTJ+rsRAERcXtCrgBFp5YntLzoAd/zhkQHkaKFDV5O4ZYIbrnv+YTzQQo6qeMjZ15khx
w4nDws85JixUEoCcDsDwkymXOxIb660diGJwfAD0pPYBKRWBy34UTHTYcnx3dzod+zDqHot33QHd
sA3aWeUpmXESUKcqb4i65Wu7+Sx7MjfYT5BTRb2T1JbqJ+HYPTbWrF1JRzxZ6gSfMBYxiwiG+OQv
GkgXSZkPetG1vwMDuz1dGyg4PMwwnzVt7G3KonItNqpBUvfCKBepbEdkaR2FyCVSEzVwqECz5st3
yEuETcKunaG1H08jWAxc89/QZrVkEvSMcLHL+YhLHoVDWdLblvwKJUQvtq1Q+3/tsRfN8HGN0ROY
CcgMy5Qxn8Sf0i3ig7ZP3ASzfefrnbBZGe57Nuurr43/YSCbXjMrDzhEnz0+nvy89ZZ3qj8by2Fy
vuAyVEBY+rEvT4t8FXLjtYNyrFfqpyLXskNxuvemkbrY+jf/xhfxgoqLahYjLJO6hPsi8xplYFk/
lCG7mbl9VmvIm/4h6dllQ14VQk42x4ybQVpVk8HFae650quic78Rx3KsaEszSdlAS+OFYFzu2D6u
9gNqt1DRyGT7wfdy1OFBu1eyRUgLd4CAljOrG3F8QXIThL0UQY1psNvEVFKdCEU7LWDx7mqxRGNF
gQTfyN5IQCmLi2bXqR7AmdMZ875Ju3Yyhzsm6BduK9dMpGyUHUTrsXFhCSpCtZCs6ujMXELgDgrn
G405eaYarbLFcixgh/U5/IQBSZaCcypw3dFZA58t5xCCGaeNn7FzPMYkJ9G8K0MM0EnFsZpSCNCD
RBMqcA2PK2OTpOfvM1WF1fkzmgByc9lazweHweTd34WblWo5IRrphsBEE0FFNZW72kmEtUyhVscb
BEAceCW5F6hdKWY+KWC/NMW+tNpfQbN+z+nmEjuUJnK5gAqeaS9TfsXpNT54gmlPA7XoA2LrQjtA
skKW96A94l4bV7t34QroGsGaCvnitmJxWEzT5KmSRi7mij45PFzfXv1cEZXzv7vjfP5kuR/sTETL
mkRSGIDY/Gxx5LGF0ryV6YqOTz0wbAIzbMLIxydYKTlvMrlYZ+PDm7/ueTsutMhdNrDkbScbaXr4
oDNkjYlktOvfD7QRYc9DB9sa4nBtl+xPJbZyawsb0do2vdSgZqM7B0BzP4mYY9K8acyuwdmTmw/9
rqj0R80b2krbGM43Fpsb2gMFbYC3JWduvXp1F7ceqW+eKSptu2Aop3QkIElnfm7ROL2bUBT401eL
x1tbbU/lWT0UG+cHaSqVsEwBgUuZRtSvd5eT70JfVgfWMXO5uoQ1WC60ZolbjA/S2AibfsIo1+sm
RUzdkfi/JAVEQRKUnkD50DIy5woPtNCSQPiRXVdJmXFI39A5qTqaD/9CCyHWcfwk7ZYUTnX5NGKN
UDirx+6TAXuu1QcfwxaWlvfobLuAttnX4COEv0OCJDzRltoKJVDqOe2RJ8TvcjAYEPmKZ2m+834i
wrKXI9IXbom9Qe88NPsTkDzA5enjrNyRIlngNtf3iAdFnzvCAG+qR18p64y7uIp1OGLjuFBKQBLP
vs9TWGPaaQBhgk9bOEjwdJMw7D1dXXkyysxMvm5RWfdvyYRGTJg2BKBndaTFmM44p3uob+ItHoBC
ghK4idjsHuvcRrBBhTuhJDTDCkpFd4n2QzPe2xxMNIFoEwXFm77R9QydaJIgMheg6v84GVM1i59Y
0SzgBR+IJ2GEHgmwalSBh8VHYhUZIMtF8oGN5cxjhxIZrBhlMXyuh7bQkyDJjNhC/wrZqchVGx1C
TBA37hHXwQCOlkzUxHV5m/fluJ0Posk5VXOrFFqeKSUX9Ynx43Mbgu0sD20hDuv2ilgpqWQbJB06
RmOJtsFhlPKXIwKNtDFjz+1bTtcSRRNLNb9/FOQbbBRDeoZphkdhMv6RTtNuQf5mwujeCiimVi55
jCc3Cz2j4sXCP4wfGJVKuYa7ex7Nt2nphyP6yNq6ym9T0Y7fEJIEIE5YY5LDYsZjXf8SI20hsHNH
vmY2DmYAD4pV/e2vBcV0zLHvpt0dhNxTuOs2AZ6Oh8/scGrTzL+QzY5FEQJ0PJzlpCASn5LSu8IS
vxJQEfwsVip1wCI/p9V3bH30v0jFzH5FGtwGEs5tzSBhymB0IS0IWMDJYWaWKLy6oCfWIGuqdoJJ
zfY+R+f5m3sGRVOMOQf48jSaEUePARPlEOldrI1U6KDa0OMu1SqYNY3/tYgw89FesUTj8N5vuqn9
PwxUX4VEoLiQm68EBrgloR68XQGPQ44FBmHK26xpY99uWMYPt4boFxJWpREjPTviV1NpQCZQ6XK0
Rp2VVrX2HOBDjHtWNQkGsmHtxCc1MmJ27BluJ+P3kmXSLjHtd/KQ7L+ythQyyOWTSezLagD00fUE
gD+ezOuf4lKPstJYBsxu7EXl7vOcnU7n5lnkxrdI/Dn1JUQoLyuxbFCRNbJ3NhZQsD5uovS7Zuma
X7McKuMHP0ZJoTX6FckJr9zrFB5TROX5xkWnypqzy9+U6rTeaqbwf1KODv8feuBCZ5MIBVXK3hq0
0oQ9eNF7I5MAtaAzpdkC4E/Y1521+lgyWN1Uasc2OW/XeQptmM1nGwW6TNuEzE3VmWNTy9nNBl97
8G1ABdfqnqtqfLu9cD/dfwN78TJDQesXiQDl6BoWFEGJ6DWBYwBQ8CjcPw+YPYQg7/gOfwuUpdEq
AtvIhdhClKBELbLVVuTi30PpiucGEYJErXij+bgJtyxbKqJL1L2KGdhBvl27lEMgPOL9riyuZBKj
ilJtBN8If/MBATE7gVtXB4iQOezOeuoBrQys/uLXI3GMj0guP5CTk1tdqyrZu8UpAUQQ35rjsM+d
bNv4D1u9V53YWxsS06mAQouPjafM32bvcLCWlXTs3fPMgFL28vpox8rlojwtYwE4plHrck2xhJ8G
SuLXi+JY7Ljeo+87M+OPctJa4CECHfB15RFMaA2V4uTUgRARBrYPs5b89pDH2Fna9T58d1pkaRdJ
d2jwvdVZKBvPA3zjqEtQk8+vogPOk1eSJtHvDhbbaNHqK39DmDBvIjydMNxDm6ULSJ+0AnI0fNRp
QHDlR4xtLekg+gHU4o5VHfrtrkjtxBVcH3pXndUuehiNADtZm5RLSEPPnLLSlTVnT1qWNO6gj7rp
omKstYkMSpSr3PdC/k4GmvN18oSoHDRRubWuGCHgFShhx65xf42Yhk0Pv7R8jKOrhUCGOfnMvP29
4DnAmdAMsU/kYc8acsU1aHAq89XX2Pw/I05a0HybNEIaKKgC/WIOBh6tFMrgj31d+L0rAqShvAYn
DCQPZcrluzW76pYSmlTNx/2PZI065lyoXlFsTNfhUUlIz+NA8xeqKyOe4Q/AIV1vzRZg6VE6b0rj
RQ22jPH2gOGg1jgO+t52MmrX6phSUNX0tgAYdOfSFIvFKhf2BpiUfuzFu5ciac2PE18gBZ5eDE/7
mcAExufKbUtRFewjEndFQTsIFswNTzss7IDFr++DJhEhC+gtbFq9KMCXRx7G/VOC0KOQxvsVrkFH
vRx1C+B7p61v2mo98snbALz1QBKqiOayiSRhViUV9jCeTpob3XeE2pv9BYSAWiiHSZKChNrr4mRZ
MG+wT+L9FChJayM/fjvNw6Pa/Ey0VaAti0kmN1EBQkvK/4TaVYnxlSEHb438nZmNB61fWx3SyyvL
SIygfne0aYaT79C9tdw4b5NSxE+s2Y645TgZch35GAGFfd6xQ8I8vkZW3y3QRR8oM+2t8w9rnBmD
8EtwilKiIosOi1GbVgFA+ak1OEfC+h2pmKY8PG1dehsd+pwIvLx0XNYUodlbn43XWjHKYI25xKxB
VUsfmowWE/zp4vqFJHeVZ1LA5r/W5TSAo2ahpJUT4L0W12oZlj4GBDSVovQohK0v0Ibli531gitl
yGpmQ0V6y0AjfUqq62EL9wmpmNP/1cw7ExCZNRLi2ncvySmHgEbi5zbWNbSvRsq7QU6w4gRGjsS2
DTiZOdm23ruHz0RYWBRpwTiuvvsVbCyXyCU8DcPkviZQHgT/ydIln/zCcWa9zNMbHAPn3nhwyz/f
bhVqNpaS/XdhQl+wNDDD8llKImhIYHOgbVaYxw1IXEr1sfGUVvc7u7OgudIZKGwbfCdvf20OG8Wj
xVjr8p3uBgT53PF0/hEWB9xbr+gMhd38WGieJC1BO/JXnfbMj7PgxbYJhVqyHnHoXKRz8h3cg+aF
u88g1vjIchkEv8YF6ZrTFNrnlgy5YbuO/ONwNuyX8d3/GPqWdf1b9v3mkuyOhysDuwgea/z54Zgv
1zbBeff+jPZWs3aweT0DsGU/rVsO5fr1UJcWM1ZrLkHVtganXVBBwD/Lh85g8XPBcsCxSals2WnU
M8TnnxanHcgRmWJXTWk1mVf9aSydpJEES24L9JrVFaGVCb5wsIUub6ZvRb6hc86Ba08KjvwxqnAQ
YhiSYylg9ZHva5RzTi/fMk5homP1FujnWhU4gKxMqRUZGttGnFd811VfkjzlY5r+XXhwRIYf1nuz
eJ976iTtk5mRTEVqpYtZCI9N75aGSjY+hPhVsc9/4silW2QjNbRwkncgv77yxCYs/EpQb8mGcw30
ODlupumeZa/SJufcEwDiIAfDRmixVxJbzIyMB7cVMI1u+MSuNW3UordeYwZ9cIWeC0gsstGY6SdJ
KtAZsKrxiddoQNIIqtOO3JuPbd+/IbXO0Fq6iJPozWHb8KqVJDf+Ft5wRWeB3KO27B5SrzU5Qkmi
Wc6VtsM6Cxxnr0nPMKHJ1BjiSLi0c8JDz0PUDlxpxAsvKwb3DoGeFaRj5XEIldsNUcEDZ2Q5LW7p
71w04h1cQIOTgdy4OP77qe02jwR3W8iLe8Jztb5awR7aNbrvSXFFqmc5K0LHlJwcaoWMwTCMxrlq
pgOylr90CuJ2RkVZJEyr/BlIj2AdZ0LxnCHIwS3rX2lve+Rtas3cydCVxV33EVZpZPJHJSORT6I9
R0ApOnYKSzEJzKvpWbC54j+HGEfe6/SrV00mH0zYZ+6UyZNOPUxIoHMPX6iMG5+g/nzGi4dL8Dmg
jaMs8XW7HyivXGPJNsXyzYjoJAtrxjdpeK5q56X9l2vU/Xew1ZmTEdVtsQo2PX8jdBHTi2tFEUnM
/7od9lLCnU39bXh37vRfLTzpOmB7gbQJN1E20QT76tst0ErvweqBLpN5ItUSqFvjO6NFvNWm+vun
zPzJgg2HfqGzgN49Ubm6x7ZoC7EbxupcDP6oia9LmY1ne1fBhN/wWpTqp6t64uT0LJqu78MKWcqF
kGMOfKRbV8wy4l6NlDVU7nWdKH0EP9n8NZEXNxh5kELgnblUXhsJXb9jb1Zifhm8Mq2LsOpeqlYL
x8NriTyuBlwYmN8TXSVXAsmor5eSeA7BW984gs6GoBsO5EiXkXKtjuVFxz7x/MAL2wNbxAgtu092
V3P98DNkQUIH6PLOEmwxi1+clADSYG1sN9+Wf6bHvWjTbjgdq5Wvnh4W4kfaOl99lzyh12piPFLz
V0AerF2NBJAxgTGA91R82jr8VmSGvi7eStyXbiNMVtBpWFgxeLKCvk+W46cLY8+VBW2Ks9RFnc4m
6xqqC1EwGaLurUNBLmUYt1rgI60Jvgq6q4t6J0BvrSxYpWeufeNYM94+A5fOPbHr6fSWn9jy6mLE
IFCjQn3B9WBLmKPi+ByMbt6P0Fc3DAF98tljEsDFmAqzcRPVdSd3RcRM5VBocWZkIXor1thuRE68
XL0COJ9ScziVawZLkfHJR3tpoFOj4POE6F545rz/SavSV9SQtIZUgjgeJEbdKbz71Hu4ju7Ua+Ja
bL1OCtCiOtlNvTRt+fhxSGVLDE1QfCD3AeYkc7ffiRmJEQNfani+OP7ckBhoK4JNXFTF9IAQVWqT
RbnYBMGQwNPMmY1X8u+3+7hVzoR0URH1JYpyf+rcg/K98sbZBA9hpLIFHQ9S6v1fI9UT0J7ZO0PI
/Fnv/PoCjG5NtSPy7zoZuDSW4TlOjSge/ouo5zGuU+gbV3ylfUzNlXM/Gxqap4cgqqq3n1hn8INr
TDtETJElMnybenBEJybpsuY/uDmG1xc+7HynXh9ycXsZgLL6vke7cJfXPsgCnPFK9mgnJs0bjK5m
WSHkC6WoxI1I1eaibAU/aX7MkqpveR7ge/MATuCXjE8fL/F/YgXx7ZcglBeLX/wAEmRo9YWWzdoX
x/SG4IAwr1I/ep0AseCPTeLyycww46qn8CQ/FHD7ESwgOegCTGoQMFryIKQdONo9pfqvNkq5WfVg
IbjaEK7aG5DT46LeV4pBiruG8d+c5nIvyMdrwEf0yJxr+s4sRb/W+wBHs9ekMKcDXL+Qo9sMc9Wg
REqIUrKCKPyaiuFGtw++VAyJhnm0DDL0xNBDMbQ+81BI/UEodLH2QG+Nc9IAWpEeiqrXZYn9YgK4
M+C/NiVc/WiJ9PnucqYzCV0ndct9/glm08cnpduxFDGwE9Y/sIAQh0LayuG1h5DWXMJp7iKyYoyW
TM8x8osVrI9Zv9676Q/WxyLhAM9hh8G4x6Xth5In+1rGZlDGJ9j81OfMSxuSEKkaxN/GE4gmZcez
qF3OusjdhLZ+tzepIWSD7BSlE4VUpM2Tt/UZs3mdzFzWOKW+Q+Aa4ox/3cMCaZQnZyZ/WRZqPqzC
a1G2hmlLPMnulcQG0yCbSAXxUtxzOjY3w9XDwy/p+Y8+OtCV8DYKqW9dySc8IQEOD5OQ0dqJFSsl
mzZEkDGxkWsj9I/tIqUZBQhKIQbkBHHuAVzcZr0VswanLFWQ/zGppdMrjIDcXBoMsRk3C6vb0LKD
6T92BchBZ7xmsidbxb7peLpBydCGnL/YtNr+gy+fXR1T3A+4VshzChUY28vDr/1j3yQAoFnbT/QY
N9ltrKopcgbkBIyXTZrhYxooedVoH2FGdCJJTyUWS0sHWrxA0NmLVI7J4uNagRqhqXNS7MtZqAIF
DwC35RMQvohnRcE4Ojd1gZyVj6F3Wuhsov66Plkp4KeMhxziq3HdZS/NE1Q7u9wtFu8+i76DxSGh
r41tNhtErxWFBK7sSUPGr3i8qLWukUYdXo5pIanSpMAB1tlYwMx1RmLLOT2FMzqydWSrwy8FpJlq
zqDWLpHHfIqNHMZVenQJb2Ei0seLuKiYFjwoZf+qzbqzUfDVhtueJx4ulZDmnWudEqw2ztPlHwWA
SYbyJdbU3Lft1KXNJT/wGbCXT0Q/x4ESuyTylW2XKvkcta/RxpoI1riyEXivx5Bl5oFJG6edT3xh
TaBH4PMsZZcht843jFc/TqNEVDlbiN8IXSWWm2s9weKDxU16T5uZIZczUCJLes2TdtozNU/F6MO8
qF+YKWvreQ1S/ZTBL5CxGRLxIskM8yTKEqd0kSpN0x0he0QudAE88DdfqdSvYcTUNR28ZTC3yKY5
ykbOHR+P1Dc/Uzik+49WSgFP3uN9h5n8faRT/5wVWZdF/RCzb40tQKbc0m8ELxBmbrIw/PHqgIfk
jYMAgc66Ns0a566Dr7w/oJbo0b+ePuAY6JA7DAppJmAdM0qHkAFyY9aAvFyDvQ+cf+pV/QtDnlkd
NeN1OOKR/eaonhZrribHFZbCW618qnwkwJQ3B3zGcxvQqLqX4XZjS0k5u7t7iPQhdx1B/ILVmIlb
D92Px7UWsG1kCfYBze/ETd7j6o70bDo/SoPTwxaigNkaj9b5zXq98emQtjM5wmz93Nb5HQczcoGh
a9SsUi88e9JTmN+E6UhA0I9VpYC34uLc5pUOzqK5fB7CYBXsEf3MJk+2jUw02Kx+MDeggkrWGAB2
RjdasFME3yMeHYZVJC9Gx6Rzo87cY+3e2wAd0SHSsXCqP7AUwBrzFtoCL0Kb71m/2Bu/QhsUcrPm
biAlF2Rq5TgZAzhE3+K3H//e9cPBQBC0KUeGyZAimonwPLdx8pUgGmUWQ2X5De4I6kRafmu1lWsH
sIjHy/ugbllmiXfFazvQ/Lx2Ngx4VrFVCuwkFKUFjloOZjwZV2mYFm7p5y3+A5K0L2JT9C1DVwD+
tOAbb6CazX7dPE+3wfPrkEPQ1QD6bAypxXAmjrUPCvwWVb38Dkv8n00dZbyxTEvELatgu1F6OV50
Cy16ltyBP1x/BrxVHkHQ/ogTpz1inIvN1OLIfz+xJoMOD1lTA/zUhB4zBSOZDcm/qm/cQMwJC9hn
Iu6Nd0k7Q3Jpmb1g8uGiMHD68zPDejNRMj4/lYBK7/I/+DsuhQ1XJ+JB7J9kt7/UiRpkHhsQQKGi
9qvVzuUs42LIjolHIqkaY+96IQBnVuxMvDOjoyhGdP/FHG0aSVQjpMxT8if+kfv2jdzZirDFny/N
rm+Yf4h+XELsG56NGIcgs5MZblfq4ENdKUw0rEK5tQpl61tTi1godz+6fNeU2/7GmqlBT+uC+vxm
ZvIM/6HGoy7PqvoG64Ovc3HoywOlHr7P4Tbx+c/cMVt0bpbefB/oI7dinLn7rGRFwo9Nuzph9NZX
YPZ3rKoJ63zThhniWoGJinQ91pUjZxwnl1WVvgrvscju1EwaNGald6eyS3jKb1hSx3hq8JEPom3L
3SBHKYdGNDeTj7Xuc2YbasOhLtkGtQZ0Nl6cHj5lAT1GuEPYKsbOhqW+Bvx3L0PZSt4EliwvSlCU
zrcdWErVoDETuJ9I7n+3e/ke5PRD02jTMkDLxoF8yJaj4O2myl2ZkGzFYQp732cIZtJ17NEEYcNV
3G3k2+mzX/mFXU+nQmG1GUwBrGiU6LXuEWfFgIY9k47LKzriOKGgCUSPcfwPi6mM0gegrLVk23oR
C86yl6d2ivDB/cPBAJU440CQcLX6BK6DpcWdRNbcoK1NZGRejG8iv0L2dbmOYtFM+igD6IbIsTg3
1SYwsLSvzoHqX78Z3Sq+NNoHJqdAhlXOg55qI9fH5RUJqfdd8C8Vb5d8OlFo0utey5G54kinkuvZ
jmfAC918hzdthbHSov4tvipTAGyqFru0YXlrk+fMVZZh/8dbiC5LzgP7DMlBovq9ttslKkMiu0hB
3Wtzhujb/Wlc5rpMSrrro+Sttu+S/6j5FWe3MiCcRYu4bJ3+cneEu33YBGdYAOopkonZORR+l+d4
iGeK9bUdK4wHXHRqe4TmJOOw8Mpc4a6BX3a5OpIT9PD7YEpk+sFR2kn8nz+Bwh8XpgTZ297IIXW6
xMGX20KNtQOzogy/JZfAuRV4Ka/w6htIZsF4VQ5dv0bz4SidgUaSYChg7cFf+Y+muBZBxlZRyP2s
me70qiZZs4LR/FxKHh3VRZoiIYGyJdXLWI0wenZbE+osJttheOk75y6j+YAqS+/4+ApIK3gpXPl9
PuZIQQDGBNV9kxZpjlu2JKzzVfMbt/8TaaGHxwxRBkoecJp0GI+Qb6h4WxSH4dd2UlS7jj9dyk8S
/9un2YGEVuP3fkJehh9xb7n8EV2mK0iUj+pBWMsfDdKE2Q8KNkxStRhTfQBoY2wOGHeM+LWqaoHL
yR8tOipAJ/MCFYFDxGMJCk1Jy0Zhx4iDVjeIL1xAAKVghXxcJALaOlxTGWxWTDWajyftEOmhL0vM
zrZMWv99jfyKF/8k9VcpTsAaDnNlyFkFYalXmIlBySkIMVZ5+7dkLX5L5jUAVZPaSJDlk5bXdGHW
LJu281ScP3FO5esVFO2UHs9WX7VyoC6SirMxsikPeBEudYsptXsWivJcTEPvDEwH0HhW/221H75E
gqY1NZMnca6OiIF17BuMUf0f8LR+hAsRNNbQT/zwcD3hbUHNSbxjtaaQR1rhWCvzAiwsgGM/PPTM
RvZpx2OSjPx9Fttd1Gbz0Dd57EyCQV+ToHBfRKJIc3zvmxscb8jFQWlrlGG67rRG4B2kdZimSCxI
x/C/Lh6SDt7pnkQtdHaKNnLF1f2Ew8EKeHJqTLj7QOgLCuEQ3lt4gUdJB67xxQmICdkBgLzish/Q
X3Jee+09niTjDXCmBBBRX0mG0Qm7EkYQ9PgblKuHTj97ahGGZtq65bvSgrnDMNfhOBFq0KkkrWbv
tZ2+v2zYJ6nFDNC4A0BCzej9uEcYaxXk8aUdF1jAVLjSeC0rTLfamk0TOUpXl62R6WazqKGeXx5f
GfmDg4m/2OGdpGF560/Zl+M2b9xczod5dev4awN1Sst8OKucgmHgvS2xys1ucDiMLE2pb89LyoVY
QlG2lo4sb2w23UIFKAUncJmvng3pQznA/ANKZtX98eFOxqIZ2Hw0xiQTW6kmaRyCP2um1qGjpwxj
QC8iPx9GQdije1i516DjPKkQD1A1GyahdmJzdUxUZfx0F+PLakIc3gF1uvkeW9kiuFRW4OeaD87V
rCLwIn05AtOFoirnkUEdoH+vrHnE2TT9zwirFC9e1phmpZtBiOqZrgXb/yRnDJA3d1B/s9YGymUq
XdaZOr1rHYPcNQ3TU7EHKKh3cgy5dEZWN0517eG+GGk8VrU9wKpOGHVouIr8sk4/A/RUo56Vk8Ui
3nSkaJVyKFBX9CrgM0DrS31PDFrwVVMN4IZbhXBO7LUhYqqSBG04pIn/FnS2diPM81n4zFSorZLg
jXI58W6d0ztHnVrQj75m8AQjUkxbY1SN/nGe5KfTY1uItFbTHBLisoI0c/9m4lhUiDEN+0aPzRod
V2JfDQKEtT8wuKHQ1zuZVFYjrEjuQX11nLM5WfIw6r/zIFC4XP44KlrZpMFhpJbKIhCQoD8wluYI
/8/kmu7me1IGRYzFXJEh7O+nSEKFhk82DiAqewHpCdI/Ln0XrNTuRHww00E7p4DH+1BqJDPhncjz
DArUc4kIHdCYWArko39L3YRQSiJ/3L6j/cC8u+rGFwte2RwhPZp9Q2XNrg83gzs8VBC++Fj6L/oY
OLyQ4EUujymkC0Hg08KlvIA9WlkfnyY6HZWo8aMu5pwfQsoVDJo3w6oZeGV2J8+Gvi9Xl4h1bPkE
JEwg2M5KYQ639gLvIw30Jw0P1AdowtSXPMFiVI4JLLzWO5Soaza6bqqkM/xlXRokn7XDqrRI6JTH
JI2SrIKIKfzCqT75ca8kuVtYClL4fdGmxMYc3qlnh1/Mj2AhcwUfoKNSjS18wcPSpLkwd919mvA4
xfbpRqmKtQ033C4Yc8mTfHPjMzJ0dR71nMDpLLo235Kd6zPcy8qczfH7jJiQbYIuQClo3Mgq8HK2
WFLzSlD144mKInLpMA4BBVpn6LDEKaFuFo4PpeRVHxTu1OMn/2JtD4jsNKV1zFO9ge5n1VqMyFF+
e1sl9leuGrVI2MMhEVisaGbWQ0NrilpPiGi07tiutdzucp7jjDfKIdN2n/QYW8zY6rhipjB7GdwN
5Y8hXc5rgEAvrmgpQGZsqFAoX47e6JCbm9a1AQ54BA/R3Zwv13vZ/LI60cKzKsBpeG1Fvz7VRQns
xPWTw0s4npgHxhSE4QJ1Esd1h2jnNHZcQrVcXFuMtLbLo+rxZInLVayXgj/tWRm65NSx9kSHVVcq
ZTYJfl2vproXM6f0mmrL4eNCVjClw74vRYXfwytDR36mKNmYCNxOkjv2/ExkTjM8wv1oRNAVHYbN
OWI5UyFazWHC9noHJN4Lu8Mv8vm7ih+NtIWW8e/0VJgA1ACShmZj9ZwtRLm2hTQ8AZDrG4MSXusy
kH8hQcOl5XDNAlCuC1wbjk9b8fAUqoykgCmxc8mGQHq1YN60HC7ORVa8E3FGTVnrFBaIylpFbfF6
MvsAge8EVvcVkzwQ+bhjKqJKlSSwhT0uC8fI4EwMxbFwAnDYpYFSNdBDKPNsfQTqnjW7dbK64+r3
I0Ozdtespe3jvKbfUtR1qp5gU7iA33CPKiXr39Cm3YIV2g7+RL5eSTSYt6nNt5PT1y9KMMOGamte
6JpNJyuRXklpZpTeVr4xjsut90W6m4WfxE5NruRcAR4zOlch7ZP7CWcZ6NGh1TtKtF34fJ2Z1ml7
U3oC03SBid6dG4XTLHSSIvAWD2UJBXsyEDKkDsCe+OKORCp25lvHBl3OH+jsN5Blbu5XLKJ4P/nP
yRAl66Wd4w+KqVVN6BeRVQl3lNZHeNNAIcuhsEfQJ8M3/aPVtwphf7TCiiWvbSqWRbYtCJxnPwk5
dsaW/de/gQjn6y7Mm0sPn3ouJ4be+ZtDX1dk+QfjnGwtVkcv48FHGBjX6pbvpFE/6ZcDXn7mhkhF
N68RO1MXcaD44AbrYbstQcogumBHCYliY9LHaR3Q62kmsU7drB516VuU+ofmgN4INfcETDSR8Wl4
Hj2EEbvhuV78JZ2tq5ulpUEhHHljqdHByKpwSOES+5YEriBz5qCKQJfO9okh4dSYIjwwje5aaKF2
UySi0e3FAwBTEuEHfu4ImNoEhNXCIwF2q+TO+doGGUSEkYRzIkOuKN2Wv3XzWtiXGwnc/vNiKxWp
XJKCa1nuRkLPEqIz/2JnyVYsEm7BpL2CJnWEsb4g6WZfxrDzxLlNUt5cbGzNzkf6He9pVZkot2EI
WuHMq5ZOg+h1Fw2gVZi+3HWP0X/aFcv3P6zqaLwV20ksbpVRfWVkMeJFPS8TTTja+OP4zwEpo8Ok
O+m7/gZ38iOabAhcqNGGBFl9kwb40G21DF2E5PtySzUGF8sZ7ThGPoPWFp3IxZRBBt5oAbVo1aN9
exZZMMIg0WBO1HIUtZ3xUChtmD9XgV8Dcy9sjUcJhlJqxbAfPDZ06IoEWfKloeOqDIuuVWt8lVbw
DxbD8HBOH6Y2UByKJT0924uXsMXvxRqfcJvmbD1BIrH3KJ/vBYyNZUdRiiYSQRGoFGTj0XhbJH4p
B6SlZRMqto0H+8JmvnyhQvH1Y3jOkM9ApwOc7rFLR062JT9PhditjadEDzyx0P+91Bigyu1Nua/+
4FMofPT+KueuXrALlH2xgDZCA+G9DxaopTOwZNg2GKTcOTtHxGwVGei0/PLYuvQvu7T0Cdri1Hsz
8hA7f+B7j/vK6/yXCOleUNhGOWQZpBZxoCdiQ16ipDkdARnLNHrkjz9xvHjtJIqoWgqEQyGN6nhv
G/FYpDLNBHeBnQ/Ffx+7HlO3r4AvIzztY/2UafKevRBt4e5uJxoYjlwGUfhpyP3pVCmbL/E0g9IA
jIFlLfJBrFXiF/p5NGOY9KtZVbykfwCJG6lUtgNXMWQS1iB6lBLR86STJ7P6ZdscxEj4+HKQEVwn
5O6sg7T+05Nva9O6otJN15v0mT2HBfGzC31CxIo4VtTNOiduKR6e9iY93J/f+V4uvsQUeLU9N8zh
BfqJZeOnaywq2StJIqVM5A9xHT1BSAdGhm6cHKoGuNHCw0iIW/7DyD51Rd4fD1wjGSIGLyD1lGAa
5KslD20sHWNhBV3TWhlp4oWeGi5ht7PJt6L8Q2EUIcBucqZxmrSIa6rWnl8lgaox6Iqcx9Y2O7c2
LFRkJFW2ZvPfioDu3wDvCR0DFgnoQXmMYTDElpbL5hekLX0QhjDEwfaHE/HPd6T5Z/Xtv7dNKMda
o4jzy2/uy724ifp2Yxjyj0VaBXFBiE14BDG+caasVKVGLs3730xhJrwYF5I5SIMfkYh/2iEvujXD
y/VYZPYBsHW3K7wS/I+o1pV7lAvRkrrqu8/18HjhmrvI5E+aGHOftCJALgcOY1FoBdx87oOq8vMc
wz+n6grBsqnKIPlPQDWZY5Ju7a9qICSwCyMw5COHn5sHqtc1VWJBv9oiXlevlXc6ZFkNf55AwKTl
DpguG3CLbLbPKKFNpFbPk6S6TQ+xsZwGaLQkxdyghBa7iEMxtm7UXZU2TXT5NvA8f459Odm0la9w
AhvdCK82qyZ2PTJ71r+4YVyBrWgyHDyWHE9rcNKzZmDoaIcdB/oKnsnIXEuGMcKMVBZxNeansCwu
kImTboE7KHkn0ppaw1FCOY0bUPD42jervUiHzYYsrcxZJ9WMFu0bWvx/0QNxljhF9vfG+VOe4f0+
78xPjcz0GVWrduKFLcYh5s2Z8DYXOvw+h01/HEy72AH59jjnHamb6PVlWTa2yzbUmQ7RipyQNg8C
k3NtToE7zUu4dyQqIAX2ECVBOKeUWDylklghZcKSJpuo3HJUJQgg4dCuYWiA1XhRlw57sZjO31T1
l/PYTYKVFCsKvvQLQ0mCOr82FrEip89+NNVIkw70tSJmhk7mV7n0tRtzilOktJRAVySUMX+jctK0
FS+F1YXk2udelbxK1BOjUOT9loJ0kkSmx1vauar1F6tEJErVWxzQmJMeI27SIhOI83PXbNR9qi9x
n13dzyZEYCwXRQrT9DeTdk3ofgUWdfz+VkMmM7qpHaGqw7bHtSj4CmZHpb2o1QH7+JM2sxKkBn1O
v4piWN6qEhpoNEdqy0yKUb9PKjXd8JOv6H0YZUZWh9SV3k59OozCu3wzemN/6GIs/5IpvOtcNsMn
igUo4dw2VHKheHGlgODDu6yIoFLgain21WIXrCWznp3Z0XDRlmxS1M96mLVEHnjaKrB5v7OWHmd3
pHjC0ih9XHYLua9UZ9CwoDKBeSady+Kgpz7CVqyr0o8V+dIrFiayiEuSLqovg3GEsOUJr/Uhg/5H
RyyuFzEv5/MfGB+eKAWGJuYUZSXFfWHc7g81xL/HaqVpvbP5yyOjXbzan2CpKb5uwTN0U38jdXz+
sJuAtTZlKu9JaNc/kUWTFhyMwHLzRyOBmfCQJia3drhZaBGeXhZZitJ3QXY13zxN0zhnVS9ITvpe
eydW+CDfTGSLm9y8tUax+FriAEqQUhAUHEtYwA/QI5jdyfVeQnIDyzOYxkYN22PGd82QyenU/LRQ
iTKCj6WSw7DwfXgpteYM0xVSAMd8vSerJK1y1flF8ZKFWPs6Uk9FvruXtV5DrSTClLzGYG5OjIDX
IDJGTIc/XKfXRENdQb6UAG+Kfh5TqMHDRMRwqc+wL72DsSBy+50rvqR3c9I9FYRrB+oqIkBBjMDw
vBqA8DweIKkSzA4eYvBQur+Y23lS2lB6FmyAqGM9d4lnk2GwziCpfvkJb3nhfvS7FZcBbsxYzVSn
yQfNaumNuIAr7IpXzpCtUR7F/yrGqYB48/p9sYsjVtaE4o5IpppQl7zD1AuPGA6/hg0GNpHZ5qyf
MoPI8X5M367zl9NZv3AcibcMTicQ7rJLms8dY2xtzg2aO9Qfc6FAZwq0OAeIWdkHu2RtGXgpDFeQ
To56F9VGc88rrbOUyS0wWxdKxO/fvsrGqPj/eJHAuKLCPSrN5Iic2l3E/YTOKds5xFciH+TkN4Xu
xzN/14yiQGuXhOkWq6e5WM+J7tp/lXgrlkrhcc994/zzlWd83ehYJ3GmjuOYk+XUN5cMKLr0iO3c
MGs8TmrtvBJnVAkEkQgGiRHPsvhg/IJYe0L8hyS6ebisayY2L2rXFzVx6VtpWfvE7vzRLSG8hdNt
Qzf2gFxTyxudGbt9apiDRSadF5z8zUDa8mvtxTqq9Y4EarM8rYpjINOcErAs4M/jBmzPmzpUMNrB
SDH5sjykpH5Y5mN2OTrxXDabm3uGaSX4F5aT5FY4MuEtNuXb0iEuQiWXcXySniejCqRJ/SkTrc/b
cL7ONHaVfH6rQV0YShevu2gFwHYsFoa0uTpgb4vU5TggBmsYWNGGyJbxvh0q4E6R4F0gtzFdxRRV
mS5l39Nbqv0Nm1/hXt2X+z08TBwBCwWc2ju7zELxnZ3OCnY44Mu/MqLCTUlH7NbNyUFniLwztJPl
5kR9CpYq3iFqGzaTPdxe1NV+d2MIUraJ/7gXphCgjwVM5/1B3bBi2aojj4siSEyBdIFw5N3rII9G
SnBGASExCVQiXzFyGv7TDsmovgPb4FdwGI4TugrM/wUcEHAcK4RUiIAsVZtHV1fE9uZl1fiOVX5P
j1IEy+KAkk8D6SSm2No+F9XODaJQGMoxAUwVqWAD1AVsugAouBf2misMLxhyI5v04yhfBHtrlfdX
6p8wZ3IPojbpNrZ+Pgn0+Q75fWHU3zE6M4LFcL7j1qI93YZommeY3bn7VSFKCnACmp1BeGg3VDgW
TFyam4wBrEsccVw3KvRncwC3lRu7NYJl+LmgHp+4lIh6z3Yqzz5R54gXBx5ZE08OghcNmnatBDoP
E2D0CA2wGBVisqFB8dOIFH0W03G5iUnF0qSa2kzqADPi7rf805FqhYdISBEwgsoGUxRqBVwl2l8x
cf7o6NSMYC/uVXpMRYmwMiWED+It97x/M3LPhoLfL1ciOOyL0FQzLXZDQ6TFWM8ao2vZidROrkVY
kfQtiD/0Hqe9eN0KtoTfF1xZZZdd5/C2LB+GCK7HK4v6nL/UXd3+njaRR6Z3DpYKAt6yV5SQbyFx
sP0oVkr3/AFQhsTDpKTbcGVh8oCYTlCydbKa6Ny6/ilKauySvoM2ulbFmZBBZOCrqjm4THKx2sEf
Ubccr2sMV6YkmMkgFuqOx65o8q5SMRC+GfvL5Ly595jrShqkfDbcgiI/c1Moj8DURKeGh+v8hmyF
TsMv5Om7M6T9gXnfWgfrX4c9nzBUk+UjNJI8wSOeMlZFqWqEHMKHM0llajnjGOjxUcFaoplhfuCE
b9PREFh77n4fDMhuAbO4UkZEO2pgfjUQkjD1LGyjfy14xjw+ziDds8RmFyaDFB1itj9Ne/lBR/t2
s2hGdvKNBnR93Yp1USrwoi//bDQTlTy8RmnDxZt8km0M0aCA2EwV7Dfvq6+Ild6fdnTHVQw1eUCw
H6zUa3dQlV/pKc4Pb8gnTURWnV9i2lBL8df5s1UWBEyS4kxNHZv/aHdvvbiY0/aRC+ZvV/xy1acH
jQNelCUqHdhnT0okp5wbMpiUB5PqTfHSUTh6NOcZ+TZc767GJa3wVn+e9UjGtJCCbiMBY5HGjksx
HU3/fgbpei25Sm97cTFk+Ccx8HLZryGGhW6QYXD/SpC8Kza+N+LapO01X7PrOI8qgLdv86TEiEw/
1QaJcnTbhjiqI9yqz43Yo11p2DNQHD40CYVIdJoLwhJnVhwQ0nVx+saSbxYWOyZTD2bjiATBJClk
TsSro297oaeoJSW2kF3E35RadV84NG9z7By420f9TmoVQsVi70sStuF3R1UdQ1VnPguSxYDGxTi+
3HaGbaacden1Spbf4Zvfrxbj3nWSZjakPbAfXw0cNUVVBL4AdchtGkpDAU6rCE1cH1nEM84BdDyD
kEWehTTCUGG8yW930rDmlYvJRSm+orUTuIZ0dqCuG9jstXZldJTSQkpSlrI/FeP1CAvegn6M0UMA
iSYoN0aq8kAasjZKjy7vUYAmQkAJcX4CvRQWc5kwN7PHF7UIpAMdKH3MjwFQIxFEsvblJlGupQPW
ZLDzgqVNysIJnBvFDbwfjLZGcLiAfcFGy2wuKHnDfmIZOJAUArGJw/iDhr6RxdLZXQzz3IS5ogzJ
LyK73r4GgJDtwu70jqEgU8HTsmZI3TxrjI5s1xeiTTmSZsVGHMAx4lf7fRS5T7sRsdBOh/2U4HgV
v4W3B+VybXsH8qqYc1Hcw2QDfUPkCK37si0ai0S85fUafFJX0UQmfx3YzYNAWCBGlYzftUvNNJ/0
CD1h0r2lIfriMaCcXLeLyGA1ZSE15HUmHkcOIc7qEhR7iN+NZZb9ddaPgSZK3TW3RScMHjabHd1W
ag7ssK9XSWVcXojPbz9EZ3Qp6b8Ccb8cpMstNxJiM5BWefZuYlvuHGDC4kA6RPcFA5pte4WiTUD2
UuIfGhveXgFfCU9Z0mHt+t4a6NERnkl5nZ0w/ek/qz6kGPWXxgXTkifI1Qoc6tuV0+bYk58rQDMG
ttZEITuYRJFVbKRplb+48lQnLgCf4WhB7T45TmmlZLhFdIuuutu8rpCNjduSpos4bPgElYL7fiza
Fd/eT0DLD/swDRmIDM9HnTQ2Rg+Yrk8YMAQBs0EajYSMrtzQmsb8qqnDMxlKSrNVOB18h/Od4DbT
hDEaipR1IUf23VAGIRZ+s+Wh1dv7R1YwL6sguFe6TJONfvRWzgynGng5CHn56K5f09NvsXXylRrh
fQH0q0BdoJobbUW2k9p9WVEbtVSwZMwmfcQs+hULpoum2/45yIX/w1F+JztLkhXWrngOjcxRe9FX
foCJSY//jB5sREXqPftTw6gn+E9mMMiuYFNkv/1m4tr39Y+lBa6Y7kfPyTb1GJiSCcgnnuVYkviq
eKA/srUmRNcA2oQSGb3Hk8ZfeIUKMjPZlzLyfWjk05NjcoE5NU8zwKDPjfMkz2e3C1XGGLsMlK9g
4Q5sdadMoqgTA37nWzSlEiTJdBiGR0N+EJKvfvwJ3b+e1jQntgGY9wOGrORPNLVXBPopqwW4Wkz4
L7vtTgwsz7XNhC00ZdYjGEUMbilFMjt+6eFSvHCF3ksfm1IR+Kp49quruusfyt3u+ruDcdUgsC+v
wugAdEcIe9DwEy0EtKncyHlgWk091WumlEQJmyYrz0FezjVNxBK4nvxUgLOfpmxMYC9z1Qn2OCSP
GTadx7XmxhQqdU1N+l3Ozza1rJi8CHzLuSaCFCoGqflPiNllRkvmSqw04c0+g6lkxVp1c6MrJ/Fr
7O03P+sQGR/dCoWcgyEMYaCjHca3RWPvz/LWTNrn6F5+5BlY3Iq/EkWNrDVtx+uBSdEFkZHntT6a
mCLDIdNNFkVvmA+0j48KsvoVukn15d/PXBtBuftUm/6vAJi+Bzn5qSYWQexgWtMKZtS1Oe3O9fUJ
4tvOmTLv+VQT6pGpo3Hd58jru+d4RyONODUQwfmWxtBtI78Z7I14r+693MHnHGBSlQtv6F3EljFh
07EAgU0qmIGDSPMczoy+ZSfY+n2hLZ5M0v5kqWtUDMq8jQ/apdpuUzJSGLgorful354rvykINkUe
dX2oB+fl0FrJiy+ivT7LpH3hqkDstiYfSdkUYq2nsOllzjCJw1JbfXT8vTPLsswy4sj3PsiOnMff
whwneNdRSgmEQToA/uOvwFICUATf2P+y90NgfQfPsSfiLxcExlVItzEce5WC3tsnmYpfwOcnrr5s
PMsTOFViWUFhu9a4pzicGQieRMXNbXxqtRsq85iRXiv8HjnKwAfgnbljGKI19iFkvr4IPcrB6XR5
rovDxwkmCHZuBcdA0dsS6eSDKhzO4f/dQhvQeGpsKC7Wp3J5W8Enaqald1lNJj+apbnx7ZuGGpWY
W+rV1gOsPLxyCFfNUmYClOM/TPlNZI40jDOwzf/yIGB4JC28ydownOi2F5v57AGxp53rylaVd38K
g5I19eOI7y3GmaVNyllfs5domRX/sJDOVtE4nJekUKV5+2LU6ykH8tqP2611/vqvogL2bypkGZmc
pMLmmqdHg8IKCy8g4PzCvlaXLlJEIiIdg6I8NrfoYoQTgD4V8TcWEmeL0YAj8hs8Ithx70oSv9OU
Vlas+4mhTts+bmq7aOFGN1WETEJfNYFVko/cU/B1SjSOC93feKi4WhI3gLXXZB/teYT3sWl+gpqP
7TUAfcjL7WbtAthbg46WB8RGkwiAfdOj95Bfjrf2z1S6rL4SEDdx9gQ0WhBgF+d/c7dek6iL+xVc
Gc4zLMVSqRkM/2xePDG7qDKIAeY2aP1Bmhj6JVHinAdvPjZ9SGUTvYiA4MN2QhFm355gzlP1Jzvm
Zg2cmdqqKWq8EBTTUwzbLovu3YbRzuW8FLUholzIG+i1mI9A/eAqNlAFWgUnGaf027BJf66yCj4V
XgETwbu6zbmi3byjmm5zINOsmbSx9RFQ7TpcZEkwC2fd2XBs2gpaT7CGxTJAoBS74OXS9j2V/kdE
sL4bMEGl5HhlUV8OTnaJWSPL0ByKTve+/6TmJNFAtAPVbcBaCWiEbJBWMtZepOIKKVf87Fi146Cg
X+loXpvqsATzRzzm/Dxl1epmMfyr9RV+as5gpizV6VHIBkaml7Yulal6SfHBeez1Uf9hffywIdya
FeD2qjp3agcVWOkkggbxvb8U22+ytZTXD1EsubdKr9RIowsfHEw9efbxkBRHLud1n+u9wyCoNhhJ
MSPnW21UWQehFnqSKvoNjB8btvyTZNWlYP7Ay87Zx8rX/ACyunfAyrbbpZVTfD8qRf/IeApUCtyR
awJHHGhPoS24hQzxcsSi7Rmz/RKuDifil2vkIzKxiqxIDfpKfzpIh2H60pVyH1hbDcCovzMBYGqv
l0WS+GL/aa42d27YH/e2GL+pXXOY0jhX28L9sSF0a8nvq27ImHTkoY7G7RLTotdBvdJQaapUBmVt
H7awvysKUnc7QS+bPPBGeAVYis7/dteqOz6+0i2xEuXBOXsl1KXYy4EOWhdgWnYRAHzpv3Z0qOzt
omhuYaWkmTX+SJzgGcelYRFBybd06olThA0Q7cJyZ3bl7RIxIrWKSS+JuQFeIUHDj5t8KweVEAtT
Rj8Q57w+kjGVCeqF+FyfyrARLvV6DsCHDTwSNc8OoXLJL4/M0rB5pc/WOv8I6IbcQ7NqPmsIJofB
juVdUOgy9iC/EcsjfqhZKo209CtKyBCbrljfSunzmHinA1a/vtrigMN07eckD/N8weXZ9uCVryPx
RnYcJll0t9/ZLviR3moanixEZg+jwSbGHXF9oZbzoixwZ9+nrAijrYjtad9tmW8GVLfqTEmBeJ03
WS3PnOGQUBstbU8nd0BsZ5FAqKRFT4nF7dllHVIlSfakJMwPYuxiNC9OQp40RwsC0XQz1sAUT5we
0njScBy5Ilshr15u0ITFNCd+tnin0yG2rq9Cd36VDkao1LbzibVHybmc4CLr7Alr+8vuZHn7qk/p
bWOnVDzx9O4SboPJzSqJQ6tpoJJynkC0n8gszQVsHEQR6/xTw7Vacw5q3M4E6PPPgzfMHiAtBmNY
8foQZ/tul1WwW8qE1UtFEIYHKGMlYrJlK6EPl2pYk9BHH22acj243pRlAJs0tHdAc7zlOnrHWFOl
bkAUfhBMCKgi533VmHvb0TE5Y4gaSTUCNJz9IAGkDMRryf99ueSvLfNry15W7yrxPBc8LGDQSCDy
I9XaIZFnpxO44Kko+zsBt8sSlGRPK7kOvZsjlMabkt5yG452JjhRoLHN/AWpe33/VnjwQ+UHiGkr
kiyjItEKMOjU7RMgfeu2yRjbYLrBMMjKzsrG4Ku75yhUfP0lOHO/sq4xwYBv1LAb+12ebxDaQOcv
onGhkAcSYsAxTTakVNG+d6urTpuTzk94Sm4AIDQ4/EaAIHRJfJvkJPEaLSZKvq086LKRbVzs7ady
Ev8En2OhyqbX7rLGJSaxjY/UHHuJJ1SXUrkYhQpodAZyZUfNrAWJvhg8q+PPuKJruBCSfJ81GR/5
t3e+fjSBmiB2UFiBG5DNO9cBmJ8BQEtHLChwnEMajZvpCzqnfMyLzpejb6WTJT97vNw+NKw1TuGW
K8s7KQCrJXcC3ll/XoENpuBeKg8LE+PGsL5/vGjaliiDc8j3+aQs0hiVp5NmnrR86qYfomOErAXB
4lMn7+IG7t+lBh7S0N8ULtsit/epTMX2+4BeFzc0BmW7MrRez3ogjYVWFMUgHCPAsngVYL0VdUq2
a1t9NgBP8UcXjI9e95F+iUtdq2ze4bmXefETwGajqyW7Q+rO6UdIEHsI5HiSgw9SmRAgKrejpFzO
/eaJ+whMTTIsrhfGiFCBOgeSRxAQWRRUmMDAMaMQ5YQPeyBaONZewMZ4Nzuf09mK11gLzSmjfjZA
98RvHKYAPzjmnNammcis5xi7p9b8JutRRuXsorbWPiAXmNNkplYY32KENhbjmHE7XgX7A0sFkaAM
LAfBaiPCvBwVcQYW4JYTU9FWbwAYzbyr+E7NEnSKGqr17WrcKhQi/aZqW/y2OjKzra3fgZSTVVsC
+l77T860XBg2A7QoxMXHaBWd4Fysy7EsqHySl0Yk2G7uyBI6ip/PSnZheLxAntYnnMImgEo/zL5S
OUsbqo68DmjrYBG1py2u4TLo6l9+DrIFRndvs5B7zei918erkWN2l7JIZQeIzQOXly1YcokEwx+B
ED53hqgblxJ3kftuIwfsX8di8uhdj2dtttvJ+OTEDg7zPCPNmD8eiBbgjda9X3qxWERQSGh4O4Hd
H9E9980NWJ7Bbv4T5ZzbcTjLufxEG7oRURBecFZ4+46uFK82XOIP4bsD3kvIMh7BgZiJJQwzQ2/T
eBp1TGmC0W7KxGSKe/WMIvmv/WZoPU4o+A10ia6PNHW+wbiktzaFwPXLpjp14qvuaNL8vJXqlhOY
U+CamsURVWdilc0gxnlkcnKaG2uYWcxag5AwbhDl6y29I1blz2//faoLIugbAIr2rSHt/lqgfJZ+
bX8YoRFTCw/kL2B1C1dP2/meJ3PN2GaTmko4od6MIyqjWDKa/x1FQj/8Fn872+rY3sksvpgbJjdq
yqs1Zp5O6ftv2PXVELGBkl30VB2oxzl8xGteWmaUFiYB/BlVipRoy8Y1NyZ30qdZRCx7PNQP5LfB
7BJF/mfHVt+PStzhWeKMtsRrkOOnEyJJxgpdbKVMx9JgtUOSEYTBxVxoJdAYu6idc5Xn9kWQRFgK
PfraHOh/ee0W6QZODOJKTb05O0RxosJbipv+HykN9dPIxoxgAwm4q9fP0QGLzSpltcZB06jrNfeA
b6GZHtVm26CF9dWajhSNSmkzZ00FwDuENt45ci6g6pRqmKv1zqvKzr/1OFPKjhqql/u0V3grxdV0
z6tDMcQ1I+VLcFSyEl9vzMuXNqdAYY13HweUujV+x8vFEb39yPQMfpqTLsPAFDmAi6YZXVgOSJ3Q
FlpqWVNrH+wqjpaRatW1t8FbQgkMTe3ggQltgb1izKZIldCEVbC0QbkQryF9BAOQwWDgtMWPGLYs
jPdNUMaN5Rh4JPmSwwn4MWifn3kqCz2KAHdsPGcIuz34Rmriuc97VZVIFKnt778JMh2CXMFsm7DT
8JccYKPNIWuT5yFyuhQtjEA1Ueiroj/SPHMMYtVyO/DNlIM76LuqxjOwawImefhMv5h29cx4dwu8
r8p92BR3vhQXTNQFen+Y1mSbDmXtCz2GHTJXxibO5Fc86GvaP3EN71RbF2lSlKrpiwAhvg9PtqiD
mlqjC9v/3acW1oitViU/BTbh6vS3v7WnM+hm2n7URvUr2vMD4oftD/0i0O4jO0QISSu+Wq6wEH+F
d5dpqOmH2I+YpqYxhn8wj3Y/8QUDadWjudc9QLLYG5RRUGdJMvbFtobadglFBAsL2V+rctOzhh9A
k0UhLi8kwxzOzaQ+X6L1w7w9U35Y38K3fMFEYaoq4Phjd8NcPbcZkgRDvs/7av1bCsmZW/vwcjR6
IT9dlHljFszZTfKKplDDLkloiFKi0aIhDM5xLqKhAFQdJnWTrwGmYZhZmuseUJN/gxF0el6Y4+Ly
VAOMuJiNIjKMuDuEyc+ckYXkjbna+nnzHvDPknCLNyQnh3SQWPOFX/gVVt0M/jTDR7C+HRFcRD3Q
jFLzn4e2nGxtf1GQTU7jVbv0fB97LTMlFdCby2ESa6I8RpTMVXaRfMKzAAUCwOZlCqOwXmpn+Vaw
UXLsOTmstaei0SYu4rKMk6jKijH5tfy+wwphW4YgSifvo2yYyYARtnmYc9ORpFyNapjmrl7yhk+9
DIT9jvA9hKpk7zKkgfKfcTNRsT+kTuxapUghdhUQOdn3zIWfO7mSoQe+5Q26QfURPDWGXqfERp0c
1oMZtoAy7PpfMLdImE0HIZSVa6gruZ7k3ApRHx243t590wAY5tIAMKln2rjhaYgrA0M7nDU6pG8k
5PoaT6S5xcutWJnLlLqQKTP4wxpu5GmlFM7g5l83Do/0LXv+P677xlrEhMKsHyHRcr6cT/gBlQnY
pfo4gP5b+FLAdaZFQPZLRq64nowljoy7s0EDbtHt01EfT4FPR0/jG2XSfOzzd+lj47BEMIXbJ6Ro
iiDOB+DRL1Ak/iGZCm1EXOI0PoR1VzMkBpoaqC1lBDN4Wt64g6XudCoLJoR1eG7EK2gZYbDX6poZ
xdU6BIRXyzTu4Ln1TULgsU2u859vS4n7rZxQ2vSiQrb3iesxpSQy8jIUSWkqtRDjJYexwfwaJGdX
ZnVjolvXT578vRTtBxqYFpnbMBOWSGjkXNCtEgGAeiRLmex06+QZmrbEhN0d4i6V9qk38HKgjht2
eAtH+Y3S4pDmPj1b6EP0hSidNge27hf1A2IYVVh1PfKYgURKJLDPnY2DaNWZ+XUdhg79uxmyxMqM
QH1mXWeUiqbvOogxKHReCWJBxKvTXmr3kcl13CMrv71zkiKRbACx34zENyTcYKqiE9re0Rhab9jq
U4pwKmuHb5hVkqOcpQhYRFgN2a1O1SCnJfhqr9bphW+QC3laEPCNZZAsv3PWkr6DfJcF/aYwvOIl
6rb1sMhUqkoLcr/6mXbt71X0303IYbj8L/NYkqAXr4RCptmXoVlIQRfSVftGoO+YngP6QxlE9LF0
Tg/JRn5CSUvilnviUPDhIi0hMd4f9oK/naA79n7pLI776qyvhKImQVzfNUtmyPbT9DUnsw12x+Hq
WXYszT/hS1NbkLpJE+lybMXKQ+PktMg+ArF7bBkFnZIkxS989RA18lfVVDFLx/WBNPFBlpgjxb32
TZ3Nok2tQivzvSB/4mbh7NRPjqK4vE+FSekkpOT/fuGC8qUPjrEmDLXndRXdQNamtz4vXvKKlylj
Md/BabXrbGw/64/mnik9qCwb0p524zl5+wRqaW+syAnZ+5YsaHojcmQJ0IyFXO9wGmeAqcoCa7CX
4qP4FIaFaBa+7nS97XQbeMtVwdGUyXKPFBGQJGaDKxVDUaFazThBiqpjwnD64JcRqj/W0BB9mlWU
ak954jX6hxjcotwFiWcaySlQFsTWrRKnsYkKjBkiPzg9Tjc1RQlqzRpHX6bbJD/ASkXpRFlVhFqX
dXWVDjtwLGY1pOZh96AiT+ftdezQ4Rn9iNigLSASkuzvsTXINjmEzTMc7HZL49xdEM31b6dyVApz
qCf/qMNzLPGz4vMPv6wtOSV14xUfreWUv2xd88/4VsNM+bJH3eYwuhiNEAkr7sutbOw1jofrCEg2
Wg0lbuGfqOw3+uXDirFFvMWT4Q4J/Y5PpfXzY4tamPE7wbuA9I1Td2lnZRTBIXq6vAXwmziLNBWZ
3VDhvsUSsfdCGrER+w8AIW1x7zI2YlTzZ5HefZJI5ajp7lG0VkzA9aQIZcYnmDsJJeyVAN77HyNt
oalrZfGnQ0g8hNjs8UvSMt2PXP6uJ45fpJFmWQkftJTp5o/YIw8dtN5lhCclg6R2CabQAbeb2URd
F9rHALL+sWZP+9VGXCLJGIfyLrzFy27AvS8iZo6/8RZatJxhBzLLH/GCmTp7h9Uml7O6zxC92Kas
FEOqMr1gCufUGvKH0BKRrEzNm2RZTci1D0Da9Y2pgwNaebwkdQknoi6x/39VU3snS/cx5HheORep
nnN95m4Z66i25uGSa7THzChXl1pGUKHStL/KjRZKg7x/76Y1DZVoh0t6ueGax+oy0zWY04/8qdep
5/tTjXGtfOf/dNKfu4kpzS3OBD9PKT+8v3iBaG9rnLYx8m8Rqe7vD9mWNgQEIvmXU3Bma1RvVXdp
zw7ucxLNIyH6911K1SSmdOT5+ivgNgstDCZ5AWr26CYHtkWjWAhwP5TgDIlfKxw5rTdm6VUa30UY
GxOs18AodvfvC70ayO8IN0iEpwWhAkTrYKHB41CS5BL1qKtQY3hLN1l1rNJJIKU8xEptDyal1piR
8O5OtCtvjAOCcFGDsn2QlRq/dJ964W/JgnfjWwPmtw1MSrs8RsOX3GMPbMnZZNvnKrW85hMAHo7l
hnjLMYHuI5BpdrzBsdbrmhl9k/NBB06uYjpIDZmMlO2ofz8ufxFH9+CThNBTo+W5ru0AAQV2JfTR
k4GrdhnfO9KRq1dF8lGwUT3svXuAQNlcKxL7pqvYWmU1OYzgCjYOqOLmx2JLb+cL65Ex6+Ckty7C
hi6jDPOKieQnlq2CxLaLJHwLr0Hbb955IX4hHm86UiSRVIQmRE2ugxncV/6CR7xsgznssdg+EyVZ
IGBrMf1gxY4zMeBB7KGEqJj0Zvwnabrh8HwUW1c4/I4ZZ5lsS4vO/kRzzUhVwXP0zqcfH/E0gV0G
94rsWSHxd3vIyYJQ6l5BPZ8h8qHckdK6ZLG8StehzhffZrdUt/9NDmXIFTayqrJhBb88IQDs0XsY
NQI0WDIkcgKKIKOiLSvnxGcX/XjC2DXx70d1dLKWdDQ+87Ub96LVgGZVj2frjoD5JwcG50sxjuF5
UjaCvmmQNNJ+uuQke3/WRLY+EMD0PtEg49YM7IQB0J8yxm2/zKcPJ3RtbyvqD4Ug8vH9ApQJ9O3c
nETKX79KMkftZ3e4EGdpNg9zyKmOjpouuW7RotYVKs9ZcUQA5h8frST/qqUbYjFGJVhe8REdf+2b
69sDW+MUS8xnuMkrRNvuaoXrOsD+Lq5ilpP7A2H62DWDd4CepiyUS++oVl86FSn2V+AlBDX4RFyQ
ntAfvuPLuRTiQdzZUELiwp7e00scegqutspn3fPIi1M9eO/LruoZy9BiykBJJPp2xBRCNb4xkG3i
FqPV+r1ooeBqqRYqgseuubm0sd4wfxzudWZ1f1V8RkoO45SntSNJ59wKo5pUBY9hBcYMFDoNUU0p
e+iDAz+fploCs6ve6Jj5uVMcQci+MRaKWTjDWFT8QZkhHIL8BbeeAp1Cf0iTqtdapnhZ9FUzQwGX
C+I70IYmLXzvGWnUKai7aJto9/lBaJndWgw3b4Oup/Po6ow56wYVgTDLEaSVwRrkm4IoTQ3wZdRg
fM4A10k3jZ3ohrqxN0EYFTk3W9lkc9aJAYKpAHGeSSGm6HEqExFXxodyXHXYgcgh9dsrYYQVmupl
ccO2G1y+UFW2wxubc0FbUbi3mfo5N9j/p9U96CX6jm8dAakRlZad8FFTiPtb2V4P4rPjvWaOlCME
B2qoLXgn6TlsNSHtAqzTVMo7SebvBpnxbxSM1vQbrc+v+3qxhWpIYvuO3VhYCSSZYzE3el99igRd
IA+eGfpdnybOFPmEUwSjsDGPRHaB5f2IDedQPpTPJgWNqF/iMG07Gc1QFUoVBg18C7xq8L2r0/ZQ
Nn4v1iayLSU2c46+yIRyP4+arOU0iM0wcjx9vTZR3zps8sTh3ZNtTz7xrqfDJQojsQXBp93QiqUZ
idYbg3GtkRiTvme7/xj0++DBmu19fb2oLvaAck7wlgxJsIyEn+gsm8fnDlsYqTtzmDRjS5xb/N/a
Vqq2XRahpdzH9sgp+NPcZh7D/RArVKFCFpQzn6tpgz7XdWBRKLq3iRb28z4o+xNcga2oceQjyRvv
Be3/BUbCFxDQ+b23gcwyk5wEclHGojY6X16i9GcdZ75QMXYPOcj3uiqjh7j+5vm5tHZZFKmhxoDv
eZjf+4q7wWkzJ5JbFFVrOzXy6a+YUHGCP8RF7MiH5YVYY7R0peLkLwf2u/pjhFGUhgkLw21rKgCe
oUVtYehU110Q4Y47l9D1JNvTt6/PEpluadMyT/zQ9LUYPJ1Jy3hHpYwC/4a7bzcRBmT7jNl/tPAq
haNmRWcQtocX8wLXa+XQfaowypazUWwJ7L/7HGARY1C7OQajKZHISAXGc7SFzlN964cmtNf4gfEP
ZodUKwq1NZmQLzY5/TNTprd0k+G80FDuaYVbC+0HcCw/rlnX6xYLJ2edE13A5Fsl2GrP3TkeK0Mm
D5fxHpu5lQtxu4sBoHwett33+MANeKdPMgN6dbuR+ugfj2lEyz2lyZdBqqppm4FlbpG8SMUUEnpQ
q/p5HiIRWiadkNsOVTCNmvfdT4HwhmBg5RBaY90Ua2uR4vH4+IOyD8wUEUn5Sms4d6Nq0vHr8KVa
h/YH2Xw+0Qaza1XjQfj/KzehCyB2/RVoKkSk+KTttBUkr/gCYZq0KD5Sd/Katocz6HSVxPiFItnh
zZmCnCEDzbD1wWBrzeA3Ysssw0FcZXOKhueCcwZS9IQzgiRDebWPomOO9n0qsRmH1inEXbaqUbhm
uxXVfPvUspk/DwZEnibRoEWj1rov22QFgE34llbT3i+UEZC7Lnb/jWSYQmR50qQra/z2TLDgfSye
SZ5kzPIqaaqj7U1pxTGQ+NWCcQ6FmMJ0KEENKrD51vHe3/3yPNL/pvrTDcwTgX4wBont5/FtBU2F
KHiKZTYq9XHk1v2s7jUYeS9YpZA6ljTqp6CNHi1dCmAshicRs25DGgmD0Zf9GAiNMNwolO5AN/rl
0KZH4dmIbh8kLFlhpL1DxM8rh+U3wswrdvlbJa68SVomwrRlJAlMly+5Y2cjeER1dF3Im0WdDXH+
/VmBV9GUdpZ4ed+4MIeiTwWVfnZIIWnHgollnPOm9SCqIPuN9zIm6oMVUt9O1m+h6H0Xh91+3Ij8
gUbF5qHTh2vQzjmwgtd4Q9tQKQMhQhYmqDOZ8SYNEJ2FM3s0Md/Bx+hspAZDunj+/h8paiPM7hIp
yT6WbuMIU3f7LC8JgPbcbigf+n4k3pgJ+BI5qw4f9OTkWC0jKKTE7FpjJwPLrPIA9Xo/OHD//tNZ
36CS10+H9QZPUorq2gRRmlvd8yMwUcEK/fVFa37FVVmVEciUmxOMascfMlx6ZEfPNt2pE1KeUsLH
8WZicXfzjIUhlCo06I5IRsAssyqdZX7yQtX0IipJR71TQMKMgXR3m2LT/GMHjK+aYe4URQu+Pkh/
BaAien4nH2RMcYFtCMI7bjor6WyCYFXKgtIRMIPmc94k8KoY0PTI693x2H4+Sdu8Oe+vG/zDuYNN
ZFvwonL9Bucv4oHEjOHqNHaJ5TjuPF1SwwmGqSUjCqA1umxrHChIdAwzqerRxwZTy9w2xetJH/Wv
buDVhv7Ym+mZveqt9fO6sDqxyBv2Sj/gIFDAo/6c21+lajjcqRDvrvwVEBfJRh/ykKQ7KsWrzuAQ
FKQE17avhGEXxqOuxCO2YEJJE409y+SQ30yghvTb1SCzKFBM03LoxaZPVdoxNKKOAVJV1JYdBs9E
sR2PM7NvESl5NI2Hw968qqhQKaN0cR5cdz0Du+vp3B6VzDsS8g3AKOlZaDrhrB730mVekOwc4RgR
jIDRXN+7oGXHSLSf+DhQzJ6hka/C7AadmrijdW6fzGLSkpzwxRcDk4Ei0bkuhTFe5ZbAS382gWoc
gXBApK7ODaOUWM2YR6UZPSymxwk6fIV/zqbggd3ao+kVuPMD+WWN5YXqTTeE9czBcN6X3So0pQOz
aiYv/RKt0O90msz+ZyoZwPQzh3suNFopOzG+HsqvnnScchjXW+NQFv9Vns7eDHZzjGV3MysDh6Uo
SsmEtnnvPq8wGZYOswJ1lCtqcmNuvrepwIpqPamaLtO4JLM2N2sOcwUe3vYyHslEQ2t42TAZq56A
/j+R+C6CADVf/G87r17E5C+RNsisGsw0+BjF3KzPblQbMhCYsqZu7g1gDLZpYvgla/KL45rMuBlt
A/RpPI0Q70+UageON5VKpQCzkNGX3aBvyzwvSz01omiIIfZYWFR1cN+HKGDzpuE0ppsFexw93aDm
49ZDyV36QxUhPVvS9A3kcBdryj4UyROOcmi1+O5C3b1P10xOJsB1pz7lc3IZ9afNjxu07M2xsXZi
U9JDAN2W4kXqQ2VuqPmPZRgixJQl0IyzcyuYfRrz2HmbdDG2za7Zkng0ttll/HZXzEoq9Woze+wh
BddhEVEkS1Bd1aT+LLIhiOVTHiTcC0rYJyy7v3bxB6DsEg7S3oCTcnue5obd+NdPKzIlxfVlDsM6
AWd8CAX+oYTO56ibNg6xBBYzZ4+B4rJaA/NKT+0SwTtnnd7YkHK1U/N3pjF7ZQDR7G2zoiUgAEOv
imPfMDSJoRRVOWhP71vVUiSLRPGKfotARC9TqCtA0uzGfXuSiOJysw12Bn6hgWhESIDts3uhpJvL
KHgfniVyRwGTz78uyTFsqc4Rlj4Txi2zlXNrciD+auopeiDQ9AJ6HMiv0NAnCIB20eY3cAjRC3iz
95B7O6U/njZge6prbpfN4cMia/XJyIwnjZ4CQ0kiqNZ/mEll8NwQU8d4yjjU/0dZFuS/z1Klzx4Q
4NSY9GrDjEfZLs4QWrTQLQn67oNjjk+diO+/jts0Qbtu2z0yiJazpXZN4FtQ68XKgdA9UXaoT//q
sB/SbTWyCXU4LBvfwLzrbt+tXynYhM/gGXeWXSsEC7lHq1swMFF9oJzkOK3gC6OruO0n6c0oHsGP
kDE70xcl0BcsBcsBxpPaqamnr+/nQ/e4/GtNAeSp56Ou4g98s6oUJ/pLfbikIurCkUmfSCO/DIAn
LF31+SBPVsNDq1mdwtOG8afL9sIff67G1octIT0vmTwweiMjOq1WTWXgr7UV2ICBkckYdfHakU7+
HF6TH8WOUr5hUg57bqKwI10PkUZw78VVl0+HxJ44c1e7rYen7vpvgjHFTtbWVJfaYlhe5ITlTU4T
rkfGjw/fPFRjIx2R1QNn5u2BCpBns7V+VBBXzpGoyaRFNDA9qA0OZhsCQZtmTIRTOSOsak1C+Qwm
AY+9AE3tc7BwG3XENWweS0YCUhVE4JuwSTiUlaOfx0zsUc2DoBYpxWqN3FDaC+j/g4VdeEvkyQUG
9yFsoSXnEhZHwAAJlyNuOxbXG4NVSVHhQtFNU2mpQyTHvIUisk4HWi04W29E1iD+chOwDlSpoLzO
Gax+Sf3Pbrxf+Zmdt/oXJocCzr0/q2jFGsKpUJP1+5uGV+reb2ua38JaiRJwlWLE/TODNO6le7i4
5NC6wHa+gnFIc4suhYC5GTouPVXdIusyONfUByvheM5aGlf8HPZTUYZXgGHN4qrMu7yRtgCBu88w
DQPmoLJPf20WTZ0GI0f2rBTlynP+j9JEId/4NY56wGm8Sfq+8uy/JtLWe1VQKh4D1oJ8GhaT10hH
x0EiGVN6o65ql9CVIP6jiJwCItu00IIhTi1p/dA4e5Shhhum35Og6DNw04eiad/V7eTB1CCbdMY/
4oJSlLuxhaxKWxKKcl2W8eImIA85i+UvRaGr9XuSoGbRv6Lqo7WJztVv9FeYLQcEug+j3fjZJ4P6
fN5KriMszqOc4uqMD3WIfQDYbSSbXiZIbpcfexNbxSGeVIR9KctMJYVHGdRuyVgNlUPfirbJp5Ya
2iEA9PFesaSpIJqXxb8+Yh5j/MBygU0ebGmHtY/lOChdmx/m68khSKZw1qtEYk6RlqxC0YGLY8Sw
cJN5XdVdkd8rgzzT7bFpQMvlgznvg231W/CazUokzjdjGC3RQVYBQVolUOuinq6w1dcAKyt9DFap
HUSk8KpTHWoCc5pd/c4gU0o6bTtbtv7m7xFdoYlPdB1sDt2mz9k6JHSCD/JsaBBlDrMlQVv+sIo0
DC2FR5ArQs1VdJHGlU4dggvYoUAle0Qd8vFVEACO9NEEC87mnzmqaxoDDc3FO9fF0G3bs47x5Hux
OSQq/EqANvA7n68o7aZUjGPVHGJ710BxuAES41z5eSqTy5HTgibKQFVrOhyGVcm5PgsPpw+NnLsj
XQlBO5zjiOKi3nQMlu/O/RW4ub89Z73EU2q7e3Wl77tiAPma/ZuAlPcod+FYfT8wFe30GlMy3Yk5
qeZGZXrKDyIBNdEhFzn91JT9/XSP1IPjhBI6eBoPTdE+3HQi60kCzTHu83sjB7maM3+GkQchYlOy
uTEbEbLDXv+X6qL/MErKbnBN24JI6evBGR/axNNwxI5jDpHGlj3Dokid1w9qXRr9239RJczhdnBk
L53YWFVFw/732VstV2UB+Og0Ee7ss0LzTdjCrNKbx6vLJRrKgUhWVV2Q5lN0mniEGfHL2utVzZVR
NKnBVqI6mZXBYV1bWhRSmDq6np+HBv+XpM6EBHmFlautEamBtr7pC1lgYZwSsKdh8n+POWK+j2nM
qI6Lc5tCc3ft290zEAhLQsfgZV6M9ndap7cvdEPWKtQtTmDyQ6GD1L6mg59yveeBhx0PvqFydb30
3J0iFOuducb6iqZzG3e+Be8S82I97vR+0A6knpdUaLQ9p3x5co5e6/47UzPhuVp/zhTB5xT5oqDu
Ygr35qAXn+3pfj5wwqeoGeojScI4HEAfjd3dcCIoi5O75G2Mx25v+ioo8HFYFi/7DHffnM8MaQFO
HtCc/F/XoleqnQhEfofyvs78a6QoJ8xua1zH5+IhRLx9KrX2KbreRzHe4MbXKsZovA3YNSPlzhee
bTTZtLafB5fsyjofKtzWwSJtChqnnXoUqSmfezxqdlmTN2f+Ks3Xue748321yDIR97rNS2n4SgHJ
j53CtBCX0FvtGwmocs+xj6ZWMUJripK3eTMwaIjcUDYcEJ/d2o44fC9oJWozjgxX00EK5SZLNvA5
rLgZ9XbjTBB/EyO4fdfaqwpLEr3BO176NaR6WA80OmF96BAtYGC/tayoS4hBtHSnrclDA3kz4I6w
FLNWZK7eJd12C4uFhcN9tm/J4XZhC4M3Iz1Y3REt11j3xdevHLCq22G5RPgWmozRDlO33bAa42Wd
wD0JKzCV5Sk//5HxflBMg2UwwCJRFW7N3OUnpipFJlM75a6XnbzhcZx/1+XkQfvLLEoYOewHvKY6
ARzCk/d0WqjyQDI2ji8LQ3F59UhUvybrDtBwt3A7wRecw0PWoJJzfyTzmn/e3SIYqh2F+3QYk2EO
PjQmx+LXN2yxEQ9tv1o1mNqFxi+nC4ZQf9bBxCyNruhpIFqwLffLfZinG8dna6qZGq11v04g5Ctt
5VYRwFioM6X/AGeEbR5SyaCn+Fxq4W6mX7vleo3SeLT+gJyGBEHeJsWmh1Xfi1aqXcNLEnwloj9S
LJA13skV3ervP2rafcI0vvV4hZuykxf4XnOAVEE5fmCl6ULBvLaKeGUKgQK52bu17ZkjExviGT3s
rCoX+TeXLVB/D9rSkmj0cv5j5F2ERz82ID5XpnxATBluOziSWQtXqE8FCvPwYT5tjBwx0qmTRBOl
4CcMnf0kmqnRw68rLl5CHkYEyeZe/6qVeSTBymHIIIfmYuy+LcvcDZpcVd5OeH9Xe0y4qP6byNxo
FxGyIVgCLvXQ7DQDZrTF4jomzQutVERsnKPUTEs8hlDiL/Uym7zwMXqYLfTO81f1NKyIuDXu1X4B
KqGt0utQ5KgylqiQI8B/xzSm240tucMRNJKncfD58M7niuCkY6zg1/E7r5ePr6XDZwSOUQescwC/
sDlCeQRaVCi2CTbIrtfHiN0PaAMRNmS67yAy0g+G4uMwSFGX4abEPf9kCrWlqwkrLFslFlyhnty9
qp5FDeKd7yoMkmMhXrXs8qnz3pq4OKprU8vOxwy+EC2tQzqYZuFrroCHGWdusdX6IBUDw1NTy1G4
u70ap6FkRw6iRNCXnFLsPx0kmsiDVXXtuN69kC+Wje2TGD23u/bpAy80638ivhJhX3/b9epy0WXj
IKa2OjCFBzWMouogwF23PT2NECpf08J7UwiRaSk9bNqoADMErUZI/N26Qslu1MECZ56aRQgyIrc4
yPTfDpEWzXacp5Ep8limOcwqpbLC8EIR/Sq/qJNmo0XQk2uu5UE1i60ybYRTE5hNSDnlWgz3Aqma
Phi5aOrQjqYESlc6PtIVV1NR3jzRbarRlrXX+LXgzKPzcojw+5f4SprKxLL4jwFOpXxkG8DF/v1+
dpXfEB7krIwk/dSDFkK3/gOddq0Bqh6vGQ6qy86vUQPKSbBgeI/8XjG+/7SqoPSOMWUl5C3Qa+gM
CFIY6afOELvcBjz8jXOESvDSZoiwcbReKLuC5oMPKEx0R6ov1yu8o35pqEE7NlvMZDukI/VI88px
pyLQDWJ+yCr9MjuC7kf3bdLmJ64m1zYX8BOWT8kvwMd7fP393ZaQFkSzjAbU39ukVVQAsofIw485
u8y3dDi5ObkMJEMGgbUcHDYPcQlhYFUuh678NhALRKB9/E4yPmh0y/xupPdAsGbtiear84zX3/Ey
6rkXByGyu5K7ZIE4mMUO6GCx/lMHqDgRR3V7E78HkpNsVmacRMjEx4IknUfkFFJyoctXviqa94vG
GeeorQ9NaRvkF8HXvOZ+ssTcMVVHwAj4r/RjctSIZnuEp+WNPoBKfQpIZg3zzdhNrw/g/4kMJ1nM
v98uRz2b5CFEdajkkWFD4X0X83ENX9pTJP6b10b5kSXcL7mupcgwZQVHx1+osGAJBS3uFWGvhhPH
VRpf2FHE6RJ23brysUdqRe7ceCwUNVMLbZ1+al5v6DzXwxSs+8znKPrACbu5T4rJHHiwD6EUQEHd
5p6G2krE0jW+yTfUs7gdhByKjCYjckWNj3tWquV1K+uRYYE4ZN4NSqvFuINPZVu5zry6J41DJNri
j9aDsD1A4rQHgz+mC1hNX5cYiTcmGImGSFZUa7C5du+miyc556szlyqsMtt/dDz7/aaZOemyGr3P
fIXuIf6sYSSfUL6d8AYb123nCHEAtpTDdLQzWUG9SB2v/B5k2kyJVbeV1iT0pQtozsLmXt8/IeQL
ruzyQQG70XmChoSANsWlR2Rk8KqOIgxUUU/tR4hwwpEG/IQJUoMT6zVUkViIZR4BlNQNKNDBAPXY
u9+ls8jeu3tfMcXphqLQl1MC116+FWYHZY+mkkcS01wKF/kLPKxxEvsOJcbUD898QIltGSepNOg0
JR/C5SNeW4yEJ1iD0Mz8kWpO11QWIakSQ1yM/5z6yYyA9hOQqQRnZyR4ntcCDDlPkrJQPOV5uW2/
QypZQi0zOjbNwJvUPdfd4UVoTM3LtxY5sBsFEDEfHWze4grOI/+OMd2Xt/4rwmSkk1QeUEDl/EQO
2/HWDTlcrMxiCF6RvmIGqM5cuSaxN6F1KdwP3qXG16guhAaOCWfcneF39z3DgnQc86Yz0R4rSl/U
SBZ48AdoJ9I3Jk2MM3V0A8uHz35kyLlsF/mVNG8swx6XwtA0lORf3Y9vw+MgWcrGDebzbBEE4kR1
nbMgn70XwxL81hPCjLhBoRIykFflooTYrWFPIb8SkC8WT+K0MZ40CDxzYccp9engPzt8LgipEKtg
F7kPfWWz8QxyRXUDEliXVJYdmQEqz0WMd5elGxJogKtITTMCbpGbA478aOXuth7VEEY6r3HxdvT7
OSWUCwofNXRveQIdH4uxoMMRhIHJ/ddLbyrM/ac8xrdadvUzpzwzY/sq08o1ZBSmlwyO8lYw6RRJ
atpwOav5f+iNmn3uOIs3R2ABv5jXvWr+OLc0kBLkk0S6Xg4OMeiRbziomiYZfjl/WcvwAT6edSUF
c0S8F8XhW+16A11aGK22HnUVrkjIlpX8Fed4GURvPuwY6pHRAmdTmt86+t0Y6gLx3YHzQK7Ay5Ze
RKJE8ceUgi6/F+/Wn4Bq3lL0DD33hT4pToLs2l7jQm6+urgBBcurCIJQKTywXdZqnyJ49Dukhh6q
7ncj3sYS60jwhxCwhz8/wlhJ+Di6rOGZIDKCu3gcReB6UusrrBPbig4IPuC19CekqvjCBeoBosJ6
DkF0vCOKUx6M28DVSqSY3QQf9guzUnNUkadkHIkZAU6CeMcqjGapbMKXbwEQW6GTU+KT//ioSjRh
TCTiJ/uyrYoxH/Shf+XXFnnQYhmnI1RuHZzdKuF8kTVhgmVY9VGK5diAmeGgPtRkEiR5sd+LHHju
vxm17zJSCvV2Kp9EFs0l8yCXqOkiua+lJBx6Zr6abfUhKnpSC5XdjJY9SJd6AR5g39j51K+MGeU3
RR1YR+tDY4VHMXz60y+488dZMoAfiGiclq5T46xuMF3VucnbpdUZddt9zzbTKxiYPvXzj4A3oqz5
FlhGn5N3qytPAM4F9xN6V5Qdk9ZLFSvzinethtZB23L8wrQDPj0NIy220VIL33mEE+nR6J3zz7BJ
cpKYq0XDWI3BkcVQP5Jd7fOyv7uavfnbA1jwWbxUxqhEQpVYfN7QRRxWqbHgotsRe3mckUEWqC6d
egT2e9u2XHw+Dt08SBAKyPQcGPdRVjRNcKBz6F2M+VxQJvl4+ws/o+Ozqq4sc7blOUjFF4eR3Vs+
NdytuZNrZ6N0Xn6dGOARuFss0pgYDFePlhpfzFA/G5BreJzF1GL2DYG+wNvEjCcUcmIYERMHP4eg
JO/B4N+6ghf2Lh7q5R6kKno2SmbuHKbrpVPxH/TTNKJ1ZdfiURK9appGbKZnCaiRXGOPn0otRR+2
RV0/ErNxMjVZ/Mnrjp6DL5r6rGhZq9r6fElFs81VDFlHd+ufKDYtRGprpRZZ6E2+c4am9FlCMF4k
1PxHRlZOKFOwkwqTG2e1R+VhY71BOyuF/XbgkdIOjELVjqR9HsV8AnNeeGmarcWlVGB5HYzZeRwt
B3ZPrlslJNNmhjDREw4bY6QbADyvmljWPRa9OiBhWuzUNdhoAadX7B7z7dIxaITUY3WjozOCrlFQ
+delPTgnR+F7s0wQWMHNdX3F9CnMW/0aSbyTrAMixcrcCwCM5Qqng0FFw1Q4CC+JbmcAt944QUij
mSbLe1ts5sOSgWQFu9+mS7YeWYUAcIR9KDl5A+vtft2XSsW+4Rr5bv4P6G6zeGIpt8WmJzBC7wgH
KuCIUd+kNXOaSpZlTBpw3QiRop1cgtqaXoNJdfCyxXj+IU3iIAv6zPubazVymeHu76GMZapsArRG
fLlwk07FfKOkZ8Anp6eWjgJCfGL2oOAFMgUVdeFkRuG0syLs1TB+ily6v6VVbEPS0fmeiv+cDLR3
xLWiSivMsor3bYTu6KBR8WsrLqC+Cc/xoJAMRAOw/WUWSXRbOi7lwK7xFbktXFvN8oAIZ+91UDqX
hZc9CySeJLMOQe7UW+UnaCqVH7TGlwvr5RNYl+uOe2Lg/tQAnRNi9nWOtRgYg4fw/Q7O5m/CmcxR
OWEJoI5jrUB/LeXWBunHfcDhGr0LxhVorwnXDk5BxV9W19bLk01ugU1ozfpC/wlx7m0Vp79sodJu
x1pjIPo2PnDTpDNLPJI/m0YO104zjh2jgfPAtWrDp4K0Hox3EYxveF62pTG+kZ1o5S7Nepd5TbAR
dgueNJjyO2sIobs8MHFbDbvkMaqXq8c111AyOcMwlFBkkbWZd0COjdo5NktBd+KwfoJ/99jgRckK
1pathHyLmcGsue/6IARfAYHU7Xj4s75764Losup2hYYDhbyUkkxa+6C5w6MMsP+79gduS2LRgCbx
YMGdENAAZXv/6WvxtlRdB1n108EWfiHxq/x7EvgXtnKBWC3SJix3YbvSAmn5Ae31+oiJDWpzcyE8
ERcU39m4WBzDKlBO7Y5cG1036LZFBhlVc6h73jFt5ZlWkNVJKWU0ZBtWcTPm+ItkaFnsTXs/6OhM
XuvCOE4yDvWln12zjwthFvXwi+8LpaxNn09lgzx1NJGBZpoW34xelSSbZxb2iTdoi7nYIw5oDVRJ
lWsgGgLGRwF89PAdDOJZ/AYGupbfgx1am98J4sUaw3li5bwNH3AFa/uSTM4VU+/zuD9UfIfm+Dhw
woiD3uvcSgd6MIu7fCVxzjhldcIk1ZwRk86Mx8vFC2RvF76NOozEpCvMVObFAbCL5WO44OTTod2i
4wrg+4t4RqgRpHU/k9JtCX4tdHOaIEg44La6rJJI2/PEuezrRSjDCLf2NoWzzNm05zk1z4Kh/Zc3
tCeOE5mz9llGpv5lOvWuM5QHsM9Zkmz4bSXNEEOWPDnMHalvhCe3NynWLjpmOa4TRvkKkrHiDX4I
hZ5b36IvryCTaWYcggVB5lqaYdNX3WjJL/nvgA+d8dV9BHCro9jtTwsQRda5VqZ6Ip/SanCr89Ih
MW203KTtM4ezwI3Mwf3ChknDtJcIJPyJZzaqvdfKJCxPG3w8sVSc60rIgU3h2/ZRVRhPIiM87AVH
llydwObvO+x0/BDkPLNFpnPW+WeaJ1kVTwdrQg6nd9VED4QHKcqAmJBbGjdUzAi3VYsCqQOvI/pF
5vcGvkTgM0iyK4ZQ8CqKMZcAKZaYb6LmXp0qfGoFJQCzs7a7s3icP78RIooljIh5jKLLf5UTDzy9
iEfonBxrO6yimGjJiz6AF3HPVGkp+MlYO2xsBPRE+cxEQzPupsDPzb4xKhOr/j2do2pRcp/8yFKc
cugSlRjnvyKvj1RP2qd9LRUXK4XYD0VaMce2surPnsWhkATelwe+uX10J4j3ih43WpcBKEONitZ+
/JDQPRC2KE5x4YLBSzTpF3cwK2TvFVsp9NRnSG3MoNXh0dNB8NxzC4iIqNSqKpCjdjoejae0Gtva
MgfVX2sja2RZPX6RGzvX9uLAttimRvr2pSoD89Ji3JD/bDwOU8JgHovBI/EAb3MqoQyGroP/gZ0t
KIf1r5cmF0ydWK3Yu6n7irTUugoRWVELY4YfNI+m0WHSc0WtQZJcZi6XV33OARD1S0Hl6OWlY0KK
MuA++7Xtbx6ps8zkeuMi51qzTf6sp5OPVY9Iqnl3wc6syIHOA9BRivoWtzrMx7i6gF/0mJqJq0r6
dEtOcmfQBCmACW8T2KkRWSQ3YOs1EhORbzdWme8ahOk+Ra2GXYevb0irDDWlwppHCexa9GhSO62g
5QgDba9OyNM2Ujgu7MX58tkSZ6NBZhEutMNJeVw5+dKyHsNJGToIpKLLSU32/ybQd40mLktduOpe
2w07XpHSY5jgM6MdlGy/b+D9BDc7NbufgIPYAHQ5GvHfiB5CKX8WbVBgVpS9+LUzx0DE4G8Ivng0
2k+isxexoME2V9p13G4vdT3kD3UaBaVXxTGOhYoLMY7kRqYWrq1RDS0Ur+dt2tMRqJhtch6t1U70
0axXGhTxOoVBNFZGy5lwf+Zkth+QJ5wUgqBtLZrflC6uvZarh2lJqSe/WypgacWSdDwDFCksGr1d
38Ll937KE5h7185WEJUs9bZcXPsQS6RkVAvDIwfHeN9PFfDU0YjlaYke6XTrJpNaSjxxSYkdtwpn
p1S57SuKVGvbaG/PuX9fgwUJON2LkgwmejEwQ38ynblm3Qne9VhrCYVaFyGrRaNGNgxbgwO9IaXX
zl+UVLxXdkzUcQpVGX+B8gBYfVmhN+jtMWFwpTxlDTeMgCP3KNlZtZtA0Yi0qzAdAocIJAc9UprX
7Ljy3/ihlNjaINi0FNGjPgawWNGEJqvOna8ocrJUMcFNl61JACOiljHAYch2W9cDi/1SUyrB0gwk
x68sib8nhCDUs2dvGSv2AowRP+RRQUgpYy9HMVhySrC2ISfTPau8vhUyZxmi/ZD8UTukopyr85yN
zEtAKz+PhDiUn/NByNajY1BRU43g1tdfcV5x7mubHBSmsPfh5AGLp0oB6lvLeO1dmAXhMhiZJ5Ro
Mg/5EhBfXZyAa/FhczuBAhETHrLLTIgHZA75zLjLxoTSa7usKO0xywB91PHaWbZYa9i55SZU1D1W
BPKn6Bx5WhsHDTu/i6A/xNla42PLLedunVy0m/lJqfvA85lwX8h8eWnVCgF/KHgl9/ciG4VmiU09
6/JM3QBAVEtqChZfY9p/IZhFQB3ye5DKaU57qhCuH0YEH6FNYf2umHnmUm9SqoTp/6Wiwg08aOHv
0WckzEO3qf4L/WPgrtIEo1Snur2VmNgUtsBl5Baj9ubAc41pOk4/rBP4iGL4rEgsnp4iy8GLc8Qo
eYxtsiFKlDGazvsIFBSDnH0Qmm03X5Y7JzctlW7ke3crUEYldNFVJjo3ojRTEaC58RN3fvyz6dnv
xouPhdPRDU69uB9AJHkDw1BWqyn/u51EPWiGw3hdcb/ESgxkioamq9racjE551MVGfRAQMW5oRiz
ECtfad0aneq/ucGFmDGE+DxVthrXL2hyiGGwHJb3ferfixQW9WAJS7WM2VABByt0EgiegNSYgpoT
b3RYcAn9dELjTRT0cIzzvysFohqH5yRJF9SBUS7sBx4qWm0RDc1YKls5cVyLFEV59bZ/LxaQX5GU
5TmMc8g7kJaMMpwljx7ivTUqIpA7SIDl1ZjDWlNqe+hiWVC84GtSxCVgvlWuijDJcJ6n3hd76KdK
X05EvaUQCxa3aUa97CG76/SzYOZQConBwwDUqC5O/0cimHChYdvQ3vTJpm+ZjtZam76NThM5seuR
7vLYTROH797TvzA/mKLmibcs15v0oNGPIWSUTWmDTsdJM0ik0gCuvbOTpp/i2I7bngrhfInrlkmi
GYBSnKjY1SxgcY1gqOUfEKCjK9iSlFqQiT4Q6tYW3420r80aW0lbfgIRhWjAuILfk6wn8XFmM/tK
qemZpoHwajOjeEv9HeR4BP9zzdulHloS5+5OG9gWOdq+85+Ts10ZEB4MYIQW1ZV/rFQ52iczTCLk
mXLJcVnR3P+v69Rl2ApHpG7//sALwJNZACqed+ne3yHRz8RWLij3WgNHZKsHlGPlxTQY3EdyhPGE
Xc4WEk6nW8FAGcIlFRAx/kbwltTBZr+KaZdVBHqCuCDZ9VhhRbTH2pO7i3nXVfnkH7Lvf8PS8UR1
ZfKRyDQpNcfvVXlUU3X/OvC6+TvnOkmmMv4GJUlDLv9+GmXho1DWHvJ4wRFgJ6w9WGcbEJNCqto7
cFmIYou81tFwlGwbxThq8efc4UTjO+fx0TxT85Wf3mpDRKWRCt20+lRKmJehKPOvgFPhnMUWHMB3
a0qeFxPZy8w6xE2WevdDyMjXWf5463Qu08fzOftgH9jLRLzUvRvCBCqSqdmKHDARQEGghMOTn749
LK1nJaJ7OqhcIv4gm/lYF4QY5vDU48yBCTGtHPfjWHi/hXQ99xJWP5/MqP7LGtOmBMm2o7qosIsE
B1yVCMeRGsnrQdBpSDyOAMqqQa/+VY67dH6eNde9vlaeYVW31Fi4pq+WOwo4GkNpkRSvVyogclQl
ddbc53aBccFxP025SWlfbTZ7ixEdjSKKc+xz8b3VK1cNLemGfGyJmRx/EFbKLCu+C5akLGLGwunx
lr3W1ISCA9AKQHPXS9/JbKRqSDkb2rgUl7d9PHZeHxkIxB35+WDGpQXCHJ9YLoMDpX0b/GkE/2Sl
z5bXDfcmSIcWNgx7XkKQDXSyg20IaGy6HZIJZkZ+gAej18yp3qo2VzoI1QBlEQarx7uHzP/M2wwj
wLlf/NpRmsI5ZwZExkXQ9Zd9d+OKMD2Q5H4srZyU3crakTTuaNfDbfq0lrEVTQ+siWN4QkV+/YxT
/ZyCCr7RQUwemFuyZfOBG7+CxlXN6YLGoSOXAjDSdexLxtSbiBjwYZ/KWB/Y2/tavboFPtq1VtDa
muegq46S57vNTu/89o6XR9lQvPeRaoEejZEGPSToAcTXtsBIY42dUJyhJdNwoupC78dXmWFAalTX
zsDnjSNEhSV0Hp9DLqCoIlIsuw4PoCMv9iZNBgo0dGcR7wr3Gve7l/PFAusRoR7egAySJMM6rKQ4
Wt5SVzcZ/MyWj+yWMxKFG66xV4F5wO71A8P37J2SIAp+RHMZU/Pcj640sb5r1nhgR/Nl8FC/KHdm
bM/4admIVFpcBhWm8+WgeY1sqLq11Q5mRgWtiVKYSiFOndnHr6TRJVCfK+Kdzx0nsiAv/Nb+0vWP
5hmv8bBTzllkrzGq+h7fkiYEp3BAY19KCGUi1PI6rgNSQcl8QvXEsES+5yOyyY5/euHchfDEWUMH
y23Kh0k356JCuAF5AmEuoFZQEHbO7bMHEn+Ri+pYvQ3TzD48Ei/aPG746XHYmyT7cyMr5xYTUnhI
pknYO58vOHHTG1i/Pm68/C8bfLXNhoKpiP3ldzsXHAG9AbEF2tTFAtP/65AU22lKTPvLd+sp35Sb
VS0Os/V+KdojImz3IlJ7Ubvs8IR/kP3wF5XqJi1KZiyXwk/BzuvTIC2ALBzZtGBJBAVe5NhT6AGm
11qr1Ns80X6Nq4f6Jadm4AMQSg1sNsJIkfMPiZxQfoA3JT+REEtdPKeO8i2MqbvK/n+PHnJdZ3R9
5TZ/XEc+9IspRJCDsCfoQ/CROXPIPjveqr4VQfL3WMQLgR3RVBhW9/Q44aPN2uFXQ2PFGNx3eMRP
unBpIl5N3JDKqBeM5/kJCWkjgHYNnrUa9KklRjYr5yLjiM7hUMWoEuFMYbYsfC9Y+b2ZjCgLhHos
Si8F13cA/YjjZsrGzknOTrBw2/67TyX/vEGKrXm+tmf4GANqEkwaMin3GtZvnAHXkRBvzoUiUFfu
2f8nM4DO1b7Aac6l7QK6v0XVPtU4mMGTzNytjzhU5Y4Imf2dhjY2sTZ5AuUyXamLw77RM6ayiYnN
vJ6oGCVpK6iD4+SRgm7eSBV7RiHmcx4qtqIiVnhiAjcQgqR2kNnYX500apHTKNIUXfT+POrtc8DF
KBdvonHdRgfVSQ+fYw5Yp3/9s8hniJOKMxi/W6pU6/Nbfd1+n4NO0syxkOi151mj3Qd6r2RwV7FL
Qt0aJXumxWW5Z0HDpRpQrSvnQQaM3u8jVEm52eJeyn2unby01jVC1syEbgMW5BFQoHl3TGnOdhmi
Yz0qcM/i/qy1oYQbo5GitzH8a3j+ssyEzBpZkXl5yKw7yBUWRWbrikQ3S8TeuZFzZNyFUbG2APMw
iay7g9BQos9O8jS9cy+V20NiK50upoH2qyK52hmVqUn9cRYuEKISCTyRA29Z9siUjKYa17+Fwqs1
EE8RjwsmIJtRfJKX8EIIWURukmwHoQ3Y7S9Ro4GCuw4rVAbgU0NNNI+rYCLnJrOPNY73iqCkVhgV
JyYYWmtTWnQVtJdvy6R6JUEiMh2zhSoALw2jLkamxAeetXVlQyofZU5jBkdtlgCwQSmHY8EYgTao
inT/Ezlsbkz1FV8YCknaoUSrioULXNco4sikgrnsvkU96CJBkv73yZxG1XzNMXx/c0VHwmzDZ/mz
lvANbqVgrHhN6YwGApvelmxUQCQM9EzHWqk3MjzJu4/P+ekJj/WNJ67SJ0ozZ8AfmkzNqY7qSCHY
dQ2O4PWZ7/9Vp7kgUonOIADRgDBpPPHHvI3UgKbnvRTnUXEl8HiR+piQvDR3hbvL+h6J3L7p+PfH
0pJO+49b50t+GItDRemkzzTrWOAPuJWB9lQkpPtMZleCcLXmT2zUGW5fyaB4/JVZDIsHIBJbc63e
/ZAYF5uI0JgHd9IUOzAITOIIgQ9uITTKMNXfeVCt5Fi/yy9D12u5nS9/Ma/zulpLLRuv1t2CWDz5
E4rxf4/T2MZH848a54xXJ6M4XxZDQO1M4e3t129hUeBTB905uDoNn+Prq6PTHgNjUUVIpn/PQKzG
SAhnTaqQQUhu5YEHhVY2euVNV8xJBPjwE9MK4C2B8I0jB0NcMOWjvljvHQfe0gWoJUe8ZQFMIsl/
lO01fE+FuD8MBgMZDIvS3N5AiWyFCTAaeSNCp6jue2Y5ZFkOEvViFsis+krizTRauE5OwBs/wG9q
R2ZPF62nvN0cMzr5bXnlMBQz2jkLKv5ddIG4ixF74uFLfnHNXzTp+AMnfl2cz4ofJvW7OSF58I+7
Va7mcAuqGR2+L2e4BvVT+KTbcInU1czaxLAKg7LU6inqlq7jqkINL7jYI7XeCQZzVT4vUxNzQt56
SmrUgYCj/l0K5wXdK0ScgIy5eyrkjfn2kY98K06Dvp35Oh03moRYg045Y1c1zjqlf0VmCXviIFrl
fgDnRsrFZNrcvxHJa4ZYuY6I0VCDsV0JQJW/htgM0ouJst/crmlLTNY570hRRH0qR8BKPQglJcNU
6Ff34K6Qnwbr9Uz266m/gNgW0tUSTJ+Xs/m/i4dAUO1quG8b/eLzZbSDDxE5mowSaUfRTfx0j8Sh
PDre18agFToLztVZNEj1FT+z/ghYLvmuK1YchGvoZrqfebgzTVzPBUhOfBcKutjadpQXYDPrTwWT
njXlqUqfvexZPXg/WhsdyGkSBTECHAyJCo6+adTV7ByRqB9YpLUzAJbYg7hgCJmpsoz8MH9yThRy
+pyUiswH0cGV7/4ym4q6Ol7bc+gfZrm5DGAZj1LH6iP2jhgRxGX2psjdn63cNUBwr8araTz1SWUs
h9SPhDJG+5dDZ/lsGhK0yRqk5k2kXRhxFPi+7NShw2lHVWAm+MXSYu4WTub0ZAtY210alwofouHp
irImpDVOzY2Ga7/61yU/oX8y9+q9IV2bJlC8KlayBYh5aO7q+93moUJ1MKIz6cnPUiOkPpdeLmLV
AGPijbkOuoBTx/jzB18xUKA7fb+fbqUEuHIvcD51itR9807H0yHozoM+/0lZb2KrmW5lHf3yD2ry
VB7BjPFL/zKhG0RO0fj7/2V3BBttbRh0nCGW6upCl6X0kAJ8ZitSzrXGyVjynIrOGjO2fG0V3arf
gSBt4S11kUh3u/9vLjNPimQJt6hMJTRDFiLs4BVBvntRRI4n1waRnl1dOQWipl5AXPWN/vWw8pmQ
I1TFWxFBnQxIt9z6aM0BGcfNpNMd7Uat5re0MMIl5wENHGbkP1yoUITxImAMKIwtdZGKD5dwR612
zck8PWsVPCbr85S5mADgjO3XzEhD95UozqMnYSsEsjys3sSnA5mSSO/3tI6hu5e5I5/lW2AzNeu/
6ze6FK8H/vPrk+0GuMIgVX2rKWQecq0EV9QMnCOfisKzFx+LWzOs289tKhq03EmCdvetLk8nfRwQ
QVFv1o7MELQTqCFrgTBunbCbH8t3O4bpmfHRvOs3QTYIC0dzZquwYLAei2v7AW20dzbxBwuEyaj/
+8VzmXp2m2CzGJicWqMSw2fZP6gYrh4r0+CDrEuT0tQRNKRhPu8utK7lf+B3CzgUIpusBpriBVEd
TwdXxZlH4TWgGPmt6zwBD9rFynu0OldxOSQlfJpKyCSKKrWVATPfdxufo4wYxyPJt5ziYEJ1Z73S
LRvnmmkINnHovEesj9JOe2U3bjAR/E87GE57wQf/E0kpLEh9yUlE0mG9rUT/T64dfVLv9lJobk3a
p3Q0Ds6skpnZAhu3YY6j084CjC6XKrnZyCxuLu10lfwwjlAOUcBh1InLSWl0uhqsBS0vbOaZSLDk
HQCD/Lh24kWiUaTDInPhSYOTY+VUjx7FiMyTWGixeRQvyQHX6wPTZk1N3WldM2nnRS0XqqBx6hwp
+cryWzqv0ArO4L//XbhHU+QGcehEp5nOnC5eWoLC8xsdM8visRbbx8XGhfZ/hpqYGglJqohy8Zg3
It7Dkp3PAkX16EFBjDhvRuw+6XHGskkdmAbv5Y6vaN79bBGgIttbP3EDlh6DZIiLzHXXaS8Ncsqz
Flmi1HrT2VdHR3DHdpVkBiOunebr3Rt8sVDaThzdX19GRMeelxaBLv/b/+/GtkOKnIOzT563gIKK
bn8kZrWP57+S39tTNpCMEvMj9w35WrTjV88MRvZqd390TRhG43t1cvSZ2sHkiP92Zt2HD/+Zq7YM
59DaAPXjZ5e2mHbbNOAPhvkWbQp+pIuZ1JbnuxpYtkG8DPGPNMdvPxKRP3ON5BRALFPvo2sZC2mG
GUW3sBgtjGCIfrBISYEvtUvPQy115Yjw1FfNrbRSKoT02brnfpjC2PFz9cQ4TdOo/a+AjLKBxk1R
KiA0/TpuYDe0ZPNJmW1rMC9bG/3YyaSUzG/HGfPjaHzVUz5wfuA8BhwVFC3owYhMGPlU2YkapJ+8
bFxI5S2ISmPt9Npaz8nHxLUc5TawiN4YSk94+FsWIFfhpjca8uWODs8cGORCjq4txrz980ajYoqw
FoAYNYbEcK2J5Cp1BGwyUMEE3Ms7FGxiXE3kyXqS6kExoNO8etlRERAjIhJMdgOhjgTRXqRUFfM9
p2tmGv50sN0sfYeUlnaB/4qO2JfE5cT8uXWTgtY5zjuzTmNqCkd9q7IRb6nH4jZPmkNDMPHGUvFj
xUK9JIFf/VA7zaFoe/J15L31b34AlZmchmNT6vNMpbRcgZ+CMgxp4FB1wIpd1/jWu/43rD3zm8RV
yViJ/63EGIvQM4vXhFUd5fs+12Sb7/gAEDZEa8EC8Iu6FBMudmGOCiBtpNf5ooV5NO6GOdOfQeQp
URjQKpvF7XUK78twEZ3C3PQ1+8UXscw84n/Sy4xGHM7gt9Js/OG2pUHCDBLzGDT4Q1XdbbgloD/F
HCCeIQ6A1PU1FBhxZjz/fyJRm0nhV8L2nEW/ylMw3QQaawJQfC40M938kuBWeIR2YSzaD1qCCvRl
3yDSUYTSXrMKTwubg2fNFCUG9Bgg2Ilrt9wtwdkTna2PNoXIp83gZvFFiYXZc643qkvErP3D4qQs
iOyBnmjvI1n6XrR2PWd3JbGCkCvXxR/Fu4PxytRCumoT9r7y1n2e7fDuP+My/Am7qjsc6HwIz0Eo
mx4HD+mJvrlu4REPm4GNqoh2BdtkTp+FRtvacvqcfvBUQLWzXc/zwl4izdTqGw7gHZ8Tp4/NlxOl
z5ms/lJ2GbSTwEij3MZnkwOlgZQTVAXrnhUrlO9jcgZbT/t1MLtjo2DjcZ3kRknN8XL3duBb50Jt
H1yiT8K+plOyQM0i2pqXq62riZbZD4Nb6ZE8THXcO+bdZUtLghY+89u7t+r3DtJlZKQTbjN+pc0K
bX+Evp5xu6zn36Rmjd0GavYKc2Zhh11AIYsNgbUXY+samZI5iH+Hc4HVqUKVa/w28svZv1s9rj76
i+9cRLZ45/UfxaIUIGI+BI9BaslUMklx6E8uzr5YE35ySL292nxeqnftky7XJpwdBsMzNXz9lE/8
HdafMOEy8byV96vcbi/t6/bNtfGog+CeGSRnJbMFYmQUpKog1JUOuy7b8h+kjoFsSzWraWJMYn/m
MREfeOe8RLflCVFBOs9mC+lalNYGvuBx49JEqeObR5APi+/EzU+UdiDW7QCIM1U/+w8B3ttUgxVM
XWpEsis9fFv7zP9hYcFROS5ahnI6LVd9vGsQsgSP0nfUqY6CaMC76O0DELa0QI2MccYd5MR4WI8X
TG4atkD/rX/5RuAt/EgD80tPHqgpxNWXg3vDV2c22gf6LbQFi1AZDrUWl/cczQpgksdAmRldu4Fs
c4tnu/w+TnyV2BAotlJktMxEGn+GjCOITIie9o5vtGeIzRjbMevhbvE0ugFrVk6SwrxUxwR9QSAU
h2gkYznOomAN4LBhvQjJkYBv6Y3DN1aw0r4e2BnZPsGn7rbsA/LMtjG7AOrDoHt4R340/6hSh8J6
yAXYX+ubjtfhk6Tjblw20eEl5iIZwAy/aMsdmHZ+EWYfokE6z0+fl5QZ/uqCVSJ3sib67Aj9mDxP
X9AQI1UZSupxsXvvPvwa0YekwIh7NJQseV2i6wpKxBsHa4iDrzf3RNEnd3M1dzifpz1i/Wunjgrl
MN1ToFwlnjq7nChiQ9T1kAqM+itgg7YPa5hmYoJCarfGQx5tdpCuRXBOYEpjKXmIINvVg4rFqPGU
4rTLCjiIlgWr+Ld/uYOWcBrhLoTdpFmiK3tuHaC4UM+4mdU4Nn6ASjSEga2GOT6G3vzxWa5PHTbk
nto856GO62wcIWD1UKDAkylViKmmEBSCyeSZK0F9fhCsL3Tn0rjkOJKLzAb/cz8AJOKWTE5xvztO
DO9eQw+oYVDUXeLaMdpJkb3Xs1LOs64eORLHA1U6o2vlCmH/8FSpjSuc6Ev8in2R/bdpfzFwrMjn
PSx25KqPWdxMlqmdU2iKS7fZ20mFjbWlQsYbynY8CVkDQ9UBv29cOMHAMwaUNtZv86/7bnNBqZ8A
gNt08y8+NFMUFsMzlaI2f4+tX0t9uWT60WS4dMW7T2cinYrh2otQPawS2uMIgy6ZE+ypmt+FwqbO
p1IQKNy32o1Qf8SnEmV1lu3ApIlTwt0L0Zz8XUL5Exly0je7zN/HfqCrzNVuC7SPuMeDBwsJkxjh
8m6aTax04M/GpNEvHPb014ErhWqXx3EGn3i54GKIJE2UjB/BwzBLEle4tX5vibtlEYLypQGmc2q0
5+Xh9Wk5/OyVME4DNu3UMGYZnP+Iq63Da25zyF1oWAIHe+6S3tKkPkS9esGsz0AxCSD8X1X0Gs6y
FITn3ATqyZV37Yggpvfvb7DBNdmHAzP+F8HTSweo/YWhrQG7xP9bM5l1Lzn/HQIHR8LLeySGeg+I
ph3Ny+6rDfykAwV5oKoqSVQOpK2bjsqC1/qZwDtJrq8peL1157ZjRu3K8SThszpwlkMyJvAt4VyZ
nldDI8kv5Gkl2gzZtI/HzysknzN/q2JdAPnbcEoPf6QN8YMtdC/uuMjkk9WvRc58YmH7O2Q9bQF7
ezUf04GNtezH02TH8vj96qIZeX+WnIbS04x1SGJfxmsdXOmNoUydJVujeNRyW45/0lqtX+nNze4Z
jIa8KqJFrLKC8xqoWIuvyae3jlZzJzQF3SCefUNQXq2657Hfm7h/wZhgYdxMdQUXhJqqENS6E4d0
n4kHAF7AHQhTY9LyXGF+EnUDGjlHzuYEN8yP2Ar4VTZZLW+EWGQl/mXwth327eT7OHx4InLPNAIb
vqvGmS0jYA49gQUGkWT3lHA7JX//xoh9IJa635Hyb2MGuQyaT7Fl57HGvZnjo17oC4+950UI+sX5
d8Q9kA1TeQ+uf69P0uXngxYza5fswOV/g6AM+rbt5dOevzT7CQj+2Gs9ASHAkcEiEgwU5WDuTwQg
kK8mioW/FyLsjpM3JRQBFBH1mPJu0BgQsHGXRF8frp0y0B3MzFwluJD63OZBZPQD7Un8H7/U0zVj
HDQKQtX9KLH/KlFMZZCxuR7nuOuYCuhhlMbIcRZ5wqLsJbawJ05hXUxNTGmMucZ6lEBvbX4rXj3Z
05FBpCw39YxTnaVXtbksJISaP/chsvZ3azyV65yO6Ly0W4/85S3iXeA0FksgLSZwlw/zUSOYFu7/
QvZH1jfE/JUhmKC7UbV207Fc0i7VYsBp1cpjpqNwsiV4eSL5mjrYk4YMMyBZi5u46fqfiOGuMBri
Fzuod3ZUafiwpx/xFRPJqI2ofgXe/aJLHF9eHAU1lmnrUmFsMRHxVb2hE0xxtt1Qt8ZpGW4JA23Z
NGWQNjJ8TqPQQryE+uAcJuq5jqf9Mxt2H0oT51cRHf9a2evk1qpws2QzA9vWl3fm6/62n0lCqh9X
OIpwCig0UuZAQZUBUsCw1pLmU+//fa7p4Jy58w5poVFqbL6Hy5QYkfhBTNEybaY3X0X+XMsHKlSA
tbitezkGXmu3sNDX+hI/lJKflbPXJO43/cfOxfDh3DGG/vlIq4xsllmokIMmrwYdiI0E5YSfciC0
Q9iEWPsYddNEoD/8ADlziPiq+SKhgUBi2FNEqAnfJBDMndZcy97kbEkJFyqTKLgkPLt6LTl7+pDV
oZMuxp8VVQkKDOVv093xPqzCQ5g8XShaooPLNRPp2LISIx54R0OxuG2a5lEzH213NIDQG0XJ450R
BHogtuIYILt4wucTedASRQ+zHI9ipFSt4RLg8If0S4Ny97itUpdPHkk6hnyb5KrUYOOYlGeZB6XB
zBEvOlgyaH4A06pQDc3eGgL3tidsLLFijfmldx32WEO9ZDLsQ9eRQah2eraMpQO90wPQ7+WSjNoP
M/nOY+kNdLo5dpQhHWo61+j3cZldZGFYevAyaO7ZB8b/aNhzrQUD7GgnBu/Blq4dxC/YRwpL09Ak
glDqnA/MFXy3Cf8YLUq1WfE3HNCa+OMLacZiuXWi/wssEjopP1dbidP+E2u8H26ZHww2sGoMuX7r
5lrnNa1AJM/pNeVk2AMmLInXn4VJCwR5RsAueEivX/8kvy2Jnpyt2nUBCylgwxF0yalThjwUoJY9
MgSXRH0kO9arPNv2vsvctkEgQv/1zaa5BhoB3Dp0Oy98fDf3jhBt4Y3dj2UZ7IY1dx71tLkQasM/
oGcJbGRYICAHR3nDrsE0opLr6gxJuICfyyMzoKtHqg8LCVZze6GXes8tjd83VBt7iYhQ7HcxML7/
jHQZHQdSBY179sC3gDpVH0WkntlICp7KSJZTFH+XOr9/8DH1rBJPCBWVPWI7BHweoPf96BEaHP/8
S/4c2QoNBGEIqIQdEErWAMhEffjPEnhy2j8X1UlFW6wyrOTgfLAEuN6eXwM7vUM0Yl+cD1NL1zxG
Jp08PJoU/rLXSJ6IFhcpiiZMA2IWSa3FDskdYVMIyx2LlvP4TPHRSo75k62KukmIggh4JRQZKXLi
1sf9zi2JPfli7z1jFlqfklVG20zOaJOxIqNyIUO8qD7nzUZrsF3FJFx6gUI57Ujs5cDZxphcfhgY
IeT7F3NcXmfvNiWE+lw31W9EIXLqUDYx+kqKeVlwu09/fInkl+qkWFfboXNZ/ZbHX83647vQ02nE
AmUXKCQk29MYUMAzUn5WDIGHMEHcAa+340MdSL5rMJBYjqcIDHZp4UISM6QC2EW96o0xP/DFCHQn
TRjlclzzTVGnsubBVLgNwyuwEwr/3VBo+P7P0z4Z1XsxT718PZErXq0dkNTacwdqA3XrIbOozL2N
jnY5nzYVua5EEOLTyE9ZifW4IG53jAUbPKj5zsgQIEcuX6ZO2E/+fRTDGu8QPS8oErzcI6WeXeO8
tQU0cchnrW2ZTmButcjrgmL7nJAc0l+Q1yiPDI1kKi7QmA+jSPbHXh7iqzquCnln3Tu7zsj4Gvm2
Hwk9toRfC4yPKQJ44NIfTDnnVUUEKf6cucYqlq0d1VUzPK1V9VVMUKqJU0uF+20iE8n6KylTnq0U
e4dBIVXJPUatqzgqGrQgvFEdolSRaY/Up/Ms7L8oIp8nQU6+KFvWy/V4gmwz/VLQBhwiJ+Urf6nZ
FWPJeQgcdZxlTA/iDrd3k5uQhNMMrA67CUuNcV+ZmCm0MtxwqCxubVjklbex8hKviW9JznU9KEL9
SNGf6mWStG2QwdZDB7SLAEK3eXScT80s5iLSbm8GsP2aWyE5vBUDQ0Kuv5T2mkcjSx+MagQWQ/de
lzOmIY593rlaGBxu+jeUgimeTcOdZZW0NYvOJq1vUk0z3sRkgkkNGWSpw9QWHl3oPKTtIrOjcn21
mwTpCicZK/S1Su8IOIIkbp1teWveC2VLZwGijH6Q6+9mrQg1w+Kytqoj0jIls4B9iqgFb+6wZmya
ozdATGkWqqr1p/9laDpqGUmr8Eu1KJHTprQqmzQ5dNOs26oYlpc1qavHM7mva4gKcizYM+JFAcWL
oP2lvFedGI4kbrnuAknG5DrAHjHqmK2CTXxDf7nl2jg6EKzcVYvGEHxvBOpWxgjmrU0yD114nTi+
SOCsRhEG4S538YSj8e1It9BKXKLVoh36xBlj7/+hsmNeit7feIQw1yiTOA2wti/XYgeWjTGvAYTR
/m16FtWWV84V3RInFXpkZ9qJ7ZrXoj+nROwFXSMO0wLkH0GwUjGAT9PGDQYBgZXuyXV2Sn5rXR5e
SyVOicWZHbXF/QSOowzgbc7vhFaJIg1pcWyANhzQW5VcjexEF0nkH1xcsyokfTPHX5v0sBX9N378
0qReAwyU7RJOAWtb5YH8hTOdt1nkkEnjpXUE/TFmrxe3ilWGzKfJp+/IY2akAmHUqWZ6WUbsM3vy
0v2ndjK/OLYYbLTN9lRCyfPtKRoUxYv8OkVv8YGFCB3VZDr9WHYmfKGE5vc104vpKs5vp3l6boLR
/zqouNtKAQBU2BMlxWeAXd2bJ9kMDzHFE1jsA/L/Dl0l4bWjwNR5K1B27Z3JLd/fVF6tQtMr2TFh
bfXXROHX11KAu4WObRqfmNJPix62uhUOo7n9EHBWRkUq/8PRw/Ztl/jI2h/vmXtKnqGr5Ac5flqP
G59PeyNb/IDn1df55b0UOTfQKiZJEmOxRfvCITkxwiindGgLnFaJ++7+2DIagBx8v5sJr0x27/kF
r4Lzi4v3FadK2J9PgFQYY7BS1poFfUaUl8tNW6ipamX6BJKj83mIc4C+3Izb2SsP7+Effr2Tb69L
NeXJZRrPeQJobepapvrYwrmfQBjSoiB380Z0Xt4KibDKI3ORi2W+37h+810gud9Sn30gE7cMLsc+
C5yT4DHyLlO4pHY2+YLzHFLCvL4QXmJkW3UNoWDjN7sQLugyp5SugP2QAJ8IZp3q6qTJeKmqE932
x77A4tIPIKyFKW8niP8emmMVGECjZ+Buw78JlVhDJuRxuC5ti4dp3g8gkGvBIXzFMkDBCLVpHS2E
gD79ltUj+6yFzAOdTanARDfYLUxbqKjJNZYsRrhsN0PLBEhZYVgOD/SZNIoDUKdPwLfaTxCl6f5p
ifWOZSzl/Y/r07qWMG2/iaeeDECNW6hVDMjf8Pg1HPqOOLcaA9bXCWymHh0jotcS/7oHLx3L+9wN
Q2JRlwR9XJNK3lsPjUXE5I42Z6NPUWnKoYt9GIFNAcyCACMg2/A6rvsRzNvjS+cIuBWneW8eVxiW
fUxHum3WLmhRwscQsSPW+RxbgfXpc233enKABOal/9WBiaenVMmD3lw5jHfJswFWj56JrTwVx7uS
E5/GmGTwz44Evs5z1AQ012dB8b587gCzgq/YGpE7+GI9FsiuB07aA2ToQBZHSBeeLB5feFGOHbQR
WWu8qXn9DfGJvFvJoXT/PLKTsCjOhf7eIgxhyCTtICKotUPSFOBqdzy4K/YqsFwTGwqjuhHZxKOj
40QqRQjSXaTcrmbzXoXOADlJ3yMJgyD+y77MdJeJUgrD9OfJdAflMP7rNyxp6kbcmE4vnKoBuaDf
eRhWzutGoZCgR0e4Qmn+AqtCYfqWR1cZ/XsZ1hTkq+u8J1AFON/8skjVKvHNtTT8ii7Ufe46ahh6
H8BwgAiTCLkmtADSUxI4l6U1tg/oC6CAIW66OtcKW+KG2ckP+TWbO19yIQvRu8sOrFC2Ul+CuuE+
ByYkeazShJGBlEDu+pE6D7jx6SqOrsc/k23nJ6GR2LkSEdegH+rpZ31VnqxfmmUUf6Wh6sBAGjcr
tSg7Qb7gPLMyM8InAtfbmG5jF8Ht8khrpg7JSYzXFaQYY2O7hLPBV+1ghgrIXVGMQkyRNWfjH/WL
wVh/yIxc9vndittTYxV8v5pM3EqqsczcavjOUZa5GHdrMZDesWtKwyZ/Yqn2fWNV4roq3aUHVcBC
oYSECdcZN2jYAYhP0L09qqZ2dQM1GpDy99rlKO5PdSWqKRRGwbVpjEtVNcg8sqTC2Z3DwsB6kD4t
uWYpwa8KtFDpWM2KfKdTUmpMDSCgC4DxiW2FSWhOnj7ODZdJ+YdEIATfwCimL9AgPVRp9MXmJsls
jXeriGJ/xsYv+cuGTEDz+W/F3j1GebDQxjQfCinrGJiR0fDAj0hHT0jVlX4P1CyOQMwoBDR1BIVh
7HqSvLcK3QiWbH+I0HQZHJT4dt6WxZwL1sfBoW+qi4rko1LMsQ87xw9qrAwxPGb0H2Y/AGXQyRRU
RKeT+OgZ7altzNcHFRqXobl78QExivQP3ra9kjMf8ZE38DXtjWMS+eXMfvu0OAW7WHnueQdfW0+E
HEiL/AZbDKQ5DYHmMnYifgUYX+VRwFhA1SDSBSL6qjUXCgP1B1Bc7oSTqLdw+tB4FBN2Gv8IA5uA
kv+Ab6adQojUCEtKVUM+yx06DiUv7C2iTNp1/v2wMV8rnRxa7hm5oey7DCwFAgT6wapWOW8TJBax
HeRO4Uokx1Cs0SKCK4Ai7LvLSAk1FDnEtnZ2H/+hcYLP2mjNRox0DRXFh7l0nwn1BGqW/SCn72T0
HMlA9IlRvWbyqdZPsAaDlmvxoHygnp0ZiTnjVOTSVSnQcpGk735wyHENwMycIxlPmoT4uet3DE4K
QXFcyctw8l/4T1M9GELUc8GLdDKeI2DqfDLc6cmXQbYRQSk2hYQB7LfOApTSiZdJ0if8qOuW5/Tl
WNU7OeLUfltch2J8AjwHULVKXe5McRiL21NxUjgZiWXI98ak1u+Rl7l2/WY2buKx8M27CYyD+Vbc
AidaGSg4x77baCIqWKqMi0tjfS8ZEhenlRGpzl9Zhph+wfF1NHCL9AZDXaGfzZydaljCDA6QS09l
fumni8YmpDT9E9hiUnzpqPH01Zc6Wk9WdlcuTdR4mYgsPW2GmXhAR3eT0tiRK8v+fAAUNhz+ciwa
KQBZmKl3t9AC43MBit9WIVzDz2ZZIlpzXWqcr/s7OP0Kf2xp3iGBvZmBPemKz94CNn/ZRvMo2ox9
zjcba+85PHeRKogsQBfUj/kx0rV9o7qUAQ0debnpDc/i7kPsrkLhEDiHbwZH5e+AjE1WryEKqSgP
92uYRV7p+krffK34rwx9G5wJE2jPJ2/4geV4Z9WCrrLUst0iWanuovGStk8g5djp/ZxD1ZoxQ2MY
MtFQjPvqXyReq3fuBX63S7txdPjUcgHr1K98u4riXHux8ki6Tzt4Gx1TKYn2Og7Dtn34mf0qA8G5
ap1uGXnWmXxPRD2yj/sLqjLCKJ03kJj+Qi3drNFEU5XLP0aVSdOHJwrJbg8pqL4iE+saG6ErpPzn
7AahVCt5bvoAE3DhHc4b+imJHBsb2Dl3M6tZ3RpUnUAKFQzNJ0vvXdJuh2BjQuc1P9QOvjkSi9AP
yac9XpSrD1ZJAwXpJ85CfeH/oHBsIcWnhNTN6pQZ0eFSf2j356eLDlWllNv1Tj/mlZ1WFuidf0aH
mpzSv9WZVRwYWYS5E5aDGP8imbGXzJbYFEL2vsoIvf1jhYqaEArPtO2ARCl2DYjNTaleBvUqTw0N
61H6R6Im/UPqz42PYGkIAt8tkMaGQBkitc6jnMDV6dLJiGS0TJJwwtsDnNgAjllvtaVBNUBW95H3
EF95AzJFGTTHdsgBAukENmPL/NMcfm0ZO8Jy+zgOqwEKzUeep9c9uxeSMPonG6uJIlU6QB15cr8Q
Df13Q+wd1NG0twj3mYN+FSjI7lGXDFBEgXCcydUnGynQuImE/kNviS7lQOC6jjznnupj6FjxCFSe
vJZ4h1s5XoLSn2ulNBpiA+o0yAHU/4g7uzkt+Uy6kkhVsdZZ9tfxOodqgml3PmrK6YSoJEPIRSfH
vSRleFhRRj74QW8H+IWcrTbXZWPqEuUp57Q6SjJ3RBrEBTLTAUzWq9nm8TaNBTK1nj4Atz+daHcF
5moaqOF1sVAOAAZg3YUFG56AhYdIX/8NFbl9KTaW5zOVSJUgMhlTt+zIfWYPdiVFRo7opQ7gCmEd
9hpAEH+dVN9rDakrq7MxuqkLyb5F0VhnAYSeW712viilIhIUrxcUIS8et7TODwOvKRU2aXEw5teA
dYYFnKR8E1q2Qhjzt64AE2xoRzyuVV24akPw+bq5CvJTzRtQ1NPDg6FqQaPoGRZ99YvozCmN2wt/
R9dIHBeRKMrJEbmf+7PAmF8oncDLcPzwXtE3BZ7C22DWPJp0NwdbzfLgt0jv/Z6M7KJx/t9WJlgq
SLl64PLAscHTf1OvibRuWMKRMNJVpDWSFTBSFj1gU9CGYc6B4iJkpMo4NMcuQmfsPmD03OSiZpFn
C8n5uUfaPpVVk9U1Nr2eYU91TNq11UKgtb827aUheXocgO6wq/FwoQmbB2kjkX/VxyYITR6UB7+S
XDjcdAFaaH/KP3skiS4tvtbn7aty883eF8W3M+kZTmWisGpebSxlQaJVsKnaYpOqEWflIGTPk5e0
8VQK5YNBltby7+uJo6wkNcXL5BtDoCfifexpNne4NdKz7zrv9i2xvLaLiK+kv2rLFBVXiqhyMaXK
j1DwOEkojXD+A3eMmevVvugrgNaj8DM3/gFmKFz6m70BjlY2jRrUIoZO3dikYsCNYQ3fh+8Y+sWA
tKVfNlpu7nA8OLbkqXWYKGXkDomS4EXUzBlSNWmyYIUUWBFW7gvlKEAjQwWp+bXTLy7FcxuGanOt
5n0FCRTu2fRjIxlakututNDk816V5dR9v1cKNq6fkKbalYXpZQn61HEEcck4QFnkeeOLagbzVzUC
uNC1bPSLSuk0ADDfr1+hHnLdBYBBMlcYPVgmSuLNx6/z3vrQSg/H06DYJEb5KveaqFvWkVmNYo60
hmWwRxsHHP7jJhqMw8aMe8b27PdawIfCneiGXRzN52C6oy7+dqolKZx913ofJz9rRP14BK3GGFQx
UsnNgypl7O/CZ5BfQXyXffiwxeAuEYMYOgou5gcEfLBgJGrQTrKcBRvXWcvi1vs1tCaFVO2JyrRp
m42ASYvAfP63oDSwj1FTcnc/njTFoTCCQ1e0AtAMzZNyMS67DVzBKWRXdqgFS6mbpl8kPO0jMW8L
gkmEw2TYD7+4JklxhUNtGIPa2a3B4G1GVDiMJFuYH72AD95neIEg2lfQdxDASemegwurJyGXpY2e
yBBlqfhsAabllPOO50iBmjl6hpP/sASuTHkqBaGVAtg9mEAJJT935v5YFkA35W/H/CNDmTe9QXM5
tsVB1aN5Gj62JrCJPF2TZIn2bDOSBFLBDNMJuETH/x20yjIa2XLskZ0qI/QOEoeKCcB3OVs7pAos
1QcZGAtKcTPZcLmrDVfNsYN4MENpkdCCCRQNCz2JrJ6wHsHpB14LBVeVJbxJLcNYtc+FJrZ1gEDo
k6M5WzXewNQziSFASQN5Yz0k1VPQyuyM7bWMNHETi/44t9Sn1pgUXUqrzglSUbQxsqnBNRpo+kxR
lNnAeyWnXdtYrza2jcqk9IHNrW+16JylEvzhFMjYlK7qY4ry8MXTfEF+S2uXug0aU5MHIxZu7z57
+LFs3Lmc/8TpHlFfErgIOhmbvZejy5Okqop+ltwHaBBJfH3MQD24Qo5C/XNaQYzjmJYlwcGR8A3f
GF281KIjk+BLCa3CmYY9GsEJ2iv+4xtK+9hAPHOjbz6D12L2CKCCIvpEgCj2VgoYGJWWHR66r2Ae
q5/0Zu3D4kKqwxBQ6LgaZxGLYzJXp5DWLcJtamLsecS9rGb8kXqQpAAymH07pMWOBXPBKy/qK579
5pWPCS7IycE2HZDyk0Tj8J0kmMUxpR5FWxtIxjuDin/RF7PnGCqTQLc/f/MK/lfBKIOm4Isn3x+U
RoiH0k4/WUrEZcn+I4T98c4vuBMpSrZynouFgx3WVN/GCM6XaSB5MmhyPWdsDUvRRLfrPihJ8k08
BUXrJcQOKtvp7AKE702YkZbguUkhU/EDgbCTHbRb0URQbl0pdDF4SbaDoSdMnhHIEYJYJkHoZ1Ya
h8w1EIer4BJjoGflhiLO3vKQ6Yhn1/TkSFSeoQraDUszZoFnVRjUBcV4GoYuP98lJF2Q33WXMbOj
vLLcnF3IZVHIid29EQC1SR5r1FbwOnGvMtRYF4+fOn+vL4BL64XavjB89JvY9NFxK8AqtoHgHz6d
LAonUdrtNbImpMUVSjVcDwH72aS/42AWcSNM2z0gaKNwbXmU3zkjo9O1JZVv42DLVIqU+cd9J1KP
xlupT9nCj3QKaLWRHNTYxSgVRsSpTna1PwnbkDM3D0cUwpBqC9R+XAdEvSBkyvdI7PV3yRs780Gu
UXCBIW3PDCrUlWQ759uGEkp086xjpq0AQQjc5l7NU8iwamooSeUih5WQ+B/1xyNe1nhUB4e4MJEV
Fx0AZ302cAGVsVqXQKjMnNKJ1NCCKmA6az88tkk2H2cjXBugL1cFPsdXir26aAVjgla/PjVpNtSf
2Q5kCDQDYGy8Q9vYjtWrywS/VX9rXDX3J4TuY8l3NabJfHn2adh9cpX7eNbcghMltbw3SiDzWWyI
aTIhCoTW6GxrD21wh/ahu7qkvpNC6yBVLMdUi2n1Eu5w6VgYlhaYYOnd7Q8SBdS+v9j4dbpyW+X3
GfPtlnsXtoIOJY8n20rLy8t2uuAkJZdoHOVokirtwLRs9AUk23Ypbmhdb+rZjf+ZtUjC/cxRd7k2
3cKdxPcT2YXO75jCH0OaJu9Yp4iFiY0fMWH0JGd4UmetCW0ukDuc/BA1PAa9zaiM1UAOCnMsEDNr
SP+Di9FXHQ0xtLcW0flWYtiKNopsxgHLtyIPYg7H5coJtFluL/PFIAIuK3qySrCW2kJoVCLeeb+Q
ORk2rFGT1tjUCvnrObVwAR6M70ETDqT+ij4uqILyVlpLmyi3t7OyPA/cOTnzR9iIs1hm8NcMKlEu
xI/GfSdOuDyV/30mw2jBWbFQbC75TdwhYacN6RKDBTNF/SAPTYNSvGmx/Y9RUKv36O3rBu28Tbo/
cQMwsbPTvAtO5JlLD6zJJRQlR12s1gYPMrhrPn3Ra9hn3WNWOD6H870Q4CBs58ypCU3zMI3Oun+Z
iGQCBpH9fDxtlz28p+M7TSqX2ff23KVnYe9KLvw+5c8ufRTtqmlFfCBLCdggW25WRL4/s7EMneR9
tWWTvSZ4F+axEGnTKjN+npK59/hcpHBdcnmxUiNYGkE8qJ6Gln2UbXRMV1xmjBgyh0xh1WOmxTJ4
UHmbLdmtZ8WwY4YY8cR2030DNhi9MoCg0F9sXb9vMN1oXL0go64kDopfU2gz91pDuIj9MaRWomtO
W6Yi97OxaaDBHCNQmSRZ22bMnsoLJEHY4+UpOEjZAkLhZ9giNfgVajOEm3Tae/llR5RNRXg/s5R5
qT7TMoait+ia/uemAmpS3Hv1Q2lakNNxkXQm+wVMLRlRb8hzr8cLNXMlx0jO3UjhBGL0V2MFXDYY
auOVJZRGinzlva1i2RQGknFuPgoFYUXhOSq33k5T1CGekjSn/hXU08gxUvxZB3yyogeDA5Ctrdyy
pYLEW3bdqbFzZHy+maG7652m/aRS4PmkdAXV3VHEpaxN2bay7PSta9QMb9uMsk6zVr3amxhVKA/t
59d3qKEOkNmROFCw7+RRWAwLEuQu8YoW/v0Df4/TlcDgLxqoqbWmLgOgxdIWwH/j7HWhjts8c6XS
3fsNdVbHqcUugQGhb7KqO2R3+W31KZap/2bDNJFd+BL3VncistFeNklrCljOEG7mnD57PCBs467C
ielR2ONR9BVb2wvIesFiubqkieRZLyn57wa9OWBc8Vq4beVgizYM9AXoQEfnaMxEoaJN0+l/ChrE
FqLXgNp3QzaBxT+Kn/ReWy6dwPsMWGyYoHsLPY2kGYhlZe5cJhOR85jg2W2H0vznAbx2XWnha3uR
Dj+QkP58MuG3nzL3n7ab8BEK9RaHfMrueFqPzRctnrZ94ENw2KBpiBu/dejl+ENYsOnFZj/2PE8g
ilr5KHJsuMLFOdWPwt0wtYMTrQWiOzO/6CTqht4by2Omvv4jDOLsuyfysxvkpEipfb89a/8TsVGt
nVUtow23nM/jEhiB/KtruLNWbL6EuTGwhgZ/xdPEpTy2SIvoqAxdjyYofhvWl4OALQ+NUX6MWslY
9t0ORgyQAl9lf5InCKjpGzfYecXyAzRF9P+FORCD6G9CpysvYqS0mAcDixfIblBXXa1hlkoKRpAQ
6e10rfcL/qj/R8L43dZ1d7NsjBBM1mdQR4FC9csEBigZQ1UYsJBAtyc/75UYtDaW/QvFBb4p7dn+
27YcRI0LmbrsyEJxIUbz5zPJ78eUxr04HTHspzn+Ho8LGpH/PyxJw6LmwCzEI42q7SEbkwsoPUmQ
z5csGXqzlzqU/45d+FqEJ24CFez9nGiH1ihUhQa9Ku4XcXOd9q/QVHeEUJpLFKYPw5LyxqzAhiJ5
A98T3KzVO1dPLk0vvsIte3bJSmIjhZFz3Dkuxqw4LttBboI4I9zn01iARSWxb91U+GEMTtaSPEhd
I2pFQ+gIn7PXUKNCEgbvj48VM81CXiQypX4bOX2jh7XT8wkpo2D3yeb2XJSbGE1B212BVndjV7eJ
RvABnDR0DuKyd41rM/nsL0WKD9DiDahjC1AiKWue+QjWCfKH/IPn1FYHIkWZLyfTtmJs6P2x/UFA
U5rmHGa2j1Xh7pnyYr0hxJ+AyZqYGc9x63GZs6VI2nGJtAH5htvEkUQK9Zu+XpB+GYDsCUEFgOF4
9jyrKmnhSKcgKWBy2m/EPuSCYyFwqjXCqRFS4KGF4jWxtmxJVGggdJjaMj062FAxDxUCG7rdyG1P
K6vX8ETcp4pyMHqmeW3C6kZhy4AFztmidy2Jq6yxlQWMddnLL3SStc3HqXBfV9n9QIwEZ4TEvZEe
DLXleoaMk3XXUtWIaRgIJKgM63wkte7ipMoJjyLFeEf1YAbwXhUYeSBBNOsLwnsaFjJWB4y/R3qR
0hcMtCs+lhbtzPT2041utiseGSRnyQly0ciTBkSITXgeC1AmUCTvMdf5nGkf+CRJd9/XnYUQ/NyD
iLSj7exMh0VC+3RQBQEeR97oB/+0JeX1QCjo+xu1aqEbEYHvP9X6OygdOjNc/wK+ha243qr2Y6W7
BrNvKsRpZzkgGYO+zKgQ/bB9qez+suJbMZS9IHuzS3CPNkp03NfZK8pDimtOTZUC/ChLNaTv8yoL
ShCWUwjlhuvFQQVMh7NKtwbVUWdbvrWpOLHIb7511zC69M4Gr/lE/mqRVr2kHLbWQYYO4qIfX8/h
EkDewmu5soaLKMefs9JnBx2Ztn073By9rjs2X3kVazQXjv+ccsdDMrB39qgYNZi425lYbLcn95oo
BeBcq9dSKr+g1Fy/8aPYZq3TkjFDD+PRnewH8jmd3CcPa7iJVaERj5Dh6if9oAYUbzTKE7LAdYxn
H2tjwTRF5KLZEwH3dW1SEp/EWfiRJfRfx0ulUJnEtgAxCq4mayl8Ve4BhM9YVLdYTA1AYz/oXffQ
7vAmQQBB/wZCSLaV8WkFLPDBgG/MoXEbjNVI5ZCjm9n9+ndGIwABeqn6JJABlXdmt1Iu5mtbVuqz
BkAqT/ed18i8gSQMNpFSCpeV70gj5K1gbYmPuCPHtblUziOHREcJ3keUkLhVrLHW96v2cOCe9Vdv
7SZuQAmoDkbLxsOHaNBnOOqNsb85ox3Qhr0ul/uRVkgsiT+s0HGgVsqh+gOfb1X1c2Pu5ufrxNWC
8wzeaNKogoYdTdycLKQhzQ75VZWRIt4O4C4wTZb9+jr+plWoUhlA3h7IbeCLmyG2Tcxa/v8fYM3j
2pk/uedr3tfrMiigknTJj1pb8cZrHGdLHX0rzEBYe2z8EDue0DwxMtNwgOeno5O7px4ADbtn8Dp2
ZsxnbRw2ob+ahuSI0wDCsiVOamL+DsIkyvz/g3PK5/+ajYEI6rI9a2u9rHi3w472UgpkmvPqa9qw
X/eZ+locWBNZ65GWPmEZ0r1KC5xKk3SN9C/W4Gp9ZWj0hDi+WTBRCZ7SjlI/LRd6NLTeXVRC6jR5
OK+ZPnIIQ/VXQEz2Q4GL+iTdi6FCD+8OxrkxoFWtCLvKFebBwK3WwIL7l5YmaWXEmJugbOuVLE2s
qY8GkhyY5pgn4eWq6ZmyzjXMsSGSOmW63Kw2LqL2SWsJlzaH2h3k3UKE0KRT7hLkEw77UIpi15dK
fRJYfDmLyO/DTHradS1YSDfWIcnQ6XNVMhxQKFFRTkE3mHbK1PIGacHScxSaXOXmYp3s/klgslh5
kcNSYEYeEZkvTs2eJ6ZbZfS8SEbyUP+Ygz7pU6td3vCGaaz8iX7SAXlTSdyYf4oUFb3C9p9Qemds
jEp4ATdVdNwuTKGD2dYOuq3+Txb82Jks00DuQyPD1AzTHNpYIzbreX8x9uz25uKn5rGMdfI6UwQ8
fIS0YoDfo7RoVzuXJOkeyojpRdWYHL2Y0n4P2biDyQyEw1aHDyQPX7i8hWRmyUWnbKAXod3UBVdN
2n0AtpvqblR1LsYy41EcOXqXN+DL47wmqp5N/mPqrVoVKVrL+K5Nw8H/DGagnoypJRFzeo5UgwZI
LtIEShuUsevm2IMJHS2C30g6E7oFK9XcbV8AmbpF5T7Yls+1afMcXnEoOqDBjwolT9PrzKEAnOOY
+vvWYcyG+AY+4hvq1Ytla7lAFkohx6xDr1eKGq7W/AbBfpszhA5re/MQ0Os51tcmrf99yGYSP48j
b8wr7v3Jam76AjQWSG+Yfx5JsJpqezGsDxq5LNJEBUDXd2dhHLAYRznpn2pkd4+VT+luEb+fgJpd
Q9YoEL+kaW0+NTECo4PP6ftVzYa4Jt2aY/DnL6IG3B7ly9VWVsWHe+GYx6G1bESbZAUQxaWmZv15
8vSNsPwbOyN7wYHCKj8N49HElgzN3jviG7iGC/o+MhXbc0pO3ezckvN1RvKWI62DJVBz2q3zW8z6
NUZVszJ4h3vDA9ImUMmM0amIbH2DNwZea8/8J+QXltOgEloTpXVgSNXO8a+abMoGJXb3TSPqXkcs
GlTjQzbKCgLJHgzl6bMR/Jc/rnyxwSlQP6iWh9HU5S4SnvQlIBKHaPOFg6cAKlmllJBNrhJjgvlq
tk0L5Xm6Stvyhc9P40uf/C/vFkNJbmEwG/O/hJCh/SU51Omf3evOS0baYUhEBnkQmFmmyYI54+w+
M89s7m00Nj7FBEAZFVXIYFdopJYiok3bxnVd+JmUgwVcb4A9FwpRjlR7JVtEM3N7zUpL6jzu3+fR
kimtoDBforO5nz67wtk1ySVIdL/fkL+rLvo5Owj3bzYgp04pdxqJF//ZU1yWlmcQDKqRwLO484qS
bHURTiFnnXUZebufcSHBXercqSVkNm53MBO2vsibCsOC4PGF5vYwVH5TQ7dtC++QZcj+YFeUk2r0
pqLw28R2DaG9SpnuEUS5HQ+9/8T7c2PSgzHPrrQ9Z6BBVskb9M+0Ltr9kKnhwPEmjRxCczZ7ux50
rzDV6ECJ7zGsxFSI/xtOi1EYbEytra25MaoB+hWVRgyk3QdsGlxhyXAMbaLlDT8UCGhyVpj0WAFT
gQtOH4TUoV4t/jRpTlUuOyuZtZFL3kV3nHJTPjNedyTVczH8iEkFPWYHQoucB5z7r+z8kpklTOpK
t7hmJbwA7HUZXjlbKpRUiLytsfoNxhZJJ3Fl8vktVTjp2DukmO0e4zWkewSjE24Kjfi9gUYNw2DH
ExxfoTCvTZuPuVzeMCAbSWuf/iTzJjzpuR4+L8tsoJZZTBoOrf180yGvmefuzpbj/DB3A4EPlnx7
98dRJBSN8zFUTAKxK/xiJQHTofkq9UaBeDm+G8FylnT8v/7Ct4oXKc2dBIdsN0l850vkfQpD84k1
z/QKFr1sGPrCpWzzOmONB5AiNFi1of4VsH7pz4yiQu+rvAgAKzcINp1F0ovVwsb1tVJtEzCoZj9M
F2gMykGeaZ14Nm20afCl7Izsfv7GhshbgOWGnjc93vNCLx7tZGeF4R8j1QD8wi6RdCCWrfDqGPe5
0KHWw3+2UNxERuwKIWlkJZFZasTKIesBvEnF2g0LkaOP9JmcynpD6ARS/vDZYL/P0pvDQw1HhSC2
25Sjkzb9gcHiopMMW/bQblt16LzwqEDVc6o+3Ek0Iy2XeSfpRUh23NM+JaSvisZ3sCLcW9tQanht
i1Zx0d9N8RtI+i/tsgzzvh1ZK1QCGpoUkW6IZs3v7B5nZI8Cim3gC3udP+TPFKAusrohfAb9GQ3l
i4zkJQbLIcIA1s9kmAE85kLDAkqfIKO8pETVW4AnPb3hTGdGbWg84QHyzZfig+TVZ1aa5Se5Sutq
gmfH08xJlUL1YEy3E9KCSWaGe8pRUCiqlvx2n4fgF5cLRBFxajKrVdAig/0dTqPWBi/mYnHiVp3J
SH16AVjfjq5kdKmo8lqk3xnL7lWOcNVBz8MXw4tJ2FHdNrBD2x2rSYGjCj1Lk9abSYtNsXUL/AXr
Fw5mS+iq3zyYU2SI5Gw+4478QdJ0VIAuuCAErs9aHbXR+gb6nqld5/0xDFuokW0mhIqer03CoGS2
X2OcKliPQ5UMskThaoqd0ioCxP0/DKHqkxlFvP/GVKRuofND3QLu+XnwCNaDRgvFVVI/UrfXHygf
bB9kED5eIDCHmw5r8OUFn15i3ZZIEZsRDhstCQkwC04NxzRQzVvmGQ1dDbw6hdofdF9OHUq5gdyg
im80T4UHqpbP3ufLQQGmU9KbPqVkwXdWYccBdxXMf5hDt7EymWiDNUMugtX+YgSWRPLnsDIAKriX
vAcpr8aBLEbm3ncJwHUZ/mc/zMZHe7yVgxvx4IuILko4L/MGIF3V0X9R2L3ygtcFgjxtdjlHcZEK
ZHXqLf/ZhJ4FLdu26S380NmLxgdu04m5dM0mCHI6LjlTWSRBKBOnpYqECIeOWEojCO744W0QImMB
h3HmvbzNnTn77wEkbm/pIOTWzEepiibRo9MMGSEAIDWYyizEV2PhryA0d5kvFB1kjHrMnvyznPkj
gQ+G16VJyAXGK89QDIIrfnwxq2GdDxqPFltDVkmKJnvAQ2G/ehLKXgaNZ6/JIds9YcFPrbPgN7xX
xEZ388BUOXoV8q7fCfkNreAmSDneupiE+yel1nWdQDnrHhcZs7bg5GEKv4S+WhnLMma6yQQwxfXD
7NYlKUQhyqoWsxY6ebWvHqffJ46cPtj4QTN32JkdRP5O7lcCokT62PSApu7nxD3iwxcSnAop/jyC
ox9WgUU0Hz0HRzerfCv5Wu/C6QHf0Dy1oM3dR/R+a/MqdhUkFqDbt+RZtaZUZW2jdH3y6XQNTvm8
h9DP1b8gJag7Nq9YpNQqIpoLDLT9eHFmS3gxofJY8W0dd428XtKWsnmIivnm2bqWWTtFTalMYfGg
/kKKUqswB3dqusw0dW4m4IxSLTnljaz9x7kCyMvIVVEyb7QTamdfk1tRaiLwsAYrS6jJkYh0tPrh
1qRLHNCkwTAsawLDVu9YsgLwL4BJrjCjaC434HXt0grEe9F9dikbdVvNyBIN3AcB1ZfVAbdls6AS
fTJVu3ahNSCaqEaayObaiA63kjjibKCwwFruL7BnxH3Wx9csaoXjiIs91GcJMk+lSTTbz8nNdeG8
N08Uh0fawEwCzKkMgbYiPW6xHCSSgsV7PV4/e/qc8oXcp7nTxMXoRVunkaioEoSvT/EJAnnlWCVM
OCE4lxdfXE13jGU4uGk1Gias66ZgpIrCOxJGMvI4haktg84TzFUlqDuwhbBNv4Ww1pM3cv5lvOJW
B9ToUsbXUDQyiObN9vQN8HJVU5wwfqkYHO63BIqZpQ5g990nyyMMZ26dO5gTrn/41/LRFXahVZ7Y
+gk12wf61kzMLadhNIvgZG7nywAO9dfE2NqNTPyUeDM6TvG0mrjDgiQ3aUwk1GwVl2QZvSMWdbTz
oPDr+QcLvGFBt3V6Pf9jruM6gwnNG4qGo2kdoen1LcPPjPgH+q/27UyHZFbViG3suKH2j7kitonm
VCh5uaxhNKv238haKqTeiS4CvQtNKDxzMETtJqvt3AuoqYvclSXS0p+/2oNOHqekFwnf2kcUebuQ
Nt83qItelhhtSMWTrawG+j/Q8jGS9fZK9WH2NONVEJAItYyCPsTSLJhr7Jqakfdzh4XJTiWSc5p+
wTThkqj5gSPcrN/InQE4U7ma3sbIW2JDmWnPv4ztc8/3oH/RZMX2MW1qRiEVS/kDBDiC1HL9RI5Z
FmfvZhmWfI0sZc0odKnDWfskFGNSE63pkM4mP+qJp/RTZ7unD56QWw0KTQ3FbE1AJJ7v/zqaqv2z
/YK7JMz2lFCK+4K+Q1LQYkfTSBG5kIFPyDPVV5M8BVmfIyRfFsjGofFlFEvTJky4m/7ZtnuPgiUR
3dMQMNx2oqzKquJ+ZUHL1s0u28URJT2dOxqM3FyWAyyuGV7o6M4PXIZWyQ8OSZ6xRgGovqfvLyuO
ZIdiQO7ZrsnGJaBrxDjCjX1/6NZbxWASVWdWMowz1jkEK9ttsyRb9RhkUPwAwWf9gufuogxvz38W
5CYQwT0P86KDT5D8bgQSVuKaTlvlvp/5r+71rli51oq+DQyx0R0VDRNU5aMo702xfRxiZ01QhpQg
lQkhV/aBx3IJ7sGjsfX0B8FuiXvpbBtsqThZCVAvlZJL//RYjVn8Ha1TEbM4DHwFi5CummOh3/C0
hEjOA89/CxfLcYZnULy9RxCVmIvTxroTgmgx0RDV9lvunDnkY0BU2cNbqzvKoZwKyrDOGaexsjtj
YmucCvRZDmWKu9vZ2V9lceYd4cMbP3vTeSWrZZ/gc3is5tXL+FtpnY1UH25iJevzI0pKEF8qXqme
4Vl3I6ygJrpVK/BWM/hTuJypvj6La3QOFxtoe8CQM0VPH3gWs5vnSUzhpKvzz72ZIArGhyXNoZTY
7CQDoV4k1p6QXLALl/7qm+P4ZB95yY8ywont5y2Fi5hrCZ28dhNodHIdZIUNRrlmcfM+gGlja0VD
5qGOWbKZuScPdImhx/66wGYRkuNycmCM8s+jPklZpkTjKXRkgFl0maU6aNquLisxZMMoFRcWNIgk
D6vahyTFD0es6xcCNwhCKaGhISaZLeAyxqiztAjJCHV3ulDNYMEu3JYSBBCJCqrzjAVZJt+2B53O
wwZ2BIbI20bS6CQuYo14gBow6xUffYznqOw8SXIybWAcxrjSktj0fUYMn3IMa0P6vJC0ASw/513F
DR49JA0z3H1cjUy+bcp1ofz2zm3ON5wdArxnNtDyrDVCSKmA7xejEypGIYIOpA4YXVLzy14QjyBw
DLNo+TclriIF1kSebi9M9garlFNCYuaUnIibdMw+sIXOQMQefU8ca7hmguO7Qw0KtHwY+c0LaIdb
xzly3JzQafZ5q2kGmOhS5Vzh2e6961Jq/l7wH3zKJZHQJzB/BaL01dG5Du2mxfVhzwQzkwA6AN3H
iIwY9B5miT6gYPoAn+O7DZCBjXD68RYbbdC9V+N86I1amIA8MAIRjS2e8ZD+RnIktDjph2HRnyZt
kJ4zGuG0aWbnQLdpQiEiZp0hgLBTbJbKAsgrCAuEauEDSLyfEjtisrwkDI5Q8JV5w7eQzn2PSkn1
1EZGwAhEaKVPwowN2iZ6tY+FgZX9wUEJkQRga/twnROYUHae6ya5UOcRGQJkrxAD64tsbHxn/Rmq
ZyYqKmSNfZkII1Nrs2yepyyasgO1bQ5Nr38zlic8XhyV8udVyHb1D6vRJ7BMY/pZ5u4zCX2/JrXS
Jc0APQH6O62tsMo9GinB82tn/lTmfytSV7cn139tab3GXlg1+FK748GrYb9WfGIQEZ3RS1lWbUxV
zFxWcG7/ty/xFkqdhG+xbdHq+nrMUzz9w8GrfroXZNxpIA9bz3p9o4EqvhQwR7Q06C172lZuOgLf
zDYYbvNxw/eHxWyIBa9GAE1f8gM/sJf4AcakHa8m/OfP3ami6aWeqsTOGb/tNFE7NWrdFbRyEbT5
sn5/XZBFsr4tDSFMie9ZRpZAkYTf6rsGtzYtX3Yk1n7l+Dm96GkwLZ7rIcg9Coq1Zh3aTawnHrTu
CG0SMtUkzmpoGZHhzeARSqVFNyRwtZARuNRqI5v49l70+HY/5Qhu/+EfKBXmY5ZRUqEL/Wp6EwKw
ynnacWH5Sk9ZLFArigJJmD1yiz0s603jltWj7e8pLLHjrJsMDd+jCuTlVsWblG6glEAFSFvytdzw
Lz7drN4QEgEP4Kv1Kg7MkUsgwGZtltbfZq77217EqeJOr3KctGSRySkN65h39eUeXfdTS1zJ5K/a
Mdv1asZGsl7iZM+BNM2lBueK8nQUdVevH2mFJXegdMVlMRb6nWCcnhCxUF17C+SQCaVp715Jsi5F
8Eg0S9Wr0sAUYEpYpC+Te0DLylAMD+Ow4iRK+GVBPPBDYOVcXD1q2pMXanAqZ4zE6u5JXMnTI3ym
jdhhUaL6WFpQyfntTvhxMN7DX4rxlDYZqLfZnECp5RQd90YZjPsPwVCxPP+IYXBsJFNaBtTzowWW
FMJczfqwhjitbZQgMDi8wvKtBfChgeB+FyLvmqrPOESjp8wai+3+c7DOduPDepYCsVRKBW+fnCEc
hLQ6En07++dN+qJOYxnatiNE/WlICO1iZscQeUA5Y5lG1Iuk+iAQmR4Pkt55QhJF8CmoikAVSDvy
xVMBiBx29MupFYqyV2EX2kd/M40BTKpAI4Kezfob/TxQNcmedwE/Bdr8su9VBubNsIjnxgXuqQTL
ZGkU+I7xollPUPEDdR6bUN/xCzP6l1JWo3vPvUnAsbH+gHlnNgp6E28sp8JLYmap9r+tvx1Xi/+M
NPpQEzsqLGUDkREkLgCy0xFdKZs+u/nM1BHQe9wh1rgPLZPHgBcYw4rTVMIrNexhl83UDZt7JVqH
r3JLxm5eR/LRPtGAXZuXUocVCNi3+PtykjrrjkTstum6yGDXLaHgGQxO5N3/YuPNcfC/jOLXNQJd
D5uc+qvMtJMs5i+HtLcEjya3jyecECw7iIMHBvWUYss4vMz7kL1kSl7ustIXwMsxpptccHdtpMKl
C1Uo16ag7EbBw8Z38TN9Uz9w21hdUbHIP4ZXQKrf0Yg75Sd82+8V6XcFUU4xfN9w/VSaZxn+JAFN
A11KaK8rSggwXzTkC2q6DjJ9xOTntpZqi3wEQ6HxYvqtR3YchIEaR5V2mmnkZ3CKaeeTFteMPwN9
MP5pcU9f+qRwDfVeH/duWDmnZW+Wa+6YLQvWsNL7R96HYM7F5y67ZbypdVg/riQf8+hGGAPjTN0A
J7mxXliwk2SWndj9rSlBJO80v9eNaYvvyW0hir23mNUXNKT7CsOblzoIMU3JY54+j0KRQpYYafTR
CByJ0NwwO6OKHX+KKvlnVrYpYl64UXKb0NOZ8BBcwXvl/hJl3hS9PWyeN1Guy3nqYzCPi6sGVUF8
znj+7+tSDEBsdfDDD6h5/RLl5Gro6xa2m1kLx/ukDh7dOkQapGse9z3HrJdjikLJBcEKs4WFFfcJ
35Z9CI7ate+KmJRDZW8maU1/wDC+r/QiRvpiV3z0m0+FwwsKySadXkgHHVUYUaEX9Sqa0mt+c5Qg
FB7APIc+OQZ6LaSNkK4OnMeBEaxHgCrHFpPSqRtbL8cYe4sWk9Q+mpElxcBU7KLGNhYj1w/T8R+3
P+kj43Xm8nH/KEfm3kWwZyKzGsEKbDutfRCbJ53nHOtnlby2+GB45mKA8hXmMz48NeSSoCjycm9W
JC/X3L0ltFBlSWzrONP0KjWdk/IjT9bX/cMM5Xig3hTSQxaTi7icEXM5qKemmXqy3L3GVpEn0yJ4
DcvLNfAalWnILeTsh0OC7A4em3WOc1yED85Mxpjq+EpEvDm/CHqRuZGzDuLHFHETe0K+48Xbh8vr
UPybzwIG9Za6I9CuxpyaItmK0MkxU2CMB8JmKSMf5JNc6YM4Xdv6+GO5+TvFI4q+SGBJY8TX4Mzt
+aQXQ/BskpqnZndMzODlPhufEaASChtv6zIsXYaHIkPhjUaYsLSdmfGi2+c3Tq76M7sGKKiyV7i0
orIRWpB9H2ZscC4KH18yQ87u2h0qBYV30vB5aVLxPOfJjVfl6aVWvdTb8yxC9RSAh9D/FLXcYerf
rgIEJiDXqkurBFLnLYJfCFN6OVAMf/bu263pbIr+E/pAEfzuw6zRTPsEFzkbeOMGdPl/v331Fj7W
Mzr1EXZASaFAk0AgKteo7XZqaavAD0Vn0VCUWbWX4BXQt1vKbX4PeyzvRUA88XHnzQiFvm1ZMGt8
41LXiXjAHXacc2DfzVq5R+W4NoSEPFNWRTyINneP4OmA1av/NnzYZhcjKkdVRbBuqZf9LWgtUd4T
UD0MOdrClbWqdl4XKTTqlhAEuOkCh1VfOZj2Rh8O1MF3usJGACOwNk/a/IUHcg76cloxY31IDnwY
PvpfdR6T9wid0Rhfq8zAAGu576WyG/ctUE/LX6AZS+zFiDv1A+bbOZrmZApcjhOg1o3MhzQvbaaT
d4MvC09owVXPtVHpzigdOrJMCcabGAUWe/vG1k6GfwDz0TPccm1dZahwGwGtzrw93y9CcD6oOYlg
y0QJq4C2rUP6IvCbqtNFOmKY5qaZdNVkifNembS6izizQCwRdLfVQ2jdfPiSR7+mzKo5c8n9niCJ
aMxivI9buNhZfdB+Fylfe+aA2O6onEqrdnlaZBmm0SzRXxk21CMbFxSrAtoJpkYjPcJfs/QSOx1W
8D8WRN9D3+9v0IsjQWx4qKfsJMgo+WEH8Ii88SvAeWgYP1Ab3Tgqz37NFZMzUF9pAFr9lv2nMX16
tvVWzFkmXA/jXoH4xLVbqp9FjlqnKyPVQ4WycaJSvXP60TgScrrzbX+JA8mtZQsy2ss8t3PWz2k7
BdkP0w56N6TijfDNYkAtNgTOxef5OcfUMeC51aLvPm7xCRGATzvJ9tXueoAIuM1KF4sG2ulPCS6+
nzIUBw9AlfZvad/BfXr6aX73nLNOKf0KhO86RvPDnmlN4rvTmcZaUitMi3N7RUH3Z+nAE1uWKNOS
Z1FgMZt33GaG0q1CgKFoHO0FkgLMGOlzYZPY1+UpWKzmyDhJBWYhJ6w24Az3cXG7OVI9dgfYjrpm
71gJIIyFTkLN4UfIxuDT3DvpW7xq0N+qqz208XXDl329dlIykzKQRfhSv29k9+pP0nOlHyehik3R
UQzz6R3T/X1usjfIIYrIU6aLxI61TzOvQMoaL6A/4UCvFtVd7HgyaZUj9XWDYBlb8vqGmlni33iZ
0P2uV4ZXu0bE3b2bnRi2ryq8u0waxfBMbtmiR5Ca+9SfZgUixA2Lsp/8XNk8IkCm/XnGNQ5ctiZx
DExNqZ46oGRk7s5W5j6Uz0SGTl+yCZ/mibulOFjYTZfbaNMHb1GkSGUp5S73JMrv9v6vqsK/nlpQ
PJ/VCYO70XDelz2LV6IxOTwzD2ETbF0dIuaVo95/BkEethY4qqLWKPjt/aeJEEIVeti8AziN5Sn8
0okqNPQCsN3lPFUgBgBNVCgZcISyAn6+V83j9rVmyuMmuCZUVne914V5Plr+w9qZBBOuwIHrcK/c
EqtQXBTEyPLal1Lycks6icVRpPBH1VEa+e7CYaAhF4CJERkQy55PgCsG4vPACQek9NNfbz84Y+Ez
QhLL4aV+myoY12P2vgP7KM21yfUOW4TgJX0xukyYdjD/9kaNCiaEHsLVR3gcNYY3W6QHSWRr6ZYb
zYi2lxFfwhhFLEqUzmWr+HNSsJDni7/P0lgkO15JPTdGRlEd10dKkdWCZO7tEP2s4RPiZSaVDLqT
uDfeAca9BhzYU4YraFUtu0qoO3lFJ8zkhaegP/GEpN8Eh0d8L+1RPdP39OmqfBGdVDSpvITNrpUX
R6KAszNk51MM9MqQXxRlvOuksH48m3kSCRBrtWLSqVQrbmhjLhoIrmDNRdCXK1dyQdHqwzU5EVT4
QaUQDFoVfo7lDs8AlQI2aYAqi7srPtfhW7uKQ9vIenXTCbnriV5dX4PB0qEc97pI5OFlywihmpm6
+lFPTcKVX33YFzKzvk3cOZ1j3SMlc5Z/yEAbHw02ubddf8xnU1cAblKcdm52vTU1drHHdi3BOSlf
OdG11k2u2Zj+zFUrwcOdTuBnAX//KkTget+wblOM0FaEvzXaorMT+RuOnkDN4c3v1QeZR6BQgF0U
f1PFiaVe5m0UXomdJ9ZgUqCCUQMXB/5mzzR5UplTikP4fw6rHXdP9tzbimATCfyfb/KdMeg/01wX
0lK8IKeAmZmhHpEjHOOL6lHJJow87KcCL3qAbBqqinqw2H0zRYKO4k+70uos37hmGREm2mg2F5YO
nfzJRPXS/dnYR4R3uE8qebb+FOI+n13s3LixI0VVkdqq8Umc8EGaA+488P/qwE+Gpv5uvvo56ZD/
XSH97OEbMkYBxmrGJ+I4Hp63rT5HIPn9Y6MM+9S1w77TJ/yQrDvhYLM7TEE7Xk2P39ItmVtJrjIj
XKFuolbKn2pEz8KUOPMOfCoDpp12FjiUG64Tr1pwr3aDcMvvmb16PFZrd4nIlARs2mjzWTs5Lhv5
H4Rmr2JQAHpAJPeihLdo5DKXIcvSH6C+iJEgJ6BPbtI7ZySjKzWpSRC6C1c+8iWlnzZjFvys/v/g
cf3TY3NypgNFjtfAQ/7l/bsZQHNkg5zqzlIwTHr+G16Bv31CmXZyjpcXDmln58zMWzq/y+R0JaJA
rInmB3UidIj12jr2E0Ty4Fep2Qo4o7mm+433JiKNvkfZB7bBUqojctULmkPmHA1K4JxYJ7JlYe4r
mo7qJ6TzvOxwYzDhIBvuivGDxr6GdWw2+kFS+Oi4q8DQxLjOeCdZrXTGlW14/3cDvWZAVk0zv6wt
SEc5RJZ5wgARZerOs3Gyi7pW6178dpCUkBgZJDKFV6TJXEbqsi29rK/hbkP173JAyRZOizgDEfcR
mkdZq+ux0oQn52WktnB1POYTmj/55MlmWN5dvMnHviNsMnRAeiLrMrvXw4nOZ+3W28Zz3mfyo8gC
stoDo6m+CyS246LFJ+JrsdR+yVBWhhVl2O2slpvpc3qEMr2u4G9832GTiWnDiWs3w3Ox8f8+qqp+
FS7hAgoK5eWCL7vniFNwNj1xon77esLEbOsqlt91fmtn1hiRocOuvnhbi9fUv008IGaJz2c9EMs6
WhUq1wkTTZQmEhWw4wJb782I+5YcflkUo7iIOnf/ro4mcMPeDKn97jguk5uP5Mlww8ENy4W8Q1zu
XyPUIt6oGZ52ILPTN7szz5kxCB1fJMZGaVJFP8kNj3jrJST0X+L/lq6GuP0RVb68WA+4e1mcRQPb
293knarxU4lU9FrIZnEhcAuUlhMq9AEG48TPXHBXraIEl8p2BNRWB0iO3JdrssZbzm2j6KcSd/YX
ZohBaQpXwX2RrYjIFp6IwFiwJVtlPNpUW+Cq3ZGW2CkH4ZSh0KhgDck1UBP3WCj4vS+P6S13Z84v
Jiex6yLmx4p9mgn6J1qZ5qXrIHMi483j5rI8is6lu71Fl+rn9pdqAIjiafivfpNGLlNnd+Bl23wM
HnEZzaJhI3upuyHc7PvtreawXvXqhxLcSRGi+gk+5QmAzkN3Us/JXsG97r4fD4EvvzZyQUGOxbyj
f2HVvsDEOPf+rCKGW/1OrQd1xU280gXEX56Fm0zTunM9bPjGAhLUfl67z6wqa3+c/nLu1ZTdhbA3
1RDClUnJzU5babhrjW0hiRTY+jRP/8PFTvgsCgvF4OHi27Tpt/vyd97JgM21c88t248OsTLpSclc
rij+DCPSh+BNEQwjAlrcKxxKXh1cFJpsk3P4FzNB/Wz5MxlL1VqqhUkDZxEdzL080Li5l2Ujya94
CA2WdHjWevymeRr1HPAJLOr3U51ScUDz0Nw8Tj50NhkJg1bkAiT0pDGtZe9BOr1mhYQXNXl7dbmT
trSRCwR/+z6cQ0HiEtRJZsgCQPZBQt3P6TYhXexj6edCLj25mmR2+c8MhlAneAFG9DKWnJoqUOK5
oytZusGjLxjnteZVTld9QHYVDnQrwqFUXuB2lRG37ou1cj7IawsbXnnutxIv/5X1nEHy0+jxzqod
iaFmksw7/cpc5BQYwUiTm6FkQrDsSEoDmx6omT1PV2fkdHzzLnLeDw1KS9V+TzePzAwesuiR8v2m
ctm8GLhLqN5oYWixPIMEm1Bd5WptEQoDNFYhwD16rSdJg4mZ12QbImHxaLfyXwLzAXok/Iq6HodQ
6io0flQqkoIyFtXRdidmJ/lQW1UWwhjFUMFo9XyJp84qbryAv0RFo8E6uN5f6PSsWzbg8bSg1qzz
V18OQyroo5EQdMFEmxIrVrbUj088kIzqJ2dKK5Mvt+RtkTNw91YZb/GvHI45XB8yPULTuj3Rt+lH
155tyzCHHVAwwlW1k3z2UcTlRGuhOInmXMllINxNq74noPQ4NcSdX5k7S9iH1vZUeK8CAvZ7fxCS
1btbZdE9kvhMnYI/Pq7QoYBRprmKxBCc7T0kpLwdZsUJNj3/uxJEyddt2TJu7QLsekQRiw8Zw5CN
M3LExJ4UHl6BaOUC2YZDiTUBxB23je8UG+Sg1EaIlIU2eQVjtclTLx1Ad2KHuJdoIHXApBJNxKS9
13tBjkSq7DYoXLVavX2ZFXSptmKBwnFl94wERatZQMwYfjfxi9HWnJiWk4XfK3ystKqccBZVivjx
+WR6EzHYHd5lMCxSOUVuXjNVE1r8fagQtakE4trNm6rWOnT7imHryT/G9i/mZi92FzxVe9nDwtTA
0Bw+9kKQJLYJunveh6rS1ui2v9ZBc3EQSPzUJrsLxykzjeuGquDwQsES4+KG49gG6PsjFF5jIpJm
gSpt1HtmEuJ9lAhQgHpVGJJNCLccUTLwUrpPOWDugo46LbOzmLgWZPP5PAArRYIO7+66mAkwXrt/
kP+aVqcEAXLPPxTT8UGdbn1xOZStd3MwrND9bSwMb/izDX6Sc0f1sZncv5ABpSr2eO7QYFeTP/Xa
L7zigRVqQQk+i/8Lc+KKr4mAYy5hY0Er2eyoOKQ/msmrIDyCh8g9eKEM9UqCKmEFpgqsJmVLMFm8
h6OlTrnCuQDSLe0rtgMIfaKXMMqnsJFgo384/69SdYqq0WOdA7R2Y4D+sDoOOYTfXpH94jLMy5BT
phvWMPMb0FX5RoyR/0VChdSitS5A1471uEeEvwVsqz5q5NIn0ge2v+cUTiXJQCwTZ5AeW4nyrl65
+Q+EyEz57AaNLc42RgB0nPqwd+nEbn1bUnXVvVCVqZGjAIm6jRM2mAJNzuh4EZZONOKnDeE4ot7N
ysSCJTyJoyoLavg4NIIhkIb3Cob/huTCaHwFV9BifUfA669o/NV5meClHEwD7aI4c6MC1ZJYWfrD
yyWeDocTZyO7jgmhEJcbZkBUrwt4T8srvHjz4tE1L1by3Vjq8+qkAdpUaZM09TWuQAFDzvLU9mrx
9KAn/5DRu8TGmEiM5v1my8MTWuqL6B5/VeAdQNf5P7UQToTLJ2KyJTVNRzuUI59ZtQD1na1/wshQ
cpc25DdEoftL/UM9l+/DLpg/S0ivR8870K9bgjHsDcu70+P7FDc8X7GFBp4ZA3HAmg6in2ywLdKx
G28W39iPX9vXpFbyUfc9J7C85h6abSCEa4VqeoMfvzNN0PrKOpPwb70VSPq9uC284ki3AwL74Idl
8XciXmtvU8Bbshk40MlSiMLjclpy9y4gJIlSYNeXqoOHpFqZKjpIXYiUy78zsxGXr2uNBqsEuZB6
UgbSBYaUSjUJvaTij38+C2nvNtUYEIOzbXhIliMRw46E8PUuObRAyiSvHw5tGDzcQdJL6XVYXZCR
N2ChEpuDeQhKYLJOQd6c1OlkPP3EVeggSdVex1Hq6VJH6lO5Jtvwn6A5cXaUIjNXlawufW93SbLK
VS0GK8Was9jRh6gadi8howQ+FrIhbooW/h5Cfc2VVQ4wF4NtnpR/EDHtN4l7aYTkeMu1zmw7bTb7
RS/0s0KziKasywovyda/7+M8EBOqx3MuwYW8pMPiVooZyIN04pbR2JuZ8+g9PRoTKYYDHfNak+xG
KDSITWYGNk0en2FuV6GL4JP+2ZUBUlWAN4ZdQV8VwDqPTZTqx47NvweBEgDOGu7FvEBaLw7kqrRl
OCaraZay8uNpyAidf1W/DqpUph4TqXV2ourcm5cGAh3cDUwLAXKlpcyQ2yHyKmV+x2oS1p6aaHJq
SCax9odRBLZsnEPC86cOyP9WgLJHjaMt/NZXf49eN3AMZwvQaBmqIJPpGBq4Ey6kezY75veAOVtg
aA07yDYvX71lE6WTuIHA3ioS42cgcevgjzGCsL7Qe9UXTTNHlHebB8pDP5S6p2+KK3W9yJ7t6rfb
PfpW2zPg5SvKu5Aa0bWgwDWeOvhU9O9+ZXckEHZxPWPD5iKOO1Ie2GNhI82/pmDLGXAG7rK1He3l
W7gZGlLbgsXGMrGUzbFE2HwORDiueyVoOatzqg7fJdMTAEtj4lyknrKPjDch07nHboSqM3GQx/KG
bYj+8q9VfOM0JNZ9QnsxfwlXEg4py6tIEzHjGgyHdLSXgvXJLa+zJ+qPEbpypdMTK1m5Ajnszsk1
LIjNXSpH9R9ZRt6KOULw3nIUd+nHCsm4LwQqYr9ssyZ+7V0TGaP1UCnT2Qwk28Xjhymfxv5uS1fG
wTTpDU1VKKDIVP9g4IGHHfQicgeuy/bwQvKl7IFN+scLWhxymiqBoh4grhpU6LZToT3QYxVE8N2o
ntoAxb9kebtfQGqighb6b7KUrf7M3IzNy5+3U0JctoXI1HO7VIXzqqZ4w/7SfLiiki590ojggOGy
TTjwhxgAulZHzz5UaTxAefqLCtW6NiqzlNWGH7SXp5587udVdVap99n7Cp7woF8trSEihHbnsmMz
+oVgzQcWkaDp/BR4mgiSjiNmC3kWXhOFm47Ik4Gndb0HKXJlzGi+//hUMOQnO/A6b/6Cl1sBvSFT
hZMPmHp49XgiH5wxnJXVQ+3UdQb+UN6NaUUXmKtZ6acI38tT7IQbX9mP7CicvoGo3O4BiRw3GK6U
QEXzDjh5LO4oZwER9fI9HLumkpYhOZCqr8obeIxZZW/vQi39FBsmvWRD0hGUSYgg0uvnKHDr5Cqr
gsVcFYTZKZLZxGlW+k18Z7+n5anbWFoGpYaEmvmQi18pZxJUbDk+QWIsCBAHeX500Ang1LknieN8
aiNclY8TPSYLiqHGZMmn6wSCEL05YOV/D7nhABqDEeZzcawhk5IHB9ABfQbde6xjXYQIhAQ7zSsr
vXbvSZcF3Fh/f5lvtd9bBSEyVTNlfAlNPWEXDDaOZa7xFYNonw9XZcgVyE55RtXIjBc1iYymYllL
P+0Vll68W/h33OIwt/R0JZyH7KwAdfAGIxUzvOmW3MtYPzqpRNFRAgSKZGiCyBbTi8sbcSE5PDHP
ikDu4bKHKU37vF9R5Y11Doy8s9EvIQXNPJTZt4T+r0QOKZ9SA/cMKZM4Izj9HXGjZ5FiU/hmcqAt
nFzffSokIL6fl0et2Ny2TOuVQiq2NxaEt3QWjW5iy/yAqDrgFrpSzuyKU6ZsyGFfkRwL/sW5os6S
69nr4WfUYKWTTmdGWfqiIi4I+i3Eu4ravar2z/vNHvEun+q8FKRUnD1mz2wRzmqm2vbPtRKm3G9Z
DMJ1PnNynrXnsL01Yw3IcakcLhRmR3gffhZwhHcMaY2iLeoWZsuP7pByBgxopWEJ84ocS7ryv4sn
5nlYirf1EJU3CYHVQRqtUqW2ImzcOqi/YB0HvyC+zZt0uV6M+gQmkOsrPd14OZuqDq950znTcG7s
1Edh8oP5nEVoA/TCMcQ7COdC9PbQpGxduvRr1M5u242kDnu55Jcc77mMseng1robWCFjPQ6fKy4+
fXwtX0y5uIhL9RrwLqTD6J80wNGnJ+oZPYg2B1IPBX46YvVifSYB3q6t/nw0E0WhnYchKdyxd1+6
TgcM6S0u778EehY7e4qFxCRof8h5PZG0lZQvu6gkfrbquShQ1nKbLobYOqJQOiK3zhxhma+BK/v/
Im4B5eRG9zowmz8lpAFCxExawcb9n6hoEFcNcADToHPtvacjHNav0ksXJNNj8xpX/Map0odDdt5v
Mj/JVySjrT4w/oZ/8HQHVK35REIQbk697sQGuQyxoI6Mc8hm7X5RXXoz/aHLwGYwTddAIPaU7WGT
R+ddbgnrJoK+7W645fTd+rqPfrvcYXgJNdIRIuLbOFuU1eoJ2KD55pp2RxNmjYSHHUGIOLIxPOPg
663mZ9jH2CZPcNOk7zHSXqc3yHT4ChV9CtUOeN4O8hdHoBlcLn3tKXoS1HVopL2sVnjbqmL5MxCQ
/ytGNu4Qzf1/2hOMA8u1UcO/D/3n4ignSb4D6+Ob4ptBgvtkugwsLG6h4pU7K9cc9Xazu45Y77P6
WHncLee7YYDfsVGTV/qVHVT28ZyfI+XjHMemftLd4ltZyNKv6PFOGLl52TRuet9czHmQ1s2FXCHb
DulLI1b9IUncTCtFtjqS3SiRSfgDzbtKvC/PLHFHxJpymi65X6GFECLwe4F+gvV8RKrK4SJeXmFx
uqKVVha+9Mjdoj/YroW6vJZacEawIOYQgju9qV2qFermlE87lPof3FFpTul0wzCCMSN/mfZeDl7j
/C9A6h0Zbh96uVVnp5eTg0VdoEUb0d3l7dYH7Jpg5PmHbl14HZ4vS88vaQHgrKbSKwpFHD1C5H+r
aa7FEpu+jiIdpgtqvHoRf90lPtKB7mIEAy95RmsLcPkz1/LehDXil/AcR9ymQND57wRztlVFGGfG
mx14279/cFYZv903UvjY9VzpF5N8dWIA7MExmeXNvpRR8LOR9CLR5UTIVDl0Btn90qsr83ocw8Mm
ReFs4tFaPNDgfPHJU2pTzaZ+Vo4jC/nRRlp41ZNSIfVOlS0w9L2HClIe7C/8+IGl9Jt1jilESowo
fRyr8nvxzyk3+Pj4n3pWgqJlYj+pI+VCUKpS0c483pagOcczigBkouFP0SZZyrop1fkE48AAh4o0
2cdOaufJ+F58RHFjfNujP1PAH8yfBFpyjfxOgjFKeHfsYF8+oz+rEeYLl0G0XUHGH4p/FBMPyYLV
mZZiDCf/q5rddsNDzFG4QIJ3pwVdJy2j5FrNua8PvsCnbAunJUovhGILfBfdElE4WtugZ98ai7SG
jpstQoPmod+kdCgB/JsbJ6g3tvYDep/1vDVjggayqwEuLKyFBo2toZD5mOmckcXYyqXyCs0BFGKs
PbzLwk+r3vnjjWYbvPjOU5QOYQyKCQfVptIs2MkPUlLESBwtuM3geAOqcPshXY/fiCRdNdqqFnyh
qdF9FwRJjlIyiCU29XBzSETcVTStXRtcHsv6KJ+Ck0WY0bH9a+H5owwPZ+cmOppVrDI1x2h3cM9S
m+engFonDYNAk3SRtY0bb8WNiycNnvScp7fzutvJpgyFqBa1hy2yRekyORTymakbP8NEoU89b8gV
9wfnaFH18Sfe64zGlBr45lpILv2oKkrmLjXfN/nhb59qAf5Zbr1gzX4HSV0cBRTRPPwYWFQSLgDY
lO4dhJhqqpnG2TNiYNAuUfuOhBdcMxMgWViakPCXhwqfZ3Q1wpuBZvxAz4CqnbnIFML49ZbvScCI
UpmK7Fq+dpFRXGHAA0NNeMsIq+QvpN/+PFdGldMUZlbvy/7+a8Co0lL82TEaKFD7c0eVkvg3glgq
jDBFmXbV/X20hzfOiNQK7XGZjqXmPS8/bfOFUwnwCQvfqwG4fIolJgMyP9nqYtuW+FEIN1VBZpzq
TcyUj4PjLlT/6/SmMoitLbq0Q6Ses11rvgrtdpAG2HyrZcZRNGov8VvaX0UAWAggGohKt4nVMdrN
zNHkCr2ZViApJrvlUQBe8oIsUu11qiKu4AO5hZCq1ajnwpSUBm54qAaUmXzCephzzC+lOcSrlMsr
bc02uVC77+eF5+tlHgna5Nxa1cDU0fBOZ+3Hm2NBv0yCni9evRgoFlpM6ZgLg83gYANadbdM4RWJ
EBngNR/9ioDkZ37IGukKN0aJ4T5TR5RS3X9epghQFURehkKLb2pzpRoukogEk4QxD4LxxyhwGkVX
nxRA7IWeYIZjZHNCNl3e1zuyLgYmy247zykaMfqnBJhPSWVErefDLlKgbGglXIoDgxntPTi4k7f6
vLZHINn6Rkm50Gcfs5tlpd8n4S5WCobGQPslfTnStlEiRs+VCMQ7BFEiYh0kbxIvbTFOnWytMU5L
bY5iX1W3ey2BzUE2nReXWerrqUrAQ+LG9rMA9/Vvc+wUJGXqz0h8WBVJ72u4GItoa25MnWot/j3E
E4oRbPes/gRv/fz6w6aF3srZb9Jbpvop4Iz3Q4ky0EN9uywbYjhSy4vgl8YuMT0r6sLH9Rz7/4P6
IojuuaejG6b1k9gl8XksqHeFh0LtNtet5qh8Em9QICTBaXyGWvH9dkwITNpJRpvGXMRo0wYWbcKf
KsorXJav/g9Lm19ANlDdJKD/+7KVqlhtuC2CgR5ZIah/APGP++LCoHQiZ04a6lD9mi140eDaxzap
bJamLnYwjlrkhLIlPop1mPosAz+jaSFSouAsefTLJOGvZqjg2gXEYHZ4+MFlDkpQ7Fkr7mS4RaMv
AtwS6Y930Yx3SovNaNarsB/dqdo0Tj5hSqcbbJpXkVfgELuQ66OVpVE8YCHwBRWUZvPsZ68fwt5v
AXXIs/LT+A1FrOurnGJL7sn//g6MwHuJTx6w8tiP9JGO12CF7UJbY/f9Ovx9g11SYvd9RE2x3huy
suNQX42qxBIwAquNXgiJVwid4wKwmVxrpiE7Z3fxWpGeqGV4D56rlAr1ZAlTD5mweo5OpYQuThLL
bCHDQJQBo9eQyy2XEAZSU1TNZj3JUbzbfMuvj6YgwVT4H8TlzB1K/3uIXlcVOM7J2WJ16YH/Lvwd
oDCuHP1FwfClWheQbNsL2BSF/22d/dWxckakgdYpwSDp5JbOY6X9yF/q3PmH/52JsMteg3nNhDtS
RF6ecpda0BLkWxqgmePxWhtUj7pqlot0uqA0bAlI++1P2G/OMF76GNZKjocD+YZ0X6z3nY5x3cn0
2D5qnsZ9wMq9xSDOotE2oAatHBuGixFgfmTPYQ5s9ceDxf792sblX63Ekjj02t1WXHh7qhwpDFSO
BUahIY70aWtmnG57xDfbsrsTX9oJLlc9+zAwhf10CBkE3IU5FzkR2GPb2qqlSO1c79MgD1O0a3Kt
Nbog+Cqi++pSB3GqASJhQAYqLDtgthNEtrnZ+LAwHKzndBIj5XmzrfUocTaDPfbEDM9kCs9eSUs6
+Ow2Setm+dlXYlSloPYS4aCc3k/eCUdGDNf0H9vqephj6xWO+E2qKf8qnLQJA9003yYcp2Rvaphk
NonMV0I7cjgQ1ghNRUpRXD0P+GfaF7eVIq7CerA6gcNpfAWeIVc7v8Oh6fA7W1GCCg/sMYvusEQU
6v4XcaUixFh5W1M2IMxO3cjkL4JLXtMRKVgTbkwFBBiS/WlUoX9eVGrDKwuIw4ACURS77Hyw2Hjn
Z1LhdvV38xSsJY+J00NReBmlypUY+Bl0eYqwoYWGp3QD+Qtyzw4WAV6aEyS5piOkaDU8bIX4sbkf
8tW+NFea0lxwl0bAaQlYG+N/SAAW4QLa4MUCF3Xw+VCXMT7YQlOsw/uCkXGi3zWNfXr6UQR6D94m
mF2j7wSameX0s4f7pbtLJciIXBFH62clRZzBrBw8t8sQ3rIWKW0mxApdljiqw+lIbImK1nLlzPpu
o18CFOfbDAw2G+5z4qa7CXd0O7HymorxzkRcAR5qBi6/s/coe4hMXJ/dfryH6yKDz4PBxRVD1sav
e97krdxXhAEAFecM/pKyjwXONp0wWVjtG7+pG5ibJTQXVGoSpfrIvp/daxfSu5hPXwUEXGdF/ZeQ
EHraVqokRwVB4j2qIumCLm4ZVw9BPd18xGaIMFyt4ySsOpxy+eqW5cG0OfhnKjjTeNZZiXauKCKw
Fea0AhGGhw3TQ0K1DoXDZq2tgJ7uXo5WifVGZOkwfj5b1CWyPgK8EljwPVtULpyrLsUXtb0dEq3x
IKUQjltwJki/Vgz8pGY8KZhdEieS2jcIYzCIhCpP5C+Eye8IxhkFw8SRWaAcZ2Ex5bOP3fLyQdCW
nFHJ87em/6xGFIlUXBQuqmetjS+PijifNxEkoV6oXl09dHE+JGsWLkYqIeuedlSuEYRS+R0nO0K5
6Im5YfaLyABnQmTesGNKhbmVFqoO80zJMc8jse2RHlwemz432OGNYn5wCjOLwR0YvzmYWWLEubJ0
pflYiCmuueHkf4tMIWtw3kGuxyeDBMVq8ddCP3N25SBL87PYc7PvIvDtxnLq5JizGtS97YyWYR7z
Di+vuZCGO1M/J10eHHWv9BKYnhCelgQeYPvsSvz+jzu5bjjDGuz4KklvhyJURoEZaZ48x9oCl+7G
Np3GNsJQ4uNpg3NvboPWg4Z3elIqV0S1UhPuGviGDrh5ZjSjoZ2Uq22wrVRriz2yTrddhs998Dri
LQCzbDmtG3N5EwfxkSdC7/+8y/6EPYkAydYsvodPrSKYF2ZgXNafrdhbyWnCsghOs4snzxsBi5ES
I1jBY6IgsQreL9th/Xlkwdu/zyR04Qy5TgYyl+BZIA+RTiol0Tmjztm40+CCYjLOIv/OTyOgvNWC
nCFovQfRILbxYzb1phpqbansUjL7q9UUaL/Zo82ebh7sNIUrbMBohapZvnMZoz82tiAFXJPRhFWG
CfyaIdc/uu4OQj6caz4bVOo5VAL53EeDfEDpEwB0bAafj6ncZU8tlUTMNtQq+pxMyvwLk2VXSp8j
cFZHEPhWiWfOMDaUiA95DirLpGBvZCkUKxVJxIPNzZWpQoLWUEWm97EJ348StvMO7DbSXRmjvX1v
nM72NFKz7+qkd5py2XSN5Gu+C4jxaXpwmj1DFt+qrMXYVVuH95IeEH9KSBU3RhrmMMCK2JcsKVFs
GJfvAJpQ9+CXG6jzMZEtD7uK2qGPZXq50E1BCSzz5vc7g4Ycndsa4SgF2N6bWid36zb0jv+WL/ms
VthJ5/Ldn1Plt6FDCugikH0E19U0UZEVEsfQEGY/vunUFLAq6T0dKFolc3H3gitrPhzCgSTuxUla
V9/tq2imFiqaJGoyharBehOt8fTBfx/ceRIyPRylft1Vh9uC3JQGmrG0xe7RW38tfKvMhiz2BJPW
q8jEQ+fs4TJUO5oXE8oOuctYy+0f1zkC/sU2tX2bZsPW2oSY4kA1n8GIgb/V+YkukjKKIue45m/A
1hA42Veaqg0RJ3UsDZW2W3xwqr5gZ3YIzl96jyMkoNCX0h7bgM2b3NpwVuJqGGxzWqGNwCOfgE6r
MMLpjb2dXBXfTftRTlO4mHK+xVydzaa0vMkmjIOtIZrQxy7L+sQ2kX4nq0uzzJZRQOqtcwRAPQxQ
Me7DzTkHKSWA/zn+fXq9L2ochHR7rIR2FXsbqNRc8tbqHhl7JGQiu8ejp0yFJkdGGh0ZZiUINdg4
vDmzafkTXvTIU0ps1q/8wepCKevHixuSztC+ALRWRpRx14rhpo30tkVfTWviem2eIa7YVab9f2WR
+Sk3rFxCl3wCjRNmvz+dZ7ZSuyo2fVS6xqiWOe+IM8oWrLSN5MIoGV/lXTig3iGMNa9clZwnjefz
y2mgG0z8NiefQk8qla8o7itrWVKVvjp6yOTDkRwwBXgPcCu6a3dNdvj4s6PEv9Ov02LUHIVoUDxa
bcv5HY8m1t/Ia58XFTBEMmfJ+WgS+8d2J+U2YDiGn1SYNliBMhWnV0yejNtVQWyONnbEHhOIOeHU
jbS8frKe/34ovvvjOBXRzYqaADhFJArz5+YfcWCAIxYdh/X9yIbQvPEmaRMDNQKXojIrVkUfLLA/
jy2xE0qvDSgfN7l4Uhik3fm2mk2TGmHAw/H0rD/h1lkH32cG/Jry6EnybxgauC5yinC4cn1ASDFz
/dS4EwnlLgnvv5dEIj6xXjP25bNj7RZPgSFwSkK3J4OihhLZA3R/ReRQkZnOvOF9o4FP+ZrvO9LM
01Ux3wjFIu3AEgpiiQznKnq4cCdC0mWzLEyU6MsT+JhpDPxLryzzMJp5DdZ3bY1IQkQdwpbUpWvc
WRPZdbAmQz9o9Sx8zry4o1Rl1nStpjR8fUdigz1nPBmXC0l8qpjoptf3/yHb6RAVExf1GpTN4PoX
HG2MNqvorJUUaJtcHSUwDWdaks+xrybfuAz/W6sCVJi2uUfuMjbn95vwKXqLUIU2FRqgY27cGKQ4
htOiXZRgjUbVrZsPgJaKNIZefuVnfe8zVzk7m/ZaYKH0fqbDCbrch9D8zXRQcnoHCYw6kcd0gJXZ
gK7ONsik3Yze3AxLVUsbQK39hU2Ck4VRZynJZBpP4kxNNbMy23qzYnmf/UuKNWyhoeSjhWBy0uhZ
iirSWxQMA/v26korNjzNDhIbVx3S82Fg7t2ci+e912A0GMlkpWY1ymIdziwMWUu8+tTqJl4YM0VR
duAEFUfspufRaKY5x3WbA+plnPn/yigj3Q3TxlENm0HH3ledi9jMAeYtFs+INftnbu14ya8Ko57X
jZoE5Vnq9lwCk8D8jCBKr+BFwzC0dR+9KVH0m7/5p66sSHiv9XoHeA184ogYfK9O4JBWNZZsI3BI
VQ2AQDWi9pQUu1svkxupSRZmZTR9eFGMQAI/AQIPzHebn5nmt0ylFh0PJx4Oc5u2lEhrmfEWyQyb
Zwry1W4cycsaMyc5VXBfFoQVVIoQfTWW1cETJjdV0F4lM3jsHoh7X/YghhSl1KElA0zbTvnBoijh
JBVnbjmVmdts2cZqCpD2AQEqIHPhbEAFh1iiCSeLSIMwcHuwZl+QOABR0H5YLzZ8jU4IAGgW+IPi
S4vg375XGcyGIe6L22tNwRbhSHCd80qoNO/im/an2bbar87LWgLeW0xgh3fL9pBKViIejSHCyTYv
QLZu7+c1p8yXuEy8iLxcJ27vmTaPkLLGHn8HEAuGN0N6cOZ7zPmcFzUZcAUZZR7OFEAoQO4kdfvE
PQks1ma9vVG4vyfTpQmklKQdbTr1w+LM4J3jMRtcDEOcgjs7BynWG8Dqhv0FFQ9thY4+LGZHdEZO
NqJPNF2p4Yu126iBcZIvir3wAHdZ93ow91aX8iKW+hTJi/+u5rufP0L9x5hxEqYIvboUSh36yfHk
FK1I/SNWuxZBMDp2Uj57owghuiPCLND06/llyxCEMEAWPCtrMBKGxlsu7pYUPVILy6IQJoImMnhE
ymD0URAT9i4ywmez9gDDIRetZmj1Q0sQmDgMyzDI25tO/r8v9JABixhXt6Q7WbJD8XA/hzKYrKHh
bbq2IDdH9XPiPSjZ9d48K9/HfmwErdLSXOEZ46ng0bwKxgVW4JoICzrq7GxbkTLbxWrKV+QzQpO6
mwYzHYhQNARPV6xSLz1AE1yMcI80NwAR3rUiVFqtMMdexgKakv14nMoWzIxGvMmzjjRNrYtjo15w
SsrCPi9FJTdHHF7XQV+9w0UOQyq6F4jyDxsc4h+R1gfLIDigsZitNx8/XggdFgjKN4oBFExDWgTL
yo+R1okSDRuXEBI5EsS+8BbRUKM+3eVlAHE2xZMH/OMjVaDpWP1DJkvOEqAExAm2RAVZXH1TGpLZ
LfV+L/vy8Jl7PamDmj4XYXrLp0z/afxxuPNlbmFKmVaQ2kg83cLFyW1V0Jf3GX8YVAK/Ob4KMfVF
IxbmPbITj6YRlz6C4GMxXyYL2qxYK/6OfwgRIMLG7xhYPXpOp/bQA4flk5j7LiLN69vpq5TP3C4e
EMUqdKEjrchCHtnafRJb2bJ/th5WFO+m8Nhd2YImcDgYSj8lEv52eYbtUI8DVoiFiWRzYnNxwJQJ
mK5pLIRkJfYgtjTk9SyukWUguulrhwCujZpEmYqglr5KBTPyLDwObQFSlmLcEW95xhpmL06Ah0l8
lJAzwED+NTjuKizZU0ylFTQ4zPLkGc0NDNibWnG3Y6k/LA7MPZJCbbfVbhoPnWOW0iFelzQKBMqP
4E8B456PAk/0R65tD2vb5Ppfw345gBnAcd46/HB0QFXkfCEy4mEQ5o/kDGElcMEJWAsi1g5KeKJi
rPOMBNZB1GotvHzK37eDO5ok25l5o7xnH8igC2hnOs9GLUR8bY2rkHxm2LHn0Rap0fXC5hEarVHI
ifaWLbQ9TKfS7L+yYwWTGJfi2Tw3TLyTZjyfIIrE1n+he1SH+cFrox4gjZ+rO3C6iLPrdmmRTjHy
DALILfOCYVNKuAHUR4FQUyh11B5IgGmZCpMAtMTrKOdrZjGMU0MDy+vziead/vcD9sTk2LSC44xs
X1Jcy2SC57kDlGMSuPaibjSxTD6h//MPndTRoIB3SYpcWXNb6WZq3bzWbM3/r+Ih80N+jLzg9xST
L1WFL9dtG58E4wPKoWrvI3wkSfSLLxe55gfCbHyO9R+dYVQ8QJF4EzRsx4bKOnQTLEQeyp/FszM5
p/E8vTO25dM9VaHEEbjYDA4gDDp3dy/zni4ydWAnRm5EsG6ojdgnIiyGn51tGkD3gq+7xCTNFvm/
btFnTpN2X/WbpTYui3NM6fWhrtsrorvNwAUJk5TIG5LZ0+8kgBJNH+H5wSIGQufHnxq4VASKVrvq
eVgRJOzXAMkyhqnERo8T0hj0/KgNy+jQIrzWVTUFesmYrUSOncYo7kYfuKZGcM5R8HvcKtFbxD5w
QB76tO4TxtCnZyckhGIEWCF236i0VKJsg8KsHpfyK0yGNzfskldwZTFhbjVwrXHWOW73p0WHng2d
Nt8gJ7CO5x/HZtXsX9oegDmuirpCmpDqmLkK47S42YcHvkFdJdvKRRMM0n27NRz+GkJSYZKQpY57
SyilG6+drscLPLAx37RgCevjXOwImj2xc4Vezc0oTqo7YlpwvbFs7rZ/Gw/SIGA8mtSAzhcu4BdC
Ef3FGrl/DEZo+WjJADI5RyjxXLUkg1YDu2DUxV2X5b5N+rCaQZ+pf9Lrjh+d6QgKh2Dg71eQluDE
lFpb2NLAcUav8r6h31NcZqA0P4x0AMCsmZ7CBIPDT3ZSwUcp5EiYISFK/OvOv6JZ8h54oTjdYHd6
qfJyrOcVuffcCSPr4TFDsIo7/OdKPqr25/Vn1voUWWatbE8L6gGzCSxzgNxNQ6MCSxs8Xu9VKjsB
sBR+tyMMKMI//gkNJVAqeRYTqTJAQAykW+CkeyEwjlkw1vfa3J20AWXBAcX3zkP/1MOfariGbQGE
3xnrgZVEjSf2VjueexAEMbJydeZm8XxhGy5aeMsrh/QdkXULunHZ2TTaPvvWlBiYRTV6+3gVx1Hi
bI9eVVjiMXHteNfJ3xNPRPhTXQ2eyz+/qyyxpt9yp+13TwGJCfZPtNuI2oXw6xKbtI9PCealMHpV
MrxdL4xTY8FnS1tHS3qSfCMt6BC2r3PYFZcV14M5UhvHKWKtAYcBAUNDRyjbNtyGnGBlFqiQ6d+j
Qb3IsunWXxl8RlqoiV/BGHKDTDzQhQPFzkTzd/xqimeiTjSEXjFMUciw6lTbbeRBJS1Hc+AMlYow
TEz47yZC5+zyYaCAT+Cd5vx5C0qBkMpRRIln2cgNS+OUHaX1fGfUhpwBGdabs6iyeKrSQFdY1A4C
UN0nINlJBKnAQzEh6LCdKNQzyMOtnTUfgQQuSgPfnTVopXM8xh5XjKdO0Rxofi8QGpPmxpu7ipGt
CUkw8rDeWkOk+8aPA5F7cCgFJYrIYfWzKGRdfMPlGuhXo16U0ALop7Zvvgz5uOz/uF7RuRHsULJK
WkMNhArsxe8xO4TAmZe7S/S8SJggrB+3giLSK8pX7Okp6uYiQo+Rlu66CJlX9v0mwpEZGn6bHCde
Drjp0NcWfS8kU1ht1O3FurMuB828ANUmYIm8HDP4qsIo7lIfxASWLEDumtAMV4P7QCdwZv10XYkS
CzvWXfQGmMBEswdlDuq6QIdW11HBhLG2n3ku528jO3YTSXk/gwDRAOVVxpT0PpuN0Az0nMN0n+HI
s2udw0I+VW176AHc3lghSdZdkHuYKoK6Ylr+RvggvD57FB/cxeXArdIHCiyAEgW0qiqwXRs3/f0o
FyEVs79xreN3paI4wkC48FzfcO0Uavy8VZDs3WIVu7QtZn5J721MUfi6klV/cNAgKwDMnM95RL/u
pw7llarDLrE4Ly2plBRHSxL2Xwl990iFy4Xp+lMMu0NN1JWRGPc4LqPB10lDeVU+msjJqV6EYznq
ouN3VLOxcEwpvQeWEE5TrE7Ez92Uai5x4xaBymGQzzFO9iAiy1AET9DVc7h/60jhdxXRK1HnDT/9
CkMfWJNpenWAVD9noeUHKoe5V/bea++qoUUyG1vEZnI48o2uN/DHV6Lnte0qH4wQwZ9+V8uHTMHP
WH7DOHrujuyQlS0Qu3Wc2ZyvCR++akBN7DQUH3nuxjA9+kBhsjATokhphgmT3TeoGvZmtk62lih/
2uozDkaqSEzN1bqQIGFO5SMd5lNWX0zxbIE/ryK+xbwta19Qy4PgUveNOPWKu0D7xqUwwN2HPiKt
knvGUzvTk13r9lRR0hxSkfrxNM4aQv9ZizlCpCP6+Uoc0AEH5fG3yF/8Tw72vY/z7bDmHRnRy4aQ
OsUg23PeywJ3iddlrLKpJAbSot1GisIZZOEGqFHsQllWKxZbsbS/H2EQavSvl0TUJBYPb3LsyV5j
i5oYhwbMxYhRsw2RWEuT0c4u8uY8PmM9R/dXddr0L76lrDZa0YkKoPweZ1Dsc01SdlQMHmzHFJ2u
/YwwMHjXgoIiRPAVcKg67pHxy2hh3qSW8sR46o5NRF0RRSo3y1fUfjiCHJ7AOWNI0OpAW1dapc4V
9we3j2AB/4i4h5dDjCyOp88vqstwO0Rve2X3stS8WCKe88UftM+5E/UapdAGCHuwW+k2pHmOreEs
1fhlsNB7hT0FFaxSmbSpTzj6aLZj5D6AmQ4O+Qoa69z8nPtuK+pg07ozOEeCPSmhmOWQJfnmAagV
bTfiiwNIpxjj/BckGDgjlO33qarTxCrzDcgtskZ65Mw0Qm+ueE/d6E1es1Kq0S4xwlLt7Bl5vgsd
AyZu3wWBBoIqo4Jjyv447UWsbT0utxCbFO6etZrqZ3F96larQHEkyv6AWGw1ye5s3Wl45lEa78ZP
fEp8/4v6Lbidu1QSo9ShIJULyZVvD217iQjS8lkexLvDi3yJyMtlWPkte49vK96zbkbX+EyzZgCB
3CuEZNv0Z0/X4gUk+D1OEIEWZHpwNYf2aG+fr9kBmFrOAxctu22AM1WZq6tYIvsK5l1Dso5Urtki
JYfcJMBvb9mSAqyNwKoEGJNJcIcmPImdFwB4TvGw2yLow3ztQAzpTfqVa0Deqq7WeP4cSL40TAn4
0UDBwgkL88zIsOuvK6rpYB0ZMdeYJmhI94J10cA1jSGZgDSwP0bSirWTZqrkCuzdluLJa6xF9ivu
UeS3IMNr1wnRUnDhyXYH5tgruhKsP2lOBxLFfNiWXUP8qqg3ovghO3e6vDvHdTWIHRq6mkqYGViO
JLqPxoxu4cRO0aSLthzBoPbLOXe1eme3gwj7VZTQpCCOekoSl722ql6EN0Bw4LLQfb0fxrF3pLJ1
9eE/JIKsmAvnEuCBfDsus1CDcHAu88EH6dsoOBc7hPgCOsVTmwO+TXPtRaUQBcnMk0pgPy+ox7uu
11HOlmbmB3weCqWc3jsgliLKf0U7Oq6evcNNZWM5gx9EHLEIUbsCotom8cjCYxlyHeVJkYH0Myml
kIZQGN9F1nXaYcW+hTB5J/Kbg5SBGtJkj0CPuwz1HbIWodeEsrFw5YeddoJVl/J3znWHXOxKCZ0C
JldiA/HB1E28YjqdkCh+FDeC+GSqLG8O+rAcuPGbhptsAsc6PojRFC/+/r/Acbdf+Fr1R+mHKhc4
nrN/YA0kWh0bzirGm9mIcOYVmq2wL71Idonip+M5YZBRxoSCJA72C+cVlXh1NyVTUUylCSvQnsEQ
Y2aZ7oqOgxKQVDiIJvFo8bdxPMKOOjNG+YLNZUS7jUbDXc+35M+wPlbb47mIZ/111oct0+mm8Ph8
Vo7syYgJl3yvdSAYHFmT/+sGSksf+7GJD7nqnl6DoNfd90YEa3FRycKWQqvgGkFOQnZQivBRlMo6
J9FsbnIvIoi3p1rHtI5PInseSbADcDOemJ9pAylI8/w18y2m3DcsihF1RH5gYunnbIf+iK8TqzfG
0VprWkaCWvhivr4/mTHXTmJZOV3auxeGf1v/Nu58Lz+kOnqE8uWHDFrq8DyGFchoVD3w4RsvnMDW
N/FyaYhsE/vhkJndQq1ktFSbeCDN4p4Ryyju1YoCv6E9xAQQafc1LFSYSkz11qfDLu25HWcK13+8
ZYFo5nJXz6eQc4v0pVe0rAbrrzphP4MsQjp3s+xHMG18Coyu20FFTAsOFDG9xaWf8VxrKFH9ptsP
eS+qzJ93ZPG0pOi0CaL6Ui6jHogjUlmJaPb+/Z3Wi9BRDPxGhsW5oMvEhaPHhJV3+T+S3J8qL8pc
pq5eCRfEhEM9/mG6Vccs/1GTi6NxdrXfeUna+yZrHHHNi/SsvsK3bPhHqe+i+0eoG6/peOYhjTYb
0gY3fvH06D1IrMtYfovbZUWtpIO0nI1n/bwpHj2Z6FkPtBFT6hhnXp/bPHaPxTBlSRYtZgRGvdgN
nKXUMSxrEkI0LlpWZ6bVKzIafpdpDwvZpm/9JcCiwN2Dl4iGVCuYa95C83KLJMpdk0GpY2s7rsc3
r22ywZiyPT22E05IWsGzFp6O949N2MxuHqwlTVW8B9emZ4fcCVwQulP2u1ZqzjhPOJgAzcJPVTcd
GlEuGStxeXv7O7M8TolkVESYXxIh5hwcJYGnEi8JBOinay3n1Nr4OHtZGvYvGsyx0hjLEKqCs8TL
dvfMlUdTZScbpBV7ifEWDNow9PaQrs7tlRmZD0s4Z4erEcpm2Jp17n3yigwt6eNiY8Rov+K1hIpC
oYaFc2yPP5Y/MDtHfm1KbJBRiOfBJPmPgnGmt9n2YkAzfYaKxpmuG81LjSNVYnehXBSVZL45IPRy
EPWWAcHWN3gA0XwAYoBsxx25vrTsd9n6w1smPOUsFIpgUnjIbzmlfYFPRVVI/aaU1+EoMY+Bi70Q
jKvZEbM839mPhUclYFW0CQ38kgLr3GOpC1PpGo9s+HL41S53V73LBnhia7w1xcbpmOodI/vCAvAf
05kcJpOSqkQDGUWEOdNBv6T+5OvYy4uZQakVGtbcPIN3UvTyccTt4PbzMhR5zlJEKS9d/478HMbX
PXmFviGpT+Y4LFvWQNwtq94D/1lQBGMjTE7AUkfwySiL8AOYBLtJbOllSHKXYSqbpKjVs8SYbwNX
nLvl+Msr+6k5YcubkullqyFdWni/ZCfeyZL+6zkA1xUAgLTF64DW+LMnQvkgu1rBjGTp8+oFoODc
TLQf+w9bZvatX2PAWxAmjDODHijXnLVfyhzcMTmZn7Eyu/8/rKwO+t21zAP/ksUDmjma+dy2IaxJ
tAymKWw+Ndft8Kek1fsbasJuKCIHxDnskHVEpvJ+miOqwG1IyXR5JDTLRhqqUS84hR8rw59kZuPl
I2huVSygWLHBhv3a1AFMMVCAgOwjRF6dVGpr0fZMZoGvTKeBGPXITRdJowX7q6ZL9UqXPmCuhCmL
KWsDDu2keFvGxjd/8CzYEDnF4dPI8Mw3O4HQy7UrpENprszOmC1oIwW5TmNCzLnJfPA/dlimvJ5d
zlW/gCL7l+F4zfGI/52WsP16GQ3IHRow5zbQrZDnsSXp+W9VEXi1f6UO21H4LJTRNNp7iZijV+Jn
Aw4DJ5JBXShzuwKbrxivvQLpCwv8iOmNk1juVEzzmP5uDZQW+2UxEzcdaiyDsCLsTiwdBnMtGbN+
59ZT3nDbyR16FPuYVg5ELjlofUgSsk7Di75R1ZSnXRcZLpgp/1R7X3wabFlcwIIyCMhvlRjuEEKo
aDjloFaHvIArdSzHyS89z/b2CaFDuUC/VF85OgkpGb17Xzz12i6VAo23yDmXskB4YDZZBlOFhnnV
B8L+9nOIrTJM0GwfxN8bVGSQDl7QQsapB9LKvEL8eJYEA3LMN6lry6YGQVQjfaCwpH5MhY2zktXg
/eaZQYXaqGYW6kgBn1dNpCoSe06Ze37MtjCrD5qxSAQDFwnrZA7VQ2J6IQahBUVPV4wpdvYjS/KO
CiOhza7Dg/YXvL2uFZXaY618Gxz26uxPSVCRg/oqdm3KojDjdQ8iI+dEwOLBGLBm3mvAwxS1Emrd
1tc9Oixz8HPjPxLSIgD+nIacC9p51TXgDDi9DNJ/pMaM2sYOiBB17IHSgBv3i36I2VW2V/62lTj/
83cE8EFoIQU2Dcza0Syez3Z+rWEjEW6KJzJylfAqEND/LJtzUuZqfRK9Ywm9aWkUnrW+R1JNQkEJ
qzlLoEU947/9bG86K7IuSwqtVmBZ5e6cG9VmdvafzyvLdL0yhWUsFVSiqCiaiYtskys3tvcYdn6l
FlBFc3Q+RowHbBJ5ECUG4nb1Qw01M5QuPp8/xN4RWKrKct2r+Jvd0KYbdQSHukipd6QyAdgctOhO
zkGzWhKbYrBir/yRh0YBuWZepq1v/rAt7uKrtBhNZo1JWDeB/z2ORSqdkk79i6yMfRGwCb1Vy40I
Qh9azv3pc2+oDO0bkMRneNSJtqqRDdn+yyeoGcS7M1h8zMSviQOnf1sP4hFcgolrFtG8iiJk3h/l
IXrJg48fLprXtiC3VBo6hIJatAFUD+anjoRIie6CsY/m09VFvndmAT2qGx61+xPgTMJb24OHhw6m
5IDowJYHUcd0rRUTddhXlmW+7JsiPd8aZVV+m13duuG4YvgJoEQtk5HbGnsIyirSa+TqAyEFDV3L
Kb8YXMA1JIxd6o3KY/GmNKK3o+e8bBo8x0B7PRu4N69WX5+rmL2kOobkcneZrqnMpMdNqJhW+8Ne
VWj5NeLAJTa6EDBCI24F1Nze/kBOoPCFgGQ234QLGoetUsjY+8rz30DFFBBZuGDEdhF785qiPEkW
5A0LdrYrYUGt2j5s9kBkblYfROtGYJMzsVisRIjxOUnqXcm//RMIs3XgMXTAzGLljGthNDXe+MdM
gkXMh+fh6So3mR/ohjCpWRjbmdPW25Wt3clFXa5qyNQbw5VQrPlivWJe1uAoFMsox68N1gguDc6g
J7+A1qRi4BIYEbROBv0kpoTvVwHUJJD8SBDapuoVUeWaO3f4FzFJLsiQowyKCT/EZ8KNa/aoHw8b
tQ4ncJjMSXufZI2uq/x2SGOb6LTZZwXd5Vo6oOHk6dCbLO1T6j+vXzD2ybZZW8cljHya5IAUCg6P
96Oqhb7uzuYZsHGGFg7ASmt85Tmqal5IXeiy9DHr0L9vhkJnx5l/ROLxy2HLt1WJzoGSCyLQ2qC7
56SJwUzdbFdHDqoxiVqF3pBH28Nwil1WOOqkTNHWuMbh+QwR2ur9Jk9oWPnWJg1HX4GOSc/qzLzg
oA7TGhfoHG8BeNQq1hnMqbppfzx9IBwjU7/1fbwcAd7habvoNQDm4zX4J4lfegWvTF9mRqbR6Zp9
b/fEQVlyabLSv8f2yTV2/EEZccKtUD11dGBxYxCY4q5T0uExgc6nzY2Y50S5BKliOP3rvj0xL7XV
ChnafOwHLLvBtgxdnsy8H5joSfesQV9gjBfBjsSeNL56Wpr0tW6NQJr1SkJ7j9ktmCvs1A501hNk
RWKNWchZWF8SUFaAiODMkwII3qcFv9xOta8nGcTzRIZul+eEoPl2rdDeWrzfwMXZkhxEz5fmevYV
bGNKjEHBmJFCGT3ifp9GHIhQkbno/9gKFQ1k01xGDQGX99KiaQofak/6d4qzrLSw1FuRQEk/RS2H
vi15DuETq6ogtOUfaBCTpjAq6l6kTIvx0vJanbhTbzVBS01+d017WN/r4nxn5KSFBanHTsG8EP6s
v72phDjrYfmCnzoqRI03KIs7FSLxmREiLw0i0YmrFjiO2G1el3BDgfGGbC7xGM7zTkPRCiDXtux7
uAC4EC8+8uYQ2VxDN3dI5flQOeQwZ2uBuJDFPSJFBQrhHL1cWnDjUAdc82g0CdMPXsqd8hN4ACS2
G0f+epLHek2xV6zeP3sQMesGism4WABMJG1ZUB5N5DN8zFFayWwardTSnUhLgFUBuOCS3MJTuAf8
gQvLQYv192ITemFLuyGG0BbFkDpcLTNIAh0J3WaGwYwKwhVKO0eIoOW4ZUmH0mfKypwBgQ5zsJEd
yOlanSTe6lLt3srSUD0q+Au5L8XMUKaLK6B1Zn0/Zj2sxrKkoCInNuTBiP3u9NgATlz7q72SfcW5
L76IRWaUHE0bLWXNo6jKbPctO47siWt7sPoSDfZm80zqV+jUO5hDG2VFO61kR/dMFLCxaXY8U9SU
VbCwo8CParCnWoU5LRXzOpYlcpwVvASuqBtrRbTO8py3Ady1vVfXrrE2vi0XJiDEKiDi1pMYtZyN
F2Vbna9/j1fNPLwTsp32Ijqk+Chqy4Ua1GCZNUFftFL6DP2Sc0d3Xw59X8T7vumOQXQ8vaA3eE7W
6TvpoRkEvXJQXNvqihVC+4ntptjiWz6H4IVzkJ2WDBEi7RoPxhGt+CNMLjI+g0IsKVRehb/CuYOB
TMVzlMsHB1GP74I92lzuP3qBiMKeLnBtuomJ9lhDA9Lv0AG/epJdcfVn1lsTEiVoDOvt54O4Njea
IlEH2fJ0P6wuhUcCJPNI/QZ0bUqN3wOUQf1VSY8XcuxGcGJPxU1oBPZ5hmy4fweHMyFEfYb3KWIv
ctQmJS/NaOM1JRbk2nO9F+yGqR1B8iFy2jpk/HkYAZsuP2Zcwkav63I/rwXN9oGlFAwYOMHgEog8
efKLiYp0C2AGdj3qKknP4bouP/LnD4MWdpCrUgNdhon1aLmEmdABTJsrLiIh53Bj9xQ5u2Ye+uMa
TwvDXmXBUCp8sMKljHaUyOUL5Pzqy8qoLXFrQeFg34rHDhYSqs87tF/a8Ueu+CklWbF6KMfF0iHp
Eb1hwnfePfelxI0ZQJvPZBv5Ahd+9jGmqPIVbBv7ofnKZDyqoqQLhs8bCjDN01ylDscRVQQSXia8
g0DitDveoQ1zwahmVCivxEaYUVF+qnfmsyG9IlOqLODU415EY72f4YS6lTq8+98OVFWnRipD9ifH
DN7xvEjJVSdUnAomuc6kaw4t/j7ZaLNyOMySrlVrJvolBXAmVYbgt+at5d3l9Rujl4yKNmrMsj2s
r706HlXRSkVcJKi785iqrR0KO0nrtyhQr7yDPJWovrIFDSyu6C8/HYSoUYVP75RjtSbyn+Mu4X7U
Re0ilFVqX0QerJc5kX3PiIX/WryhjPbats5QSz7mz+edCLtmJLcCW0KOCWdB5ocTHiQYXPlymaC9
ltaWaqZk7rEapOsq18bKGJKxAb9txWgRE+dQRjJdDyz4g8R4ozxJx6Js2sdpwhn1RRGZhSEZcXiq
mkybGQT25ZbceW0KfvDIlz12KoOnJ3lX0cXbrtZJPQz0S2xiv/hF3kPGMCLSh5S6uaQMLG3AcHRt
mYGEeQ+01DTrcbbfuQJgXLKoPNlA1HYVT1eWaXaq/TPUmu6BvXUYiq9KrsDVjTZ4QimKHdjj1rp8
LP0Ib6JAuxoO5qHbKlz36Vp/b3bJcXMIXGXiiFetBqQwY61nfvllPPr6B5zB8Zxmb0Z2ZFB1cwH5
26y4BZQ7/iSDSkyZHY79dZAl/LAfeS25LT4mIGK8mv+3IeU4gaUza0z7ySohyg6OBPu5iC/LkOUV
yin9hZKTvxF1VMLdj2qxSySwrrYrAe80v3RGf3tDAHa1cvvyw5Kd7mVJCHAn2NLaY0Xj8tQMp+QH
96NhEt5VEaE6LLtNHUatnDwcCDiNpqxhbalODQZHKpbbHKAYuR0am1lr0ZwkVyifFk+oL8Rwhi0j
sKeq6Sgptc+898YefD8Xe/Uz2BHkx4skMjMlTDTuL7wpI616vNnFB1q9ubS8tmsNv4sBuTzpixg0
yfboBwCnnPyz8rlJ6LIpZXtZMY/PpIA7VSkDwYLViMvgc968ODB1Q4al/9EI03X/8HXgVJx/bw4Q
u8J3kkr3VX+VFseJkJz3AxVFqwyQ7X9pBkvf1AmmBjDLmNk4HKJxUm+jHbo21eZDE16NcDODvhyp
ry1egG2gnV0h1OeQ7el9k98Hp03lnUPpmMLwE06t+olFQjdCJixEKEG7NmLl+xrBoWrwfkuwO0mu
5Vvgx5NRieruTqSYAEBXQXJ4dX9k3Hozr+jKGhXRvFyEWsL21qWsjQ9VmWk/Bj1MAEJooKo2yQgZ
QM5y6lZPUnMSDUnA7bC2F/rjIlLRgZQea/1DSfwP7RDq1MG2gZnofObd4Q81HB2ynjPe9rvIc7bn
yaGcfpxILlH6X+2rWw95kl8RIwIiFtdEqvYg6kiv7PVR3p5p1EyUPoVSgXgxRKEJJoLYMK+ewpxg
wDT1AbrQAHR8h3DIDVool9ChbPgPFu4proSVHCOmhvD7JP0eCx23gy+zz5epFiXICILk0JP7BPWM
5gmActjXMHdZfQDNSJJAsNhyxCPVofkL/J9S//U1jzn4ek3lm3OZgX3K8jjK70lXa85fKjaqkGlN
7g3/SfDYmEsKOjsF6mhxV/xEl8q0wR4RrBUML1wj3a6ddQorB+5M3WEaYjeYwHHcCPb+QHJAlcOr
IT8Zdxx0Ftc6yfLRqE0mGFpgBgKYlkQ0Ak1hIxVcRZmKUsG37mvw1AFNQJfp8R+fc5x7QBeHZBJx
UZ7LeT40gx9OjFE1nTyuvaOp3JI8kb5DIUkWtjHNKXQ1iz+Nf7rcNrj9o4T1hRATx7t7u+mRlCNg
cFQ4w09DTnB+KZAZiKNeeuO2MNjP/VVKoysUlRtUe/G9y2Y6w8uQG+U/X65qBKFX6J6gFYjcFSwl
YRS3kKQh0/MizCzRnHls8QROeWbtxwK6wbgTG9bQcPYUZlUuawLU0htjRPi5Ycc4oL6LXN9FTAzF
SjuC2ZKR4+DC8YAWI3w1jHYWQ6YCoQcQl/2ax5xw+Q4gUMlHgaEA69siZRNv5pYRTT6aQJMTdIga
QbO29CqBqQshvmaPmN/UajQ7+YVmmJ4TA4alRf4J0FMmlVVNLndfwhC89xDPSvG/byiAQCcgL9j9
MKS7Lyi1ndX07dNgFu9s5+7saRwqO+A/2MDOx4rzy0pT65WS7ss+eeoKuJj6CQC6RbuqM29kTEXa
iTGUmkInrpLZIo3sPiVbd2vmAp2BUAhSPyK6nUPxQuwcACee9ZP94gILJVLtMhRLMQqpYeivqpE6
vNSgYWL3BiRFDYPNworRfdHo9BmSlEWJ1gCyAXYfTkEgEqtCa1QRa+RqxE7isqUUsrCFbVRT6ion
gF/3IlL3wJOvJwCf+0KdiATCQUDMzToYo82yCF8/ZPIzXLthpVwnKpR8Hv9ASfqywV9SoWnSECW0
fYU6mgY0PSKh2eOS13kjSFcYGYfbDTM4ftZzLPfhPcmfqQ6IJQ1m5YhY39DVq1l+PZtk1JnlEIiG
+KUu8mF1J5Fqx+QUfJdGfhMy8/WiM6DI/c/6F9N+AU/7z40BejP86DEPvP5MWRqjiDByr3iqDkyF
TSMb4ITcRER40msgXxPK91JMqgWVR4VxX5fCQuE8Z02Sq8vaf5ZCGTQSNCscUzTFYiQpklJIqU5L
jzQ+2P0E7CJk2RuFaoPZ74DMBgn+FQv+iQlpM8oCD6NVJVd7nxK7taw6BLiG41SqDuzVGhwR4+MF
cItMZXlp4nNu2CKMTg6E6A9kyDu1U4K0roaf6Qd4aEO4MxjRgow4Y8Z45ElpxgeDnmLS4mFslt1r
bEGnKoMWl35xQ+Nmi1F65lWSG9vLTRSmEci9LL/AHaOHnB3cS2nplSucNnAJtyynn5GIkJDjS2c6
iTAyrI4z8KKVsODxyWNgTdpnfihrONwpg+rU72wgLh6xUd5iRsHT+8SYAMR+1fCdrAhnlnfAayRk
eUfusjgWNknbVLEjke/1OY3pWXZz+ty7XVSVaLgkm/bIaeXy3mryDDJYwoxHxN3WR10pjUOWb1jG
GAYzokTTPXRch4HTfnQI0XahIu+Ci1Wd53VV0gEGqLUGel9bB2E5AvDCuSgKl34dl9NoQJ6NVCVb
ertYzLhAYsy+QtgcEdKiULelwLSKhvAXlSOAsTkMlE8vBb08sRUBI5v67PaYzmCqBj1/bKpBbJ+t
w0pB7DC4avvy09wCEJ/AQMZvyTKAAGV6jDYFynNlh01eVFeJbSlS8A9P49G1lXNImtgDhCEPcKEI
PzrcgkQJuBz78JkaNNTr/ok8zHB9il/tcGFXrDwGmEpTCzXBO6j03sBj1vJvHz3m36jR3oEqd/04
rhASvi0fBHzt/RDTizDS9McbWRtg/vnWzbMQ42FHtMH6RwgeP0BKSmIPz2cwMlZ33s5E96IFj/yO
lqX64T9B2lOXC8VdMHL4sxkgnJo7xF9ew68ylAApQZ2r0kUNfbUh7xV8L5ZT2NhGtx/wO52w7OtT
yU9HdnNgPiGb2+UFuHW5rA74lMG76C2NYvft4OJiWo5yQSo1keUdCgo80B6wq7OZ/OkOXx8zU367
qj/TjwNkTbJZ2gPnvmwn8ogJEy/2CTwgd6pxdL7bdu03bBrhA4clp6yW8ZGYi6j9SLlJe0nXLZ4O
Htl2w5MB1uAby4xzj1ODO9MhXWHM1V+Y6m/qSiWwcNgpvl5yPuj8ttIFU+RASxiN8/4YAMZxdU0i
u8/6c02CWVfg/mKLe/6etprxhw0zWmPe6+0PEoFSBnpVLbJAPKeiwQGqly+0tq8IrbeaBlIo016A
r9KvM+kI1rOYbYq+AkUDeCs5hWCYMvDSh9jtN6CvKJ6ccy4e67flXmzz0IWItIfdXS7NTNhVw2ER
w4ymXisS32hIj2EsSnmobNR38KysfjROrEl2oOgp/lsED+uTM18C0Mb3siwl1H3sf5dNateVKcGU
CrsV+DENlTfBidyc8Ga1qwVpDGUEiD4WIL9KznrlvfMJJ74LFD5k1PqZZsfpb33zI0/bkMvqMuG6
jCGbzEZ2z2Qg4jrurwVnN3I7sV38NwyVXctNmgsZYbwMk4bRUSE3P6/LKE73YT8EliNhJUYxaVZV
2YhSJTpdnYs3C5xSDYt0H06UEnj5j1iCRAcekDUCwD++hQUnUuCDvQ9Lrp/HkqWMy1PouM6RsSN3
GZ4FrNe3uxIB9il8cyxdcQu9IaTh/1fBuxbB+dfMN1nt4jQb71S9XFKFuW1mN8xGfDUKidZfpQew
TdSl25GVSLtTK0Rg8gxPYubPyBkj0IQnwBlfXW2KKEFg7gsrF7627fBacQ/5u/PaHrpQbcyxFR9G
Eu6rKN9TYqxKqjFC9aKu1mTKKpVoG02ppcaj1fyImSyP/HDq6aObQJI0KhMwW0nIAfntoaK+gU5D
VLJwVQVu5wBgXdXV5ket4Floau+fKTKbmW/fhR98VcdZDbkgh/vKbHM6tyqzmit43VvWD0s9SLHR
ZKmy38rFNBUa2iQGfVEr20uyHMR3xEfbzAuUk3NjWzgCdulKL6I7Tyj9Z+DtqTeHteP1pAORVgKf
AYCUm5nFH0ij4+ohi7B2euJcyKUtx3prYwlkWDCJYJ1zVpqWpWGw8+bmvoRtG6fsw+G+2FIJ3uKR
hVllbN+cxZ8/zffcBcN1HjWumDZZPPZmyyLCERyaLrr/VI19H+EQ2BFMJSSTeYVa/0gTng5Ng3kN
ozwLG4bVnXm/OuMcGzXpDPTS1MfqFPTCbCLgq8x+QA78UR82nvnjygMAVxSzHxONbXoS9KN41UMz
aPd1Znhh09cepxRD1gkoZRuy9qafhx4z1tyWD8rXBLZjFkMI7nkkCgmsC+d0V8oub5X2QY2DRJHy
P1jjToC5lVaW7mzSaTz/3DQCdACCwDu8VRs0Wz1APjwuQs3fFthzoK+DAMufw0Gx/79Ekvi3I326
gAWGSvwFgxoOusStWybVAnNZkM5pZZLqb+qUQ9k5XnJmQZf87Wy7rBiEuCBruE9nKtapn7WA96jM
VKIUYhA08GKo7j48jdiCWKri392/tgYlwHbPu+kwCN6F8NSkQsYYHBUdYkkFXxuuVfyEvpv1Ikky
6IaM55HqOfEmLHEB18ppk6zFlPxuQ3Nb2yaoxVMwv1J1352xx3KuMXGs4VQJr37tgWlhow+6BLid
6HkoA4zXogFjy0dQqcOXDl0+In0YrUXy2g7D7K46DN6yC5xBOZwYqVABVTTMBMwl3gNkT8qUSMEW
3J3o87juz9d+jfacaS9rWDkNhPbLncRMajimekMGA1s8gQJjJCyFxd0dci51+RljqiA4jXd0uZlK
Qg1jWcFgr1k+kRwPs+PkEKmUlnj+9c1TKcySVlrsd0hbHQv6ZA+vjNlq73zQB8YxoVb3DEiU1Zn5
DImX4SgdNJbY93zdlFQRFJ0y/hHCASIWdFbkMJKU9nrqnKNPuk2MT+31U4lItMevzJUmdmwN4zpw
uCt1JRSWgiScNr8rde8auL7pOjtHHy5DsslT+i813c0ROt5v1NYUtLa5mPoQbndBqa+2HNZ8v2vq
JRtoy9rRWp9t5VGI5JRuMtTq5F2m+cz0IuplYIl1pWMLhgDDGUx9IEgJtFAYpICmHBjBOUWHI9+f
Jb1QYSJ7BZs5wfPnCjEvmVGrJYADtqJ3rNNXOXzJfLhXI9J5WFakwCIpWZA/3pTLbm8jggqFYNIC
nQHlb2QYD5t5LXt/pyyXjmUpwnNxEMXvC4Uxw4EwPTvW0iaAYbl45qzYnTrvgJlWd75nLcKsAAoc
xvWjGjxwLEyUEmbNEC8Cv62n0gdBTCnPMtsHZ9OZNCRSW6mtlgrpKVm6L4DqHgz7iYPNjLLG/Dv6
NhY7uDH9Q1N4nHEt94INV5yOXk+HdK2iIXXnxeHVVtzJ5ZSrY2vlCU1HmlNstJxNi+sE2AUWs1CC
FyqNQyieDoLx1dOyhOTDU6N4Plvk0lCFdIEAV0w/uI7+AjIAvnaypZDkycqTljZ2NeYxzZZoh0No
Jekcbh2PmNsb9NCuNQ2fvqMXAcJPyZx3VVh5xGlnBjlcOz/+YqjLnFsM6fF4nfZ9Qa/LM5XHriG1
ne3Z2b0CROZChCSF5Vq8LwDXNxRKaKj55cc2+ONG2eIOZ9Oit8Se02DoY3v5kEJQFTalh2G24Jif
xeMjcAEAWrScS+4NXX0/XVwPHsUM90kdRvYoLsSXCGv/+0Flx9txxHXoO8cMucqBW3KX6w4/MW/2
UEm5s3Jjj0VC1JBvlusTFsTaaQAAzU1vwL7ompr7MEgf7CMtUTsp1ffjlyEgn0mjvLWvVpJiU7Vn
YwIis/ZpY3xjMLMGT0Mro1C96VluYodEFoQiDe9/1Mdi6iY4QMXHSTmjXraL/q7Nnk9H/5DQj0Vx
q2UJJf6L4o7nxoF/GzgiynBJL9nye4xtRIEN731woyVjDVEAqxUy6gl6TteKY6oSWdzPVhUeXRKX
ZpUgxJYib7AblUpYy1QSBD76HFBaMjPLFgJOztHrP7mxQOJpWdJzZSrIgSqY28+h3ITJaM3qNzuW
0GBiPP/bxSZh8hEy9CmT3yiBvnyi9Uja8r7oBwQkOsUw1HeHnsJi2fhWox8EFlkLEHttWJAXrdqx
v3G81a8l4b/TZkBtPj2aJ7eUfiDLyUXMSJhKaG7d7/20MWqYPwTH7x2L4TKHEsbXaLj9MoXah6Jt
McyODmugaNf0yG/Ud35sb8a2TAcD1I0Kw05alZJB1g36ZOd+h7N4ySA1FWSZoNUYB6gRFBI/G3ga
YAht4q98xWEICet5z+g2O6eyC8qR41g0ZJ2250I91nXIji4xUvIB/HhmZ1Mtfq2GKoD+pi+qYZN0
F+g7oRsJz9Ih97iB5CCIX+NKVa28cSL6Uq/x1v8eKR4biaRT3+gZKOPVG8VnKiOuMTvKTwr5Fm1T
uOtjbI7iAZmx9yfLsaKmyv8aYtT+Tpn/AWvwSNkbDUFfF5UjO3W+XlFV4kFuC9aD2iCqxenspUsd
o05atMXjlg9zNi1A8xWyrOcXSDDlf+0tdGfE5d7dQt7IgOYfDzdtsKvOXS7lVT0ndNRBUHJGgwkL
g+KDiMGbiZCGnnoY/SDSPZry99vTqG4nDqgbsEQEoZa7RxrMuNKEEAmTJ4YQhOL9jECpLTRrcsnL
dLXRVydIodgMFos1wiT9Buf7nB8ksL0tIZIa2k183QAp1Gtsmn0lGHob3XwAYhw5cGRm8lzhJgtQ
aCCNkmBYXBzn0egPrzVRdEJotolyp2vGO2GBWIoK80o5F3fh/S7oGT8tNqAaFSBkE+ZZQP1V3pwm
QMcLOJyseEZ6rv1EsXBebCiewDzcLNVdS5G2V8HNl1Txf2/KZxIl/XUJf9DdPfo5r1OHivt5IWM2
EguYLffygHbpXh/Tb0cQ9Ll4ID3OmVVn2yPgrc92oiEQe02cOKPPHCDDnC8yLCnYZge65jy5GDHy
4junIfeOs0SgKwDywr3V3lJk47d0tTh/UpV1q+jmkjg0UKV3WdJATisy0OvBaXeTpoIthjho6MGj
ojBZ3y4o2i/QWkUA5U0j6tiea6joya0qwXkS5Afa0IBwU3olZDrReo05NTA75LfcdbhYd1ik33PK
c51x65iGoOLTzl6eEyd4/gL042GCJen46D55T6eqxO1LKeRUjcNMDQkDf85BL1naeCopb3ayadtc
JTIDSTXs8tY2FZ4lReZCkQpa4Q+P4nsWVjMx2PHR23gID2SMOD2AThcA1Lc7XVyODZqv90xv5iqu
JDD88s+aomaasJ85FXGYeMTFii3fIWckG3cstMwyNRaloUAn3Q05JmP8LovJXhA6v/AkNkvppSNB
cJzl0cG9SKsDBloHc5twg8VWaEDDsy/j8UzWdaMErAvspcxcJEZfAfmSWSlP7uxua8zOSQkIA0A/
cEAvOcVt7XvnneSB4eaXq5Iz9YMZ/43IDbIJsEtNmPHSYS9ZfQnQKMoJpDs9jVnMWnO4v91sB247
sy2fQO1ytEvz4QsgWeP5ykaoMzHULZkZz1DNEy2/5kHgUJ4U+9JG37R604JxfqM91/w6cnN62X3a
FZc1KJr9gvoczk2lbzZmCfbq0EO8Bqxi2k2SnO3vysuls4NAEI2MuKm4Emtkvru2PU6cbO4QGM/8
mlEbc2IGcD55qafI10EqdxeoUr20jtfxww6WzEMLsbcr5nohesthMX+Q3joSumnypelAoT02k6Ur
uMyRiSSK6xqQKd9npw7kCR7h1e5sm3lQGd8aADraG1h/+OMR1eKznBaXD5ixtYxZ9K9Ph0wUBhGe
rkcM7/uVpFVbHhkcX9WAUEkMHQnjKzj8A5JFGNjDN8dshJe8nm7sutxLngKeZGyTWEa17cTJU8k6
W2+xnBnXbaKxxtukEwn0Q3Na6ritsBBafu1wgpzByejF+u6zOpSbvf3a144Z5lWgelZ0mCS31OHW
ur0fSKehu3tcMvXEx56Bc3LYb131jYHppa1C1gmN/OMlIvooRWzWivXkIu1YXxocql1Et2kghhgR
2sTCIDtVjXDDhqnV/oWdwW7+L6EKB6PMm++ILY5OY4JUGvyNZoxWBWGoyu+FlmqNqhlhE9OfMlDj
fJz9yWZLHtUc/VPVYkSVgopdv/8rx5aaQ8IvtbYDGj8kGAWgB/K6o+6FHlvpd+rpLEi4v8kdSzE9
BQuHtbrN6WP/kn4DiKwH8vd55D+o1KAle708Kvi7ZiBotoPRQ0au04zboskLSjGOdYh3bptVhViy
mOln13tZk904hS3A92cmdYewgWPcXc08phdp7QiP+4CdrnhWbUOEr7AG/L3vvZbigvJRtLrj4viV
clzEW1SZy6ZBx4OZKpTtRFJT1E/sZamJGr89LxCrPkWmKBiOy5th1cXHIYj8gY0/BAP0DOHBEtAT
+L5CabTKBeVR/SUt95ArWhop2Y8TOu+WjMBwkp/KggUJSLRBQH/wDE+f4O2nunwasr9mAgxj9Nwj
AY4X4HW1aVX7XJmhwvdEvbW6aCTTc54KzAtloJu9Bk9iLHTE7ow34PP7MQaOrDV0SojvGBz35EZp
KSn1uHE4Od5suhr9T9hT1/MXrBmRAYiLX8UYk3j+fSwPs0KU5R7EGJ61SoHJIxCl+Ndb0BPqxkKN
Epn7QVSuPhkJbs2prbxjN7IXe8uPlMq7yJ/Ub7YYeF+PEeUhSMxVAKE1hSAnnBmhzArL0SOiGHSH
UJwpTVJVFOe6s6vD9vdwg0y1CoLBAR2IokGT/YOtenYNtzKxrhfQ23GGFB7YdQYPUU7g21q9XFZD
NgbJ+zXoWIsV4e82au6pXxgbWgjkmxbPiqkoJehB6SUSOF7dNnYk90l/nc8X51Xgoe9l+tK1K9L6
01FvewFsRLdR272VKls1G4mFPyoqj5NCufcYianNuOFYzFOeH6sdPo1WkAISHZtfmx9u6Yxhxx/e
gy5Rsm/HEfH6HHdcE4yzUzGyAAFLZz78Y76fzXA5sR8GEu16pSU1vjPRnIC7TttoWlNfL9pQWKMB
ODI7qxrQMx6+NUAi0H2d8ms51aniB5hAMPbYLxCsejbbFM1gD31qR03S7PnMes7h0FBCzqaBs5CK
oQVXB7xWUd3513hDVYBNYirlK0r3Tq+vtPOaRdcWdS/4UQ6mXw/mms1b52xRijX7FATAM/tZf2rm
D3biFyEYDlG+PbW+GDEeBhtUgjedHRTBMoLiNynME9TI3LwrTw9ARm2v1ur6I7qv/I6kKCv0/HXo
FJZf3VP3evTcSnIU1mia9F4fAaUZuaZKoNKn7dRfs5x2bykyEbnV3gAhpYoRyBxGmOxV47fS5sym
zJKVM5OglXSRkdn2M2NOu4jkZduU3CRfxaSj0ok3Q5+TgKQeHLtZF7CEFAEOZKww6bAjsNpnrKl8
wYfr0thNPk7eIBWhG7piQvw1rjzdZDV1fF9j5C7I+2UaXwXALM/A82sJ/6Lljz0mpqE2yRgGWjgT
ZotQInbd03zf4xEjEfmmX+5KUGt7wbz9n9YpqmzlZ47p/+rJ2s/6egP/qQA0+LAszmZKk/Hghskq
l4CVtZml1zJhCoglnxazU0RdlSWMvI3h1cGGneqHg3FH/qXwu9r1HPAvNGP0ZXRmf8PuPBXDaRBB
rcQT1TdLPNSccAVJ8StbqY4DZkDzLMbaRRh4SWcsnLzfgS469YRA/g9dYTOwFUQifdZkSehm81Fp
YFnayBDDXGT6wNlDlONLQ2rde1NTgiyosjtEMpLKlpv5PECbihhs9aU18TV+LZyPEFgSK+iK6wfG
AyQERfxwScd3XxQja/Qp/05I0zvgz5WKVZJJkEOYtymBBCBhkQrE2KIMturmyg1HDWJ6op4Y9KZv
9/qt/rQOMwQVIX6kYCxlr4ccQCZx4bwE0v4OjRe6D3M2cV4agZhGEQ6dUc22DCEeT3y5EkpSuICg
bNmrE1VRHMJ4gZtlnVr6t5gkG7BplU7XkaDjbuDhvJfhrV9PjDlS2hmkTg0HWFOrwl86PNdxDAlY
SG6w2C6cTDBfrZw+SMSko5FQnJQZq2WtRfdtCb0P7hvf5SK/9VYjhi+W9y/FdN8yqFFDuOj+R3Kj
1m06oORHsZSJSgIKI0bgH+J/YnT8sBwF9yk34t0dEZ+RAwr3qVHo26LbeJGJac7Gps9xOVbvQBVt
I8t/qU9vDaBZN1EWyQKqKwcNPGp3Vc4hzHyCLLdsGmYpiZWOkzRigZwHjl023/hhdeoYIvtfClw4
x5wcQcPk7anHNy8KI/xSMdKzjpTcwqqnKIBVuUsGHNbRZ2KBz+AX8o0zfRFFkv2m3WIHPsTKD9n1
lo7Qx69zgDH5Y4qNkrdjc+DcDwJa87kV3ZC6z4PgKp99n9uhTMdFDQEfRVMqRnpuXuL5qkoBruA1
/4ZIFHC1tATQGEYqfB4JCaZGq3W0uQCU/iRh8h8OyffZT138Rh7oUsAJ5+6PPr7vkyO4Vo+aGP/v
9KygKXfBuQ8iNuxy/iLrkPzZZCqHQF4GMJMu3l8ikqgDbKYQ/NhJcHnewUP11eEfUxkb7zlYfg2C
MYD5iQTlcccCaYxpUl3/DZhbPWFXl30MRSJ5eDFIheZ115sbKZcOxktOuvbu1/ZOi+n2sOOLvTEl
57q2yr7NrZi1nKqlU8VsB9iR2Sj1OJ38TAlM7t1lD1O50G8faId3BGGdoiMsdMPsuV4nbSDh8NEB
KY4mdNmSWT4RXLBjyXS3rQbhV6RvpEMf+xi9hJBSwN1IBfxpvHfQJjIhJSToVd+Vnl87wzNxL+38
8filUJQopPQjCP/L7nySWOY3HqNibxBnjjQSOupW8qhyX+5WOhv/xNGUcU/lWrLS9S0lBDn8mX+k
gEZRq2bjPGpw/mbvPf2os8gkPYElqOfnygjkBKd4dOO0ZeZ/kIoA4+KnEbUInlGmj+fhWPiBDugx
3rLk5XDhvE/WnkyvHkzcmHXGODQeSSONZlIl+DbleXaP8TeuxL74BJArOplAaxvq7f9/qxW9/LkK
OZzqf12DoifvhdY/wBmvCmWB/ZEA2T4ZzM+ISADk7we7EqXPDmb99BFFqU6UniGPrMgZJUiWnQL8
BALqG10TOooxFAKkckM/7ADvLM2U15+iBU7qBJHWmR70nKpuPZMPPZPWDIKUygsnw574b3bEcEcI
+Ei2f2dLtToGgldc27o/TssvUh5Go06FIbo1+HuEV8uoKi+jQAwcRRy2wF83lusqpCATuo/I7qjM
gTgw0is6g0uedQF8FEtKrPSG6Y9QTi5Tyre13EoWlI+UfPnuuF08lXaZ+NZT399G7Ac9i+cfDbvK
rvsma1LWX3K+JKWbjjl2Qkg8WGBSgiyytHu6nrRWA23dU32D0qF+4VQqp1qDsy+sDDBj4UZEfs6A
GUWVlUun1/7d/WTsNXaRoza4FtXIZq9vAVqHJuOusfrm1tai2U4orv8OyiEEZ1KGI9wUj9l5Agrh
/g2rjMSsi/ajEbsKqMqptPHK5fzX/hyON2X76gOodok21Zonx3xM4YD4gvafBCB2mo4rFL4fzub6
KGYbKWys7QWdrndKWUI9o0g8m0J0BPPQmpe6kYkq+IAUuPavojJWHU0GpCI1JVaMKgrm8jrrQQru
fA+5sEdGNa25xv0JtIve5l6Cr/9aar/H6hUNKmHmeQ8dIKP0cZZGBQaWKO3YNhG+fNb9pPDJQhmU
27XuvsuQlSI9q4jyq8dnOlzoZd4f+fmnvWIOcWkolroMswScZgQTXd07uCNRqH9u9kyB6ICITNjz
Mg0s1mY1Ret0ztmoiWt2yKftFkX77FwDlCNMBbSV035Un47X2b1oDsci4tNT1vZN/obm2ELzQJjT
Zwhh5IINivsQjPGgnH57XMVw1aXmN0Vajjc2HSD8aTqUhAs47Pj/45kBEHlPJU3PcY9zKz5clB6v
y7TfpzEgx1eF2sOEE2tnMFkRIzBHfiwus/Uz8aFAFIUqTjiOhNSQoPvfyvhLJ6S+hI/xuGHUDD5B
A/x8DbqP8K3l4sF4qjVI8bHUTcec5MIk/cZIAQgVQHSp7GHsOim5F59z3wLmpV+ywBbNdxkY00kZ
SXauNnoETkz/1ByF3SGiYa2xVG5DH5ZCTFoPnL4aWc2wR4vAjWlXFed8MpjCTlt8PdPe4gMS4Mxm
8Ao0itAJa2eotlKz/D6OYUvK/51igQujx6TItk3pSPQtVyNX4y9V05V4GxUSQJXToQscGZWqEZ14
zakgC3RDqpOUh4tvGAxjKq7B0IpRuohgiOvxdx5ZVSn5R1rx1CgiyAU9KWyoSoP4WGJYNiTpXiiL
iUWaUVXukmu7fVoMF4iznwCaHhDJe3wzykFKY8CitnXorbFcplmWSW4p5Nj1ewj9YVJfSOYa7GaF
JUzJpShbQRB/pR+O4evXTBYn30tbYvu7Oc5o9vM/rpdAEJsOrJsdU4mCpd3gB0fPieHgCbD259hM
CxPnT5onvh4MdKgWK7nVaoaTaWqIX3qP94gMQjMlO8rcU72dhdRUmKJWazUtsKP2BoD/r6suDcuf
gvCsEopJkmrmEdZfo9PPkLEMYN78ImCL5QLHI0Rsv8Yg5JjwN4cwFwbOZeTVgYGFlEuiGbKyZHEN
6uz24ew1Sqcfbq5cLK72oBMl8MsdZkMCNqlwYERy7XgvqwlOoQQbF6jXboXo3VD2DNqoufKQ5+BE
oYU4663gxfXaZvEUg0OZ+wVloiCI1h9ks7xF+MklGHrtnSUpkKLR9YBB085dkpnCCarD4SLuGpj4
jMt95EM4dKypW54YOx/tz9mIMc0RsLXaQ2wTlRDQKV7Z2He9YYohqgAmgr3HS+vJii6SXqyUNaFt
QCpMFMo1avyaP6IMtz2mDcNgZ29FZbaX5jJmcSzKTIodnUndmyt5zdcLhpDJSUbK95w87/FlO8D9
8WAVzfuI7SApvIFNi1SVqH6uICw9fOiRCwlIEnDxKXsXPUPCDkQZtuaZ2mTogUii+6cctAa2dxj+
Ur64bXtS+O3ChJPSJIyqO409aPqmmTwNUa2wTA1lgB8eLvo5RYDEZmIKQbSeU309I3QAxTr0W++u
uG0RcxxOq204Hs6tROi7AtdpiKyFGO/Wps6W3OJfmIVi6BNtxbpmMFgELXU355wfeD32lTy85Sum
+ceqP1raNQK4nOS4DQkWr4em+XfpfCIBGR9flOSwCpRJ/Z0ec0GIINVYXINMPkGOqkpfx18SKJcd
/w/pOxvTRa4MWR2iDR9VQfn7z6CDkZ7YHYNfwX9gVWES7ZOrAAOo1Yuh+dqi4yBfG4Bxr/lVjAXP
1CKR7GzE3OKYkqVcpOwBo/huDoBhegahhHnob51gXe6uYDkR26fAmhUtXGXUHiH+HzqeBXGnp7Cz
6mv/kq6djGSWZXeoReOCWub9/Vm1QPZ3z7lubQpgHAoUTJw9KN/feWspYZ2pGCIi1Ey54vLrK1o6
r/z6EbnU2OfJBXmg6zn8UeLqBaxZYED821XFWZJRxytM8Qfd0I9iuGzmclxC+ltq6JNNEagf2RFM
1mHVHc4fklwUIyHBceJoth55Jl8RPbUrkBQGJGm7Jpe3op4s2YS1jN/3fCzZ+wjyxq7j5vR6AtZ7
t6XT979EuD8DtdphcaUz2cPhi0ef3VGhiDPc9J11fgztqZhp8HkjC/eblNTypMF0u1rFOCXYK39x
r1GsLQM7DZHTu4VxmiLtL0iDeR6OMfmnzTZXoMm6MENLXV27sTU47N1rZ6m/1gkhDDVrZ4A8WhZI
ZNUYB5mELkRnsF9IKQzamQ1z0IWNco66hPgv8wS3lQOMoen9LdGDTZGV0wckZfQfeE80E1EMUf8O
mCmLBFwyDsipgQ6UbPkos/wT5pF0NeZdrm7TZd47xnkHj4O3F6+lPedTsfKSAT/5pxRKKwvETcyr
wLFo7CBJEdQ4YZUG8qx4t9iODanoBQwImAaNTG9p/Kikinmb5kWINZC+NOqeG18lPLTqoe5sqD4d
/T1EcBg8OZPp99o6Z0R9T2R6ZP2+LpLUEMJK+tnuWDfCNyHqrX0ZjVC84ALMBERInRUYpBesvhXM
jQn8Rp5dD9BzkG83t3Dt2ni1eW1pTI0KhVnUro0tS3crVGLQmieEZ/D8J4dNcNHxTwyKipuU74jJ
7e2Es8fPithEHfOj5i1Jm5CfcTUza32caVDJ4fkHinrKG2ny8VVUyfS5e2kiDgmqP7M1PVNr4P9w
QDzIX5+0we084SUefhRVlYFXpzKzP5ebAchMipicbBCaTDELKrTYhc/K2U8MZWaD55z4PcF7ksDu
qIobCZGBNUZ9a0DILb1mXQhs0v6EeGySWcEU/I+b0OA/KkT1YZ3Q7tDh7RjZZExIqSxnD0Vlixmm
IViyyX907o2soeGZIG7EsStpzAWWQ7aqabtfTJLpSMmiWkS5sGBmHKHFAGd6FAWbtxWUpINZ345T
lAQiyyVO8EU9vzwBnEbtjNmoCIfoXem2u52+5tq7P5s4dtV984L2eV6DWlw/Usi+/d6dUlvsTXOo
5YTEVwmfz1apFR0W3z8sNx4SY7s9QnZw19OS7PyLfHX5H+Sb/1IBVw8CYoc920p+cevzeLPLM8uM
/tSa+HR3P5TY22TgvcqnT4k+gWxxKFvXbFUBsf+a1KC+1i4rNDI6kNbZe5lOS81c0J4VHNHWKVjZ
rNPNEVmryfmZp5gquvLjCHdxwZ6nX3qYj8+VxFDM0FJ0GxM9SAhU399AsK56In19KO5uMIG9dAzX
TetEMK+FYN2sbpQu478xoXzkk1+JRhb/iBzH4DTDiAq1V8XI5LYomqLyTmAXB0LBPSy7ZkPINB57
ZYIhr+SQy3X8QifltIs8xRc+21KBa+M2Mt1QZgA0zYcFhD9+Ae6ZEHGOF/Riyhu8NcGS5z2yHQoA
VikBYVAWCkp0kmeMt4xWFpZi/mMuHNik+PILAlXTdPbVSmRMLdA5HI3lW4Ppovd/svDL6V5lqezB
ju5/m8Idfra3VF0wRw5oZBTLyp6cOaHrhWXmwNunpoWxFu0Gcv7PhkRKLyQXsVd1eNqTU5KeBisv
SgBu0gljzMaDGW3IpwaIKl4wfHn3d5yrX4iAmChonhGqr9p+bC8hGRb8XqPdbQmX763HQdtiunrs
lNnt3IrZQayIS7egFmyu5Tp1jwlc+pPLhdpKAeFWsweCgI1d6qHzRN/pep5RRPL67/atv0J1LYMP
PiAzm1njOb+OQQDzUi/nt9Nbonv76o7lne42hochdH8QoKcGlfw6uOOKkWWhyxnSEfSlnyLn2KDp
sCbhOtD43hL8eGXOerutv84v3+cUmwDB/t1J3AgOXL8c2PeH3/bM3pYtXWLjkUUaQfXWj2FtP6so
LdZY5m2uizSJqKCKxg2pzRm2kSkaXs7CvFza4GnK6LGtIQTu1uRHBi75pygWtAl7iypMQbhD4cyJ
iGcF7s0SqTC6/WQuaPxsAXfu+LMiJAtdEhpYTpk3NbIjXRD/qI7VtAtCqK5+UqYQ78QQv61LUcVv
MKHX5EKPqSSR/xFmEjwdxtwKCkQncYSFb2XgH70EVG1obX80RaLUXx0LvNiUdU48P7sAqMrPzhWz
vig+3AO1l/rkkIitxySOE2XXtfThFuuPoDDEbq2bI6QFibDydbHnL0mBU3l0dI3si90Jx8w42Ur3
jf09s4F5emVTDy7nw5fBHz3uRiUbIjkZv52QRwH1wzL+Q22OB8XkowwgWKYeQ9XFyCb8ARtdewJG
kAz9hXP/M2zjyGCP3j0v09+O75Vc+7LmvWuB8zTLtegYCicF944suehTnfv3VLBgBRl6X5CEsCTG
zgPg2toWH+W1q6VxtS26ZXsmTQC5zRxiX37Fti/7FdL3MbPiAzBg8pz2WWzLYHBUevBIr8bpwHiA
vH8zvIfpmZT9Yah9m6u1Et4r6ZVHsL2wqdh9vh1+Dwu4fUPK0t64OONCxDA0rxjBGLg1Uku3enT8
rh5kdvnAD9CHmqvi/9zJcPNDnvKk7yzZuX9bWY13Vyl1MTt+Of9kicxUIG+vZ/0n1LCayCg/cImC
+0JTZSsDWcvJBjDg081OgeQGWlkl+kbuvoDHyIjGqIN6FdJejNJIIauM0CejxpavunjLgWDSanuL
OQAPLfDpA0FFM+yi35S8XhM3o/sIvgKDM6tj6lQR9XBQh46sx+xh/e1AW75Tb0lDCuS/GdykKs4m
OJ4JD4c2HGmyS5Zcrzvu2cWInfLFlsSTqfaWL59lXwE6K7NdTe4THBJiU64kBJN5Lus4gOgZ3O2d
rQ825eUWsKLUXdS5dQkPpXsW11ErUFL0BuMNxRfkFPoMhobPQMnYqQQdo7FLmv9mSF9/NxP5WqIN
WCTlDte8aj9jxRNA0tMjaaCH6TrtcjjspQydsprh2velJ08oP7nHxqhon7epESqCFl00FOpjpexZ
nqiLu8E45EW6LhvK4zWmlx2i0mGCbPOt8oGaoTrGaMXphzK8xWXA83FLR4T/FuRfQZ4XfIHtD1sE
htNSpi0Wha0zkWl9tzUPrsn00VWDyNmj0Mfmnho/RD3bUBTIDZZvXGYnu31nFmja2bHtNv85ECry
iREviXLxq+SLWQZRRV6W/AcsP8xQjpDsL6ho8qD68qlF+CNH/gVn/0rn8gprfYgB2EYk9zB3mgH1
+eJPkH07W08vXGorrnkP25RFHkPHRjHcVQrF76jafgPM10hrJHPQzH6y6t41ACz7yEdEiwsW3lr7
lZXuWRnm0GQ0tDw2kKAlmRzC2rG/U1jNZ8fv+htorbnAUTlIDJlxSu1gx7TDktX3XB5pp5fCh6TZ
8PhAfUVKoaqG2iAs9BZJTaA4fBmJDxWcrHgSdCruDK92TtucIu729a3CvgpEhlQfRaKjuH1K6FF5
nl5RXFBjDkhn8xIqPQdG2+fOJGM1KT7RLVsjyx92N9oxLRk6NzVG/xufVpPQiTsd8bVu0rhT80Rt
8cr4AkTm2IQu4oqdfD2SuGLaHQTpc9OzmFg8+rZq9b0HsG486ZCMvsEeooOG2uJvpBRK1l2K3DVd
W3+xuPIvwzfVYSJxwJYYS3G2GBFRUIMpB+EsQDLMSx5wFgXISsbaRx7Q2X1/4ZJBA3cEcXPRCxQK
zKh/u8PkP1bu3gUpYjyqHrx0ajY5o6/EOo1LR9ppCCuBq2UZgZE9N3pga9uBYPQE1Jo73rW0wLyv
MVrkSwS9Q8lde4TItKMfElL5mSCRQ3+Ypz9R4VYliEsQcw7jhe3j1dyKnZ6KBCToSW79LYbKxN+J
N8yJkVw4nBTGSGYGpb37LBaadCo024FPRmTTmdR/YlXE49SPRgkdMQUFzN5IVoRkyYaFGHephhmP
G0pFzu8XIJEnQt5GdTnWXUjkBqNTKxbRyrdqYDlbyG9jPTxMLmzjd6b0V0I7VNghXo2OQFaqJ/Rb
JWSrhU1qocEa2I/psuqzY1rQWgjUeU0t1HLPKT1rGh40jL9NoT4i9uKgU5DX9UCBmByR9cPgd/Iq
07F6dTc8pKQR9w/np8yDCBZCIDg9DKVKOwkMiWcE4v/evcHsH437LkRiAxGHsZZe/UWHXDkKqJcO
Gd6JNURwsYKBBOnA78XuGBqrv+24lCcbenolmDlkc1ngyKm/p8W6pxl+JJq3lV8v0ZX4rutFbKFJ
QemefH5SR9cowLYjHy2PjXx00HFw1OnTsaBX0X7+dB1N+OONx+lkD5GdW4XujtzhkMw2uCUpmF/1
MobvF6x8a5H7VVDsfnDzZtu1tk+G0Qes8TOT4xHBcvEndr1xx6BkNRgKz8pEi5eM8gIq7dnbDRJn
BYxKy1zWloZdK9B2CK3O1/S7aKAdDpJZKYGdxpdkjiHSUUQwXgFhJzty6guIqbkwP8IiF+yKryFj
EQvOjpXZcbDReoVDKz1G2+1GOh3CM9UEwqLuVsyEfGVasPyPLQUuy4H6dJAaLh2WCH52vJScLfk3
Lb/A7syHM5oFQEXLIqOFrTNUCK8nIMpzC/ZyuFKP+/Z81zlpPQ75i/qg4/cCXguoMlkR9AtKymDr
5sKSyVnpvg1QS3HepcoWIDY9mR0g07EpWx5ZpCuWL0QfFaQy6wRloRmIjrgcQNDo5JkTinPMEuuO
WdwlUD/jPuwYkxCMHGnSRQfJiP7QYns/fj5TIUooeIgZ7QjyO9bvOgn/9nStJgPoWuPcYNVGuUjf
l/yMRhtiuFYOGiQ/gE1Yn81BhJPjXei8KIT6jxYmRUlSkzCpdAz3xDGhG2jbhtwlQitkmu0o/7Vr
cmhuIksR1soGdR/4isAkyYzRvhlSuB6X+EU3xhRm24/rD7uvO3C84RL7VdX4d1+69uHCuIwf1l8/
PZgu7OjY/bTGM9kChOJlwtHx743xWAYJGRbco+b2NHYlkZOttAWJAigP8+/aatbP7r8BeKlmoIjG
dtPoFgvrqDK248vBphl3wULta/KGnNeHhptkVAZnLhMCmhv6sA64Mg3q3DuTEq30SqZKPVa+mqSV
dPKSdsu5TsHCHpxav7DCtTVtb4Op7wcyqJEXD6/4AAipCxTuWYBIesw2Y+jDhn+8lBzhBzt4rB/H
D9dWYe1JsPj/d2k9O23VH3Yh7vZvnq7Y3SugC0e5OdN2aiAspFIn8C/GN8NbxmKBbcRG5e7kn+Ff
cRjtEMtgSuZDMfDkbZ/WOZbhAGxGCX4/Z8OQ2SVcogpGgwOpZRT+S/CydT0z6CnDiOLXcb7PP5mo
LKqJyY94UjFapALIvdC2Rcdbg+SsYl2kwyyY6q446Ljc7hRmb+jooMKohuNVSbqD1knh4GU/EFPO
6s22BPt6qw/lvm3Oqxf/jdl2P91pQ8z/zK5+SRMKjAY52rN/DLh3eCzT6zOg4HGFOKkjQ4uon9mz
trqFQzhzWMPvutbdJK+8kC1NaEB0Y9mLcoOinmwJA4DFBJP31PYNQ5BKGcfnoJSvxKqyla11Z6S7
xydFxs3HBJPDFIIK7wb6MVep0uHxZd3D+UdpnOva4/nimneLatBGRt5XuxZXLlELt9+Ew2xvwizB
G9YGjTDUpDUK0yIOvK1VBAPMmPZL3E3jdCjUJfX0Pw7EsDXjc4MwnWx0AxZFCHcycRghAKfEi6BC
6zea9yZhY2KDpYzq4C1V0utFjNqa5lemBJGe0us41M2sMuUDBhHTuTIjqWqthLCq/TIChcl1uM23
i6ZTbLwtESdKKReAM60UbETbo8O9LBLxFFW/azYEhoYuKX0gTpyDfY1qqhsXA/jQUwT1BYum/4st
yuJL4aMgr9xFnnIJT9CcpOlpDpx4Jbiy6srIf+S9ET2LW2ywg3+BAGoXhUdHS6eTkDWRjZvrToyY
KhUnWt98roYmLejox/k/XlBa0KXy0PHM3gM6GKH9wtG3DF+NCUobz5Wqm/CKZp9//d1os27+qanx
jc6DdBZcsv4j6Wrbsq9MxVcmFiNmL7nwNBDI6ttW6dxkhhKlbeZ/ZSjsN0H2dv+ukcMD7dE0ddct
Mq1QmMWsjgvT4hvKbG0Goap39ZHLSY/DgoSIDvFWP3PoMGJjMGscHPkikjeZx4qo+1b009H+uXIS
UUxiOdJUk7idn2kV/vBLz74XXXOM7GlBXxq7W1Z4UTMmy5OS/rUb+4QgtZcO+Ae0rsU/xXDC402J
kYye+4bsI8ZYKQDSuRwB7g72NZPRA3QY58ivRaiSh90kFSYXwEhTg/0bVQdhFumG0vzH1JYk8PQN
hSn86WBMsNKpNzpog4HtKPnjEpziGhjRBTCr9ZVnAQ8ThdNyFcanosdV8ZRyY82SOdPMyDFz7dMv
+OFaPp/vsSuKWhmCycNzir0ZKrtpT1c2K7DWqJJxbCzmcxvNXdlaZlSiBSg+osdSTrNVethUUXUg
smVeyOoMMvIpyF6c8NwmfLvGyZVUveOfQofIHFKuEIwylI6eBHlkT7XBVvS+Mz0vCNDkd9ES9H8j
Fy/H8xzqpFnbIoDqOcVKE6708YlhnXrgtM7Pm1JuD9a6jrqX+0DVrEQEc3H8AbCoxozVaUKWr4lt
OpEy5P71VyMyZKROvIz8CqPG1jI73NqIDIqIY4RKQ4o8lIzMZUPg/4Gs3We5YHrnL3PfJJGoSHg5
YxGUB8/yXGTxFmLlyZLcUavIkDtgaZHlzlEZ5QSIgdzofPqvC71jH22/Rqq6A69hFwwwOsQHIn2L
TepTtqRpDNTV6RuNGu94sreZRxuaLOzQIO19x+4KXoUr4vJpZ3A9QgqaAhpVI+YY8RM6n30Z7tz3
DaLfOL8VFpWss6Gei4XrEO8+ZW5qBtBPrpEevUVKpuhv/xWB7B5JbGCWKEP7REjwkgsix6d/03IH
ty2yXzBD6KgbcFeRq8Vc8u/YjZWxj1SvSb4LXBFvIrWXNvgR4V7ranTW3PMXeT5QBWqrTcLS6HZE
MxX6l/u4tSPngZtzXM1pmKiDDS8hqJOKgDlVhNcHG3+W73EMthrRvDpgzhBoceqK2O0qOMUJH+kX
OOahrSCG4aKdQTI1cyMXFT+LMJXsWGUmhARMQx9KJyvm9jmU5SDbzV7dbQT3kAbof7oDQ/KDnBJl
jN4EKax4Y46PL/WxhbyQn9rMw2jDfELGAOgmOTXMdCqV5lFSRgrMkK4SNqfQaGWWJZChibY7XqV3
tUQXB79IE1RyktIVbT1uNIgn1Nw19yTvxz9HMfq61+HjrTVSLpiZmlob5Nt4nthh7SFKqLNmRUJv
r8NkRtVIcVaR5mqrZCW50Itc9tgEbbbEO98F4viteDmRNa50l+DQ+/hr5nASepros7j8rv+LnlFs
Ocirl9oS+AGjXHHqKQ4QTlzKFTlxFDoHmpJlnBCF+Pm6gumI3cP4N/KYRw9EXFGBhDItnsLfLaXj
a479GzQokRUVfMFHFTlx2+3fEWd7tOi1szOfyIoTaDXWs4EtUHZursnEiGgdPoBZZsnpq4oXpSmL
mNwzZ03nB4EojlJn1UAP+n+9XFdfXiDm0tPPpBBUYIeEVpatg50wkr8gpeKZEP9UoOwf2PiPy2W+
K4lm34WfEaSbFjTtWcg6KYTL3q+t2iELBlHWlb3EQXn9cXkvjKXDJkE1GRt97ziePmF0VX1L4d5p
21zM7SWh2oUaOCq/siR6yR9WUqjPM9ldFio02o2fZgfXhA6/Cb5Yc3TrFfRREAXZsB7qBrxVxEst
MHior7uX3b/M4SNTY7J7vqIaznx9AUOuXWoiD3IXRcZIMO3THzEEqIEaeeaFsDNOi/Ui8J1WMSiy
SFFq6MQRfSDotLPkIbxWhV61d7aEgGHBiC7OMb07CePu27Dx74zWiU58yj0zaov1MTMpK/lLcUgh
BZq6P+GZeGYNlRGXFfE230fRtKtgRt5S3iXzS6Wrn08iF2BPtBTY8csp01CfwoT9cbpW0uty02Nk
qgCQ7GdlyxGjtOSIC3Qo0P5FXO2ghmXhJvQVgpryWn6vBQiyt4EzXXxZjhgz90VTIfzLgxwCpMx1
gH60W4FW92KkbhhCgsFc5Sit7A7I7/ofwGvAA2zpZXv4YjSySYtkziPXQfxcTicFu9QoAuQ5e3Uu
mY3db+tUaXqbzn2aBbJMmRp0wivAHci7JblWaa7nIIROan89CoZH2bORhmI/wggKl9lap4nT5WZu
0htPrlT2ngjoEuVPlpmEBVPzqbk6YYoB9ste4IdRp0ZxTxEuzKudKe2FqE+5raTXI91JcZmbzeRl
FxnLm7pd79uJ64OZ4P7pOIM/o7WkNLtPtth7VoYs/GS8/peYDYFGJYh7e9CR8lm62y2Hs21eOL/Z
l/nEhks27Ibr18/oO76JM+dUiJ4TFpWu3PO96dKuW4E79ory56XIknf77Z+WvzHbWku2PnpOXjoU
zypjlfAxIi6c9uyRJT9YPisXDSO8bOMLJoDYl+LFwQNPllHHvNAqHtHVgbE2sNSg7FaG+AiFaL1H
QtHCwepd0khaCk5c9WVTwGtZUZSZB3fDAhWHg1D5lLh0kFM+eugebXL2G/ixVIH4qoJTpCnqoozD
TynDDiwL0HvP5nqJ10cFD5EGLGMvf7comkrgtkpzYe+Bxi2lzmq0oSXzqo0S6K6yJkQ2lLawKxGn
YA94Ouq044gDmJ8HIpQBMvz7Aqwa8a552yN25ZFJSiByjHBTWkaLK1vZT6JxTf7EbZUlMuQoUG5V
DRPGlrWiXzU71JmS/oOdWMHrn+AQWuQ8qqKVWFlhplllE6mNIRhxXoBeYogkZvbl1ByZy9gnDjOm
UJXP0VV0YDRY4qCewxdpsuusqK4VLCMWNJuWiMlLxeS7lmfAmADO0N6skHj/EO0ANYpznylha/YJ
A1Ar1US/XJM9UKhbmCBX9TdXkTnJXH2nYKXmZQqP5OtOqL5QYOdxFJb/je+mhdyDPsxxN2IhfKxj
nMe0yLhlvz3I+B1b4ysi03A8oXsApC+UX8g5SRVADS0j1XYGaJmjWaU/+OozqEkn1OYqmt9l6KfL
EOrSKliyjkNer2b3NmRaNTi7w2utdSK4rLS8OZAuowpM+Wh2G4ZW5cOklDwUiJDcjGbe9F29O4Pu
7TN/fYe4zauHIokrPx3Jx7cOLcUIy8R9U0rsFPRWtmOvtpMxAf/g9h8MShjKlVcKx5CIYm4D/6n4
gQOSmqz/lr7ZudA3LxEkavkEeY559FGplHOPc7LdQ3bcj1yzE0DfrAznvueCbyUxxxj0P4bT6mrC
cvCHxpzJXC0nLR2vaZA39IHxszvwTyrryMv7Haxnw8uX8F8y1Dw0Au24J8UK+vMIU2w5stjJciQn
Y+A6IhljrpRg/6wAhr8PWLB2hq3CMPWTF3l3qP3cmGnpjT2OY3FYSKH2KqZ3RmxBcCNo3oKwhUdy
L4DIXtFjUOosdMt3EZJKqSk8Lig8CZBSyQWMhBNmjbn5b6HV5fRtDxcGvwKeNBVzurRT/EdYNqEL
v4Br5aF8YdTzmga+fftRvG8mYsttjCbG0n/cRAmcvkyhAGYcvN+WcQjWcPGVPfgczp5MsjZsIXCI
JyDmH47/bz10/LqEBEJhF/4W8muZBhaSBS8EodNCQGBVC7POUoITE3V2XQHAaGUd2oR9FCoH8H+R
/CZYs5A/yCR+D/HDSpeslCtnTWQVuIA8U2WZEVG6PuY9gMHcpNcdy4hkOFa0ulBILvrWfeFcGWF9
i9p0QGM7VDVaAAeFc5kLrnzqAQ28a/4EdB6IGCtvmoAsHhiFUW70/P00oM/MAVhEPrfJwGaBTmnV
FZPVm/guqXbGGp6+FUhqAQm92ho3YqA+1VjWm67Yy+46dPf3YyuDZgQ0ruYTUqnt6PtUrzkYvfRl
Ov+SdqkokwDmbDSDIoE6Q8tGJ/YlDIjWXSTG8iujpSIA71dIFpONNs82GPwuVYo0d64xevOVSc+7
GLrDBg+0ZQSmXPv/7ef31jsFzZEf/ZI2Ogi6wtaNbUizHuLu1OgQyKtz6i27f8CZAbCN2jJ8uyj6
S/kxRkeym2oXsR+rWF1Yn4yE3RQ4dOb2LZYa0uv/R+Gd82zjfofvkaq7P+qozefksdDACfYaGfg3
vgI1mttFRET0fYmK9LToCZZodiTtZqpGdhDGEsJg7e0YqdGNV8l9R4BNeOqeb7qiRQ9Tx5o0ZYsP
+N8Xn0YxE+YMNsg3qHdY3b2eauicIQJ3JAf2DTJHcfwRInvhugMK+bMItA9T22QyLJjN8Vbj0mbk
N8fMRXU9UviLoMYLxz2k3+S4kLPZtRPfBD9kYyXBVt9/PkKiGbiVRAczyJ8DhasvO1BwnduCoIKt
rcozuL18oZ8yK31ZPHDGX381CVKi0sNL/0dBdQ8NjKaXUFn0GuqTUIgI5xTgceT3Rih5tdrqnlXz
pWV62blCwmSBHthgrIzZAxsmO+9FeJTPQ+I66ra3mL7SLv6ayX/EQIyP+I6BGVkoXkzpT4unnx12
QGIrgoxvLChtgdYBWPM3y170wicD54wdT9JuLR3H/w+bATnX0g2ogZgZCQabXeU6Zlkr/Glgxd1n
z5fD5bz26/youzEE4RoHMskO9RDf4LnDBUvXW+sZeA55/MgAHD2wRzwU2647zebPPeJ5oGNkoaya
Xq/p0mmix7GI+dR1gDJsnutJnFSOyfWiYG/DIhGXfN/Rd/5WwF4zL6TCLuozdTXlz1XXVED4VeyN
rPnSzDnj/4w+Jd1GuVZ5hMmQ2zmINd9E7Jgty2+ZXhZMq/fKziC0fJVvf6U44bA2qgAoX5hBrVA6
AR1LoVqkO32cai20eRAh9V9DS1qasNsQTbg9WFn+ZKZDuLiCb7t/SbPTVICHGW2hdx4yqXG4RbgB
y5eMNeVxrRt6AlqH3ZUtQ9N1pc/Mr58O48F8N9pwe4r7ppg5V9/IEc25U2oAfrRrXA+FIL5fnsor
G3HDz9jmFnrIHXiNvfXMcHOW/bjKSIpStSLt9FGnuOV6yx8TPKNNmNL8WNcqiQFK+0LHVZQR9LYx
PjdXKdM9tTqnn/jSRlOviA93iepUS4yu5PSizKuZQOyhycmLYVJOO65i+e4fpTzsumbSPaL/DZWs
qNvTsIZo6D07BuRCTQIvZuhOBnZ6TB7l7Onk0mw4frG0YJXj8+nYLc7fyE4S+wZdf8P7bBjSWFQk
gm0TN/uB+N3eVv/jiAo6jSApSmy91PZG8LaF2ZbRqGjCAaK7oOKsY6xusNyxTHoTx9ybHOy23V3W
ptat2HGHoZnVeMQ2at6Kssc8afoiuM/fIG2163qJhovVvwZ2e5Rn9z2HDBHTrdm34M8heiJHhp55
YCuQL8oAmQN2u73pt+1cGwOuMZucw5hICjGHDtMypaB5IhfICAFUtAxojC9QwffAUok1CklMNR7d
iPHcB3XfoiNnwdyW770PKZxh+KPrTNC/bDa6DQbX/emcyG+lapz6jMtYME1uw5e7brw5k3me55Zv
9QacLgDIf0eiRV45O2u6bhGQwORc1kGw9D1J6hLt5zYkTzvuzaGi807HqabyT0YNQw6SoEyhLgDY
VdcMxnJ3LBm27r/TvfcisAaFZCk20Di1NmIk8scKpERhOFInK21ZED1dPwXbLxhd1bEfKJmCMoVk
GtdmdS5kSrcy2kMV6gxH82b3DeiRpR/cX8asrlly1MvKWhp6ZxLBYf7jcwtX/OdVSZ3KSAQ2kOa9
zL+KgptYwkW5C+r8b8olhwLXZH5T+4UPXr8FOn34bitzLBC2nQRq+8RoTW3FmU8TbWk4tRn9LsQ/
7E/K2R7zieAnbome2Nesld41Zolch4PS4iWAhlKrb7UQJV42ndz5Fz4nOe9QDbR0otJ7c40GIF/3
XOoFjptsYgs4/0Tsa+v+C5JjSYS4KWyoUdfD7SPBYEathoAixuQpsfjzqD5osJpNXlybnik3CJWN
uYvuU3sJFwKWBj7hfbTwfnrRE0T+8c0E+wVn3kfDZHpDm+ukAFQA8j/ArIqkwiYh47b7D1dccv4/
pBvuRC3eeQntQS60yenomh55nx3jwHtN9F5QA7PabMkDwFaZWaKyi3Q8yiv9Ur220aENXjCLsuuF
QybhO5RkldHedSdzOu+M5LBtiNC8FqSsi9DqiWkejIe5QZ5BJDaoQPfznZpV0EUkjZRBbTF2VFft
AACREKmjNMoUQfbc9qp7BmyF1GhjhmaNFHrs28F5qWhylg80Q5gp8O0OA5pkrPFWhkYqMqCGmRlO
yRxedZgtJDbQHBtbrKjdRcOk+9wBRf8Tuq05Z580ghNYKsjRQCbOEsGWIWAtCEPYfn3f4qL9H8/Q
uG/VzesKiagA6wRqUaYviZjuJyPMiUXSFFKHZBRc43/rvdjpYLXM/BXLzoMwknvDNIy8ULjnLyE7
FzYRIXzvlA+bSPEyg+Cgyx0Dqm2KEUbvShkKq3uuEhi5rOrzl3GTlExQGMtP1c/ez2PTkY3kslk3
hweSaqw2NRIaGV38eL5itdaUE5gHWGn+SO0+XrERsmsqgTcq0FAENvx16fhEOMn3vU3NKCIFLvFR
swdcP50xwxJqLhd+bQpv4nuvjF6kIULD5uIIXx/noYhvQ+LV7rQjk/Ahmb+4jP8osu8F7w8+K+dG
C0KoMBZp7/dCHYqVNIe6upUj/H4jhLtmDg9Ke+hsa77T5AFXEiEpqwU59ASDUg1Rj2lc0cUDGYYR
tyCmQOYtPk71k6ZXmPiXqV7jmCcZ2EOtaN6oGKh8zztqRgZ+mwon9M4zpO2ZwtZ2XsYxcH+z4v0T
+KW+K+jzzaDByEfwnmvzgx+MTpuo+94yK7F0o8IIkPkfpHthUGcbKlGlgIS6xEj7NZN3UTkEKSbh
oxugem6uTVtj9DKKAox9YeMVq7356DB5a+BG9/SXES+2oJDuK2WMCWacXA9+u6mzNLv1Zy3sRz41
PK9FbjikirOhyD5J2VLRjsPn4pDT3MVmG/erwl+K9+JeKcgcJVEtMMSjcC++o4FPsE9Z6YDJKTvT
8V9uXy8A375gcmsc+IX92XXzb4ZJMsgpEtHYF0qJjfONNYKVSQGwbJaoxxPUJPEZBIMa0rYOoE3d
zGqL7xRfaa1uucQIzKi45IJf+/ENkeB2wUoIiGpv0VpxTDPeZDqsZFFYaZzPLHvM7hggAqM/B4xJ
4pF73gi1Bkjv9z2Pr5BMEIPdbP+u1Fi2JaWdhkqoMvPHankrJQrLXOjQfxRjkz+sWb6wEv+Ok3pd
qu4LP19KYE52/IEV0cqBVEARl2xpjNOBJrtGzf24psa4AJRufEUj8GTYBwYIHJho2nxdOQ7rigCq
QTURc5CdQRJqeZQtOKJO9TjG07nTIDLHgLJfUaioCCEIiiKapYtT9e3wJbbqXHsdiUPiklNhgFO3
Yl6tX9IZyiQThWCxOuZTGdPtPe3Fj8z9idfQu5qnlByqgW+nKIz58vDTNmOQWZiGtD95RU1AIGo5
K8vVs34mnFU49imhh0q2v8za8rwjERQwsWb4j3hJx2ONGKmX4dAN60lJmc3rqQl15de8VvDS6DaW
B+/ZVISSZjH9eipP7/w11RTo5cd7bM4KdUbq2plter+rttug/gdWYQqupT7U9Jx0OTI0lHHYskhf
izW9bcD8K3QoXP2IwQMq+uTaS9UrA1MG2ydMGl3V9I9LzjrqnJCuT1E2F/0N6uEZ32zrEomO7j9C
sT5VvYGpyG31hRgfmQQ6HLczndOBRQjDZHB28rrIn4EJhczBH+KBo+pfpTIFw7upjXsnKxmTp/3g
PUYvKw3s/OJGTbWHsItCKaQpe3L3DFbcVSYUQKgiOviZwLfolBo4z2ZkSRxh+HCcTXW06SqjhkVs
BQ2DIUGfNwee+gNpXeTtp+5QUIr2DP2XtFysroRrIq2cUA89xbvQS24nJdceZly+WhqDNKIwwixg
yk+OMBYlaT8SccyzPIoEUxVgEoukhHRwFFFKk4kXSbGN0ZZ/7HCTvF/WX5Py5pE2nofySf99LR2q
06F1kaktDEZXIs4vo/xCvhBD4ccpt4cYwtjsJSstmVsJWOZKaBOqq1OK+GpNS4AnwlDHykOXZH44
yD4TngvjVtVpkpd7TK0t40nmxtE0qDR37wp4t131steY430iVvoArklc5P0JqDYq1UIDAmdoUJy6
aQkTVMsgDl34PY+2BBdQ+2pDD76vxIzh9clv/doavQWKvS+D8Ihm6YPmF9N8tc/tdf8eooBPqiqP
ubG3bsToCGwmvAhiZkO7oUp/zK52/qj2q45aAG7UMzOs23hdpac8YVdOpoItfdU/ij7pSBuwCAfN
asv++Ea8rvrSg+fTbMIYTeub94yIiP6Y6CplNTXCVxUNvjdi987oe1AWvSOGbODueXHrbPNcecD5
uPHSVSh0floCTDp2DlYrz81iB+f/dmPVpWHjGEzhhzeOO072MON4WKqrJZbm3Ac8D89vmoeoRnor
/kyfmsXzwZCJDkNH/L98w76v0MwbLWMcZTLilIbH3BMSxxFg2L2pd3oxcIAvUV0shsUuRi10UbW/
WASbydSwS0gKH2+iUovav9TM2FaSYtSkuLaXTsHxC8FcpQvSZSr64D7gFE3tN/8myrfz0NfonSow
BRXzhrBSzYcTVV+9dZBmXZkyxWtdi02j1UPTZ/ljKxT9lLI0SULO7Go2q8WZz2rhwIS9wbvhx08F
JvC8hHvb57pdwkuSKSFZPp3Q7SBKtBbqLwvf1bszvJ7cwwJ4wS0umPIOIqKbWyffg4q2Xq5KsrNT
eHv+aBmIoHVJin+VodWD4cY/zl2bt4V3YHF7DmFPuhJeDDhmGB0MNAOU+WuI4YpUJ5Z7S4hBDdBR
aruxSoWp3POFE3LKYSXpjG95wKx3aHIXgethc6DhaO4L6fhAYyKk2enhtLMvrzuraG+5bU3pNjm4
mPWRqTGDzLMhZ2k0Y5JV4ik0iDvoMXUkAIiq28vSAln+KXPGpjnOrjhMnhtG1Kyz/fAW3FmmCB3K
bZQObuE1Rc7HSWDGBww7xRYl2ik7X6wDPU3wplqrusJHJIc8+eKdXGOtpEKBQ5cqX3qHbM9VacWL
7VFHGfuSWuDsPxhVLdznc/RsZcFxP6LVMvc4IpYkpssv18fuDJptOIMqn4yQ/n04uQBRMIWjjb9s
07QU0ZJAMWQ34gxHE+u9J+q8G2VCDAJHe2jcxuoaIivbBb6NtOPTmMUHkdexAtl4C4kK6cW5TDvJ
SKVDZ/+IQo6zg/4npHgqDNt83lhCjbd3J8lyE03WhdIqLhuTzXhdjk2USANFpwtMl2B0HNe42G4j
47fdISnRy/c+jBlIpG2MIGIwT1AhzelEI8lLQ4b4AaF/07fMEnvgoDDpd3Vin9PqB0J4MaTmxsr6
9uXoQSSVQ2O4x//PD6pt1ggpfIGhXaMsost59zJZ2GR2MRGfdCRe1zIu/3WBVqNezs9hYiAoCIKx
8DWXd7QF9HDiD8R8UFuHt1puONA3TPOC4qWMtFyXzm8PoPXSkLNu+B4SLjrbjwLhzoa7Juu67aYR
pq0gx1zF6yRR0BGwsMF+hF1zW9IV4oxo8XtcNeDG/3K8PwZBAH1xo2gmTHiYxM2sEnkI0ggfZHVf
8eAz105IzhYUSSMq8Gse2FCyKLWeT5gUhcEyBAM89LseQSuEXChU78ZGEgLo5x7IA3ypuOwgg5e0
kj0RTLHz5MW1Aw3IsnDyXmMmHJyC5mBQQKkOEQPI7n79rJZHnHKXnijn6ypMV9eAHieWn0RUdr7c
ubFXBqdFeyYIpQgbVH9GDt2Xph5mN4OjTh5wnwTjP6I0dDTPyYsBPzqMelS2zZeXEU5ecb2a/vCB
CviFaTTrKsj7f3MqafjAX79IE9fyUdgPBSl73fnHZcCb5eUuQhhw1Tz3ITppc2robLb7Css/0Lvf
9Hp67UBVt7om2GvAC8YjFyQ5uBOl4BqOFpiQz9JSB2QF6sRHyBFi0zDv1p/ziEI1YEw9tUv8cjJ5
3+OUE+ESjz7RbYndqNe5Jz6ogLJ/x3xpLcpjqNAyyKNZIM7gNLr22iQkY9Xhy5PDy6r7l0xhinUn
sgwlLaldNVI61l4+d/sUUOYOTMkPrOrgfPMrrAlTKAyckejmzzyIwFoPIA+SEYMC8y91meMjO8ZA
b8E9S1guT5ZLknFHBrZAEOqZ8Tjx7HWoIrkaJjo7IJrTWIcM7hNiypuGDWw239aw0AszPEukDtbs
t9YZC6adZcmZ0x772CegK3hXB+WvZOVy9qAiGcLsgu2UYiprY8UCcGJ+dKHQci1SfR+XJs+2GP34
Es9u8ZZedOQgMH8WpU+8eXjWdGwT0yEFMiB39/7urkJQ6uC5CvVY8i1SYHP27wyY5Y7OxB1Ti/Vn
VbcBbWoKz+tjuoTkCY0uP/1Szk6nqxnH6QzIgT6+HH4AIGhnyLTl/Qt70E0E8VtEhf5yaBxhtp7Z
7dJinLtR827PJLsj2P+oZ9+jSZIulz5Nl65RPvNXjNLayOnkWzCbN8ebFaI5CyW9iOKHBD/qzfQc
WZ39tvl8TLyOK+DAbvU21h/ibiBtgVFyn9e/oRanvdTI/ofjB0SkgL1FigZ9/soPhy0ldIMDWCw3
coOj0unNbJHcuBuQ5xEpHDgVkuoYKgCnZZ12MCWmK/qB4GtRQx93Mp7CbtuaT889Y0a44slxuDT0
GUf1mg7V+2869nNjahVDvTtgVIbV6C12zKA6f2bVj+ZQy07UC+BPkwMS/H7Djw7Tv7mPPfXUlXuL
zHbfjOw6Bk5A8aClPDY6Th2Seg/uMk8Hl0lj/ParqoGAk5j8r/nCOZgO40SiRsOm/PS7NAAlNaHe
dljweeGuCx7dCjjqsfBksjAgpp/FH70B2Pxe0U5Yf/8GQ0TFFklr6sKq73fZTUq5quEGIfkJl7DO
3GU0iHfNrY/Mz/l2kN1LPp411M6XNzgggGUFZO7NVijO6Dv0VcG3lDrgkP9ITTK7BfYutVSBHA6M
7EgieSNWWMIsFZwTOYm/9TdK+zXDQM4XVtR2QriKHlClPmeEXQqeG3vpxD2DO1cxMYI77QuQs5Uk
9jb9x2v18+SoY/TPThP/XSM3m56Gtteum20DHHjhK+7IupC1OOpw/Q39FWanGCjnbQWuvRMm7bls
KSBIAfvxVa8dACFPqwL/lwDzoEJuYzxFSformRcQmrIc70fu6JOAzP2xXhvLUPgWl+U8Fv8/d7Gy
ePqeeCAsr6Nfjwo6zDyndvT7jXoXnpiY0DMM/otCwPgs/dLZAFS2uBFB51MoPucccfi31uXQkIW/
eluVbKqrtP58pFQiMVVpuRqLxj8kD1gGhmGhsAq2CKcv//e2o8BCbNDkFHXUP4ykyFt3TzIsrx9l
9pEXKJIaDgoazrCpFNYGO+cXF9nqWx/YosI7PMHPUFv1bD6v4R0T0Bs+RBRvZnUS4h2jX+a0kuRM
09mVgXmsOiCBHcO1Om9HUOTIWWZbfxWZAduu32N+k9hMqSLcZkmg/M6J/tjeN2CoRu2vWFMiOCn8
w8t0+3/kpMqmfNxzQvbqSUVz7st/Mo3ntUgJgh/Kz7/iTE3JJixmsJjqg9bme6sQNoTtyLuJ1tAD
mta03H+LvVjP3g5T6Ey8D2fZuRAr2iBcvVAnruPNUlPY3a8HaKOQ4qgTq/q4/Oc2Ye6gxqDnuiR3
hJGM/Jp/0Wv/A5FxdMQm9SM67tVsvrYuHyqucNJnLoHvzdx7ylJmRk6Odo+HhXS5NmRJvcZCBWwg
5nXwqXJWChMH60g/CYqcr9/zsWYCTInJLaB0hvoJHJ5i9XjtlHjNNsCab4hKEnag9jgKz4faJ7kw
a74dhbnoWh4Jh+w3BEPsnVyfA/P81YUk3BpwL1mcVRmDGhVnN7co+X4I+IEsFtbJta+4ocIXY+sp
ngBl8T9qiydmL1FE6eEp4Rbo9TFtQcklbP9rGDv/UeLg2YDNMfNKXOoG432dLBLkxSGbfI28PDj+
FUMVXa4NmNsOoCllS0nujBpk0uuSaqyqZqHKdc8u8lcsLt0U62q+3Hh0IiSETeARLTiSD9BnDdWR
OOKUX2G5mUvQXeF8h1mnPoyTRrUmQxVu9BXB8uwrrfJDYOZ6ohVWkY3oVTDU4MOrXmgpx6uX+ESP
27fWzG7CE18tUlYJ12AgQC4mwDo6m+IwGJjXqXKCy1iPJrt2/LZAFg9Zz3UJXdvX6kbHsCoBidsK
40LkX5fNeMk2lr/si+oDH6sfgeWmsMcAJjWblkAbFFcgATdAO9z7MS7OGzor98I6SN+3XlVkE087
2XEeDKDUvkWCqy5iW26iim4Ve6Th1mOprtGfz5icGBnF1D2Y+LSEsnqZGHG4VA7wO4b5l8TORXlY
qyEARHUhI4gwhR/S07/gmJ8kBkhdG1Tq4ntgXgO0atlUtrb8TMMZZr78kLxtPz12+im1QIBsEpHN
kVOXZbAloWgtm8DN/B80caKTEAU2SMblw++XspeXJ6OyxQtuS5DE+189aFwQ+uT3juMuKYGnZYgy
fZa+wMSFj6H20/v4dD2X8SoJwJc8kW3k7VXa+eqYAhmqbxvwDY5iuYq7mjuOlB0l0Xgiq1gcvqgP
M9d4Kkvr1aI3x7luuc82Y5Ox07E/ZUcD5rEv9eO2zgH0YrZGXrqlSHkN+KyuWWoaIIUlXFWzP22v
jCtOOeaToE8mzFiA4e76pNONj92+CJH6l/L6hcrcYH35DB5FkXyYpRodO8aTFBfqf9UZZ98vta7W
geYgGHk1+Cugu9l/Wg2JeuiN4C9EThXj4o+CaX45TJ8MSvbiCU3TcaP9pd36gHvTUbtksvQOe+Za
V6FBQ4jNgnFb6l+9mhF50gjiBIVYIq60XQ3EixGB8Rn7bXAIueGFChRS94U0z72eJPE3tyXnQdXV
TskXrAVEqehI8NVjpGlRs1uklIPLJMB/xNju94QpVmWwKZN9J6I+s/TKhatbyoP+dyz9xZORVXZ6
kqfzlb6npXOiU9404tX9YOjR6MoElQy0gUV04xsUT0qASKWXVc7nRPANUbka+cDFCT9o+hWlb92e
aGoamlnYOgGu8Ki5+7R6hJyGWHGtIbTCe8LeMKzYhzEpsGALkGb7Y/uo88QIDXO0zWKGO3CEuS+i
HI+xrSOYt3Y4v6kMYxyY7TY2/8W1mBD31hGY70NhMOz1gQ8paNqZahO5U8vYKxRp6bZ6rR1y+oQX
+tRP3YJstFiyHkl1JGHNm7IxQ4FkoOhdflP3Wumu5jccJGOTzjH/tlekNe0kOvj2Htv/CaCG8qTF
kR5xBWYwxHsPHbK9WQN91WKS+bw5vzZcjbhvM7vNhpU0cqsQCRa/GBNaap0B8I31PXJFY7+KVm3d
7R7Nvv11qr2zpSUmMvFVCpQw6QueVobnm11XxqcVoQhx704e3E/hAMPxyrN4UoVHZRzIL6n0CcX0
JjsnYplZtags0oHctg9GceCy9Nzjrfxyx097hB0hK+ep2F2XgbnNSGMQA057+yTGY7v84MtqgLBs
C+VDWnhlFGS94Q1SlGaXnVsgMRKNK3RY1Zz+UzSYPlbrWcgGhurvaM6H1zL/m2mbPEJG18Om72C3
WGKAmxpw1chO23147Z4HUocuRvRJBKwRB8fuURh0t85VFOLkLIIEpLI+QvR2YnzWKv0QdnpTcgvi
mZ8YfbZET6E17yvaIef6Qe5yHl1vuxbRKYrT/uGxFhIjGkoESEKLaix4SEm82/uJA9mWhqpeSZEn
3cu6EdCzYsuq/XADrOka5sgjqM90GpbEPtBfzuEBxQHLemnYETWm+15JubGY6zk8dsU2PtU43jv3
DqNoX/ocEKP+KL9+gJoZ9rAWkGJ+TVzSJKnC6jcBdkZOh/9WdOFC0mE4ryMZgnJAXpdPFffMkyfQ
jKpNSOOexYiydEccIoI7mj5FLrO84SYNny2Z3CqLw8gC+I3IkRJDys8gVNc9k5XExW8s0iZnYIpm
hdtNiqPCE9Dg1yRrmZSs4CPpGzRp+Ng/DY25O70IooTWAIakfUBmwEgHTLRdmXeecb6nSQ2DT3g2
/v+2i3bWCQfzHZMtDyxHwXKhP9cCzSjDhWP+ZnsN3hFUIaB5J2k/bgpMKBLtpKCtjb9Lb6D9aUyF
wkuK2P05gzdS/93N84vZnAQUO301UC9VteE8A5rAoaKt2wHUW0qF/vxW6aZwLxMvBWmFusOL3scs
G2hZ76Ez3Qn04BRu5eOmRxikMRlukJW8IO/rSI7cKcHSYxusV9XbXEfnYMpUsOzJslqMFEr+lhtv
0A5iCDfLwOdLY83gkgeGCz1BVVQTcPWMkHQB8Atmebv2oxYmh8rLTY/IzPHEDSJ7BSQhm2jJD2N1
ReWk2Mp/KbXya1aM9fbDj7Wnuig91YRfA8vVN5oSZ9gT4SrVYIniJ4dWNrdZUS58oRr7xu2flS4X
JPKW/c41gYVYFg+weoE73nQwUXVr01nSxhjIRBi2owSdnE8VH/1fb61+YycmrjIKuWCe5muMhf5U
PODtmDI0NTyUBu1tEU9lk9rp9c9Sc5SshvaArQraHZ4COfa7J5eGjiJE0MxEKI80XQHdEX1nSFTQ
hpMCmMnrgElDavVUVQMYU1mU7ThcW04GQP9BtxnhIhcdLUvpZEfXdz6JE7TgVyxs1Znb/w8rRHLf
YKYSLnzxEqrdSFqd42egSy6z4Tp2T14zLZZaKmPXTOf2LLhEyGk6gsYejZUGRl7NMNQJUCmz4r1A
M/KMqqsP9QeggiS8rL98JUsy72dFHSEebJmJC6bihlR6vJloRWZKgGClqhpEqEEDWcI/UhLsi9Gt
h7UfbTO9HmuF7wEuMehKjYg8qeLizn4HsO9SrKCQn4mv0MZUD7RhmyRabABOrhoiA0ZFj6+kkaTY
wouLnmedH1hlM5cxo+hXjVwRCe4Si649/14qP5baXaWSIP66bvxWBGx0HjfsWQiAO6IhVsr8QPix
nu7vYZHu/I2PozAxSxgviZ31BOf5NWlGYk9/2MsIiRwzCqVsYnqSmZTpvg2Zvn7rhpqRyvhCGIPT
ZmwVANORR11jdF3/ujEEIHl6SUOVwFojN5hjjEiWJBNyM+rJQMqvgdcvZbKEGUldq5jp6ePIJQ7h
6ZWt+C0mxfGix7whV9/lfWAI2DgQlbyHWlaAE3z8dSXuTlB6ZR4YYErGwNpHVdX0CmGmwpUXLlyf
Q300foZBIYLpbYSH6H0FLql2enfdgwwUvMh5ftGFTLACxwG+eUYazUwMnBQI7tuq/2OcqP49eby0
nRD5l8wzS3CAAbhFdCRUN+WskawYBRDxJuGO6nw2Jz0NSqLyc4oVNb8gsHrLKA6Xh0H98EbwAZyi
7tjv2t1ZYteNDzZPYrAsNru8Sh/hPnVfvD1sqP3aaNeZfnYFbe51TSGEtWeYQAb8mQCTFh5MouQr
DNbJfQqedztJLhXt67eeefD5FduG+KfJqVHHkVALXpF/Cs4ke7j26iOVZD8DF18ikplx9cDS2mf+
KjFwQFtYD2BRQK4LsrzFQR6UrpBlJfmNdezqk+20jXxmwSGMO41wiw+ZUS+dSu2C1hbE9TZyzYQ4
IM8U5aEyqQjzrud+yZeh4xV3SnrsbHu6QiDj+K9f8uAUYICUfk4l3UbmTVg+JIKv22ulZxI81M9T
nkeJSwT4jz10ziTtUfvg09jHZix6MdW7W/rNaHYfA+aKlpk42Nwxunir1ZOFheZIvxVVh5wUYFPS
HSLbdIij5tlY4AV7BSd0ciqi3EqJUwmq5uiLs170KFBbGLJszgQL4fx7RvvUOIWDrUCQjg+i+Ojr
iuzkdkTd1zWfLq8o6FmPqit7+hUcRwHSHoQST6mHSrMRbhx1iBQHwf1jxnQg5fu5XmOBcpa1u+Ys
24CIVd+j4vlx0A3+bj7GT4HgiRMXyPjVAki9ZY45DP0/5Jz55EBBh2/DiUdBdIq/XKT7BS8BouZV
ndR25i9/rH2rsao28IQHgLdDnHSFCtponHxyWkNsiQN9FZVJu2GxyPd1N3rgOMx4YRUSKIqp8kNT
+Sax32jsHLTrEQaJ6QkO2hEMDyQTozBK2yJhMsFCgR52jD9Tg1dSXqbHD060ppwc3sbU+BtnSWln
EO4SsveozGjP9dm/cG4qA6lCkCJMWw4dTYpxgNx5ewkyMJyxkOwuzwv7W/ObQZxR2D4GfIvh3F8E
ihfwadOULhjD55BmL2zYZvu5wQHQYsXr9CcxwKjAVzxz+X2ind6bxD6EqOwd5d9UTRagcvNMNAaG
xi7K9BzS6LiTLrfr5uvsR/lLNykkXgSI90zzPmVTlewj5IEzL+HKShWp4gjyL1NY8F08JJRuA8rn
o5rNet+fd/kFXtk5LXqKCAZUAO8ZqtcqaAw3wcRyaRMQsylXCs5MR7I0Bb9CtHbJ60H0VvpkJ/ze
A8b18VB6RFKY9czArnaDl8M8gqNPhnsPe6fMV1GSyKJmyH5myMVYncakMJBs0rtKM8lkO8qx0idZ
UU+Ih0Ni39WXrxB4FXEVoymd/eRqcx2MHf444Znaaw/Wpp70QYYcpvL/YT8FTyWWEzZdW25dho/8
f5BacakywlQM5J9o3l1ynNM+UWDpqe5lWdQnS4svQu9r4PMujyOfhKvaXsuw8l7CNx79/YkIkhMH
4syMdy+c7voj/0MhBX7UG0Fb4kczZ7hmeZ0SiClFfsoX1GuS+By9zsRzmykJx/xpACqBg8F8gXDU
xnd7W7BVd3ECmc2xIjWLYDN21WrKxu6Bqx2K7hy1KvaROz8BLSKtpmDIYcCZ2hB5xn+gg7I8sq7Z
yvl9aQfYfk+eq3C1qMOw1bp9CB66KL3d4/19ev5VCNvBwON7OjJR8WjfQ/BbbWqfAmYbRneEeaRR
YiQZbt/lQ1m6MQKNYnsG/E3DMYpphjPUtCnQjmWxHVjxgqha6q0p/2WcJzYqWZNb31FB7JUFtdPA
8U93iQzmOEOZr35hYERbRjl/Zjaj+aIR9ZfIoHU3VpHTNXed4r/9liZxokGK3xX04s3ym7S6cb3t
3PLORyCXDcMd+HHw3XyGT6nnQ2KNXJr1PoMQKxX/lAIGfE/0+1eL+rgJs13Ar70Jrl7lIwf4eLW4
o9/xdj7sRc2GbcBcy+R0I9mKRnCCMWKuQLWJLRI7RzcR+mRRJ4+SyyTQrdCd4HmOm5UrWYbVEQUL
qlpIo6rq6MYDkeFKdB9p+hw8b7/pwt9w02TZwJCvyGQYNjkoAb5j2azQZn5pFcN7s1iJ2DyczkIP
8g1jQIJpNkQ6/hV3w+af1TLMFIpCH1WXADyAHZZ3pEzNej8ZmLoKkdpSpZwgGpgIpTmbsgoNJ7O2
PlTy4BjXunuzoBAwwzVQmN7Gf+Oy2dq2jXi3dMAg1QBYIPu4WEjZWKTR8SAHrdXWrowkPdBuMM9Z
JF7W9HCE5RZ1CvPvSWZIjn8nx8uerALFg1cKwRchsQ5P+4VpwZjVFBxVThSGgn1EVePvJU9JZG/R
tLXLLATEU1ACXzOkq2LJSLZ6RcPE/zjeuNcX37KgWJRM7EjlupsrjEvDKUN3Gi8VwvveySrygW+g
bEXLb5L0VOSsMPTt3RG9GlEjH/Yhn/flfYi0QyjJWGSdKjsAm9/IGBE2D1QRmhCQW1FwIjkdn3n7
nkXzVz5Pg9QRaUqgePUNuhELyZ6MJneg7t6eankj1ldYir1r5YN/Q0FY0q3tSnjBMi4hFrOl/jJG
dImHqCYb6k+9/hvhGQWnlXw6e2aK6d/Sn1WiooMCKW3R58tTXrhBU3fNYfcsGPOjMsg6NAIW9hBD
xDxSEcOMDh0ZGrVe2cHA9CSRT/CaiLTas56nPCjC6eT+1QapcsGm4VqtHLiktOKqAJZoeT7bL6QE
FQbZ6/YOuEiCmTgVfhmIiCJtc2VO02Qzfjfx93r92ZSJAuJTSgu6jvTLXMjs5BTVUf+Bh9GqAKuu
Zcs4rO1nX2Lfd1mKGcNwVfgKc09vrm3by/6llQyVuA9K4bEm9YlZ9MtiqXubXjvcmFTaJISXAdnD
6iY/0fyBeETJA4TjrF0WmVa2yW1D56aFPNV7KrDHsarq6+w+af+8XGL/0IXXGvGye38rI3Bl9THs
XI/VaMvu5dNcwDSSwsiPe9/d5JBrb6u3C/xOOoVAmKh7rLRT+46SpI/5nRmairs2oeqnC18MyERo
pEomOkYZaMTsA7ZqRSCkyyh4Mi47lcqq7+nL5PEot49zyLUpniyRb4kVOaqiu+lhGqgVRGtVRf6H
BWKn94/Yj7re+ZtQX+Pra7/F+H5jfaRXT0EnyzinnFLUPJuwKcaPxRb+P17iZcIwIuvshgZIb1Dq
ZpzWdlndiixDvNomv28ki/VFHEPigizisKXPup0/XGxXSuxTNl28YnMkx/BZX38s42EJMBht7YEM
2iBbEto2ElY2lk1IP2f8GS3X+zKB6IYztTABjHzF+EzvovU1IIxEqeW5FHVRErxIMylDSpN8yP83
RKynv43UiCV8y2i6wnl8PG6nsN0a+u2gU2bS03IahNFycnVNUMwmCz5s5tJD8t7opBXt8nDmGca9
hwyKp+th0nJwA8Ry6MjdlcPW1kXnpyvCJg3KP5DR9zGc5P4/LwciWXakCr8ihuS3GUJnDiZIBaLP
y6u0c0oDFFYqKXMv04J8iTsJ9DOxpkielPrD3nIbkfR/1w0G9lYGy0KKMjHFUcrbp+G8Mxpr46v+
dazYWatzW/rZ3Vfu1BJkeJrqP9nJa1NvliP1DBPLcnsOoSdJpYDs/feY0Bb4vxNNaf8VDgHR0mnX
qEb+2PB12ZzlA8V0ztEKG8fxeq21iQwwDsdCaj/OJBSE+QV/4CTLLv0tKK7g3GQxzOOLP5WjTjQP
vzAUW0vkfmK8xy/Sx6hijP2jAko/OfnfciWYcv5q7zz3B9zhpGHblZlUUS6/DOi9tgloaXBS4Q3C
FvATrI8UCL4Os+K8KGnVqM6kXrWFye90rBraIWyjgl7grS0ZWiiBPv3dYCiKe22LqGyzscRhaBF5
kJyKzQ+dh5xaYggKdpDrpFva0rdbsV+9Q9zkxQvpf62froDpFLCXJ7N9E2d4XSiD4wuQ3qmo6mwI
+6Nv8JW4LUFuc2yLmGeGDssqm17783vSNAAScebLCdSX61NA7g6hXDibugEBM1sezwskg6feLwYd
/cin5kNF5dO1he9V6GpQ2npV9a6VMtJzDGjmCT9gL24gsQd291wIsKV4hQq1wAwFNuNrRHkh5rA8
bzpzzBB0JXOHHHEi23RMLnhEDw1A+fcgw3+9WS8JGmawqZcUzCoGdaXdOcAbxZ6KRkyNqnoOQGBo
FWf0JBmdTBI+obi7SJdPCUhfvAHq8ReSkKyuv3C+AhNTegKT/6aZFW8qhxyFf+rBrunaGfXZbyjq
LWuH1HRtHh+BlrgCIB8zsFpZYUkJRi9EOmpqWqxT0zgJOysIjMIYR0c98YLTtRuKLe6kiLmitQCR
lO9SQFu3bOvXKb0dyMM9uhYVUBaRtZZUCl5AqXG4oKzmuMl4CqLIsvoytf2Ii8+KwyOx592nrURL
azmSUTtq8JIudGGNQ8YNQcmvl8bQhfVWl3sEmySpGQiyXE/6LQPFykOkcnvksy0gybBMeLEk/BYL
VbArcG94+7avqVN1F6NRC2r148jggtpmnykpk/kkXY8xITtRcJmuf4MqGBs86nMrUI8fge61Loa/
m9Q4O0LV/JxTmOt8igO+8EF41/UeSHrQloKTSvvwRhLAjp8S9aNcZFceDQqs0U8zFojlnQyyFiYX
Cgf0BJgUs2Znx/CrF8EZWc/DnCqxbLeZqz0YIXkT/bRq8BXpCxQFXkV0nghXJqxun1ZNMncZWQ1q
chtfYf2IJAUsyYZkZPJ2svwJ3rTgEMd+yPjUcX8jiHfIQgrlNsz2a8IR8Ty6KetbD/xlLz93oAqT
cbCLtscEKxgQkgutehWeGYR62Rlaz/4HQ+FdkQpp4SLzOhDtJtyz/RY40KEf2peTnMQrSj8cfvYL
mjybPnekjvXtVpI8X4S+1l96k4uWYCbiMnr7DD8Xs6B3hR46uF6RQNuVecFXCsbih3+zTOf486vr
3fCcagCxl3hSljx2l1eNLX0SV5LT0JQkDa8/luNNauPFA23G4Q30hjZWITHaXvSLy8vHxbFyoJ9Y
FGm3ptM4maFDNuNrYVaP3ZGiPD2NF44oXcMSjeM9z4VecM8WJuH7ajWwPQbGa/Vn3PMbJl8mPJv3
CUyQFdt+cgGze/T2FJKsz6AYaYZ87T102YK0imnmEOM19xfxl/r5CulZvHsIAoU3lhS5681+UY23
PoYkPmaJJ5E2KvEfif4YcQFSN5dImgAGE82XPE7OploWdba8PaG2UOlUnl950vGjX64D9PgYzjzw
U9Ub7wQvpUrmwKzlzhwAyBLvlEG/+fN3qC588aEnzuMBIyOMOYCGdiaBzbRPiTexoTPJBFJASEAT
6j95TBMtU3QigvCiQc0fMxy+tCdTmYoK/dwWO4heOR7ORvF7nqWGzRgp9goWynqyCWlGAqaNDRxg
Lfh0rX114qw/LTZulSlORVQXNjSv4N7BzvUK1G9PyYyIBRTRnX/lCO27DAMofeE6WT7vDPCQWpmD
w2ZvrVFLMl/01dtcv3919p5dvGE6c0nqAUpSPwLce+CrwSYwGa12lUzvPMITYd7zcfNu9OC8ZJQq
lmWqBwPnOHLXYshN6QrxCWKWfIv1cHRsEd9mO5hxhNOVxzTyc5CjTIwTF03kPLfUq+Hf4jBU3Dkq
8ISlSAiqQ/yX/5abFM99yuEQBDdvY2AJj25zPN8X67wIA9dgahDgOPtY2yCDa5p/xuJlLSwFvtsZ
lnsMNh0GjyaH5zwfWT0AmCUXOhEIumTIkZKQyEQUt1ucxNKr2dxps93BRoAHdJmXeuKX8HEI/j6J
/vd49x/RjxLGajmj3WenOj5fDRk4DgLYbDhHsO77RClsBMu3J4sPpcDbbMMXB7d/ZzWP3F8++gw7
RIoK3nVH7UVeobYX6v8oZYQrqKWqTTnPSxCtHYIDcCgL3cxrhf9DJyUcn8SlKkbz5KriClp61xgR
ZmvyqZfMXYi6BETiOtVsfOCg3AjUAnwvloF4LXvlgd/wWQc0GLZyAMxCVRxsFdkY3fcc+D0P37Mr
E3jOVbEe6Z+2Dmi02xqPAk9tfk4apCYJrBJMdlPp122LZ4SikpRtiildA700rUmhVNnSu+zrwWcK
mx72UKC1GBz/HA+wq4iLwKg3tRcOnTGaqHZuMSLZRhnofiWAvKZZWauB/Jyyx+5fvTIMvJaYrJt2
UqejZjWddX3lPhShH6K+A8i8y31wOsq0S3r+SIDrvkzfInEkuYSGXDAtezAd1JNOWtzagJbWBdZ+
RoXlp4REdFzhztLegKJQ5tfipi3crAYmhUkm7K63JgNIvuxXFubcsxIUh+ugK0lVgJ4xthzaDSZN
jZv3yH7IU/Lrgem99wJ6QiRWklzTa8t476gMCcWZ3vJFc7UBlLA2ZnNYJJLQQ0bi2h5ZlXgQwnm5
DVDP8b7G9pmGOfRk3SE+lv9ZlyjaSpSMb5L4luqbp9nJXxfpwlyWqa85+cNpB7cXxFwzoqwSqbQ/
FGqmpdSBwQcJ6Faiak8WDceZSyFMSFk1EP4FSSIhjuvRIaV4cGUNPFewkez4OvTSmeLg5chz1c3U
HOA4FHaTqf1lMphkhSOT1dyb7y+xiYU7jvtAggeRQLH/IcNHMeiQN9xsRmJLJfnunT3GOqpX+ccR
kZQU9J5Qfsck8BG6YM8+HZ5zP3D6211dcz/xa1JYP4RmpEb7V8H4pq1PqNDGmM0oxYA7P1Yg+FiV
acm453E6fiwKjCmuxurLSYBbnvzhdbeCpHxwOG8hULyEJ+amA+bsKcdR7jPELFxEaQSTYefF5Khz
I7YsQySVNPARNae6uzerFi8Zm8lcCgvZ9DQZVX1jjpnl/HqCSikQ4aWCWw7Ouk2paLjVF0ywkatT
UjqEpcIlqH9P7pLlprJ8+8CwgapJhRR2ROVFFRbRSnDs/lBndqlsKLaXYz/0wd80rgVRbwH6nzC3
UIEVlDkrXWnMVLEX5V/m9xhMvcVwPzOIzpJ8DZrPW9pUVnzntgAgqKctOgANRV0wMzZ+jd0v2ZSq
jCOkxWDYHtj7YtVH4AB+EjaX/EIgXByFqH5QwZ/F1P96PFdRhPYODsHNjITei0h+a2uDynCSKV+q
Gie6AU1lKvNxOeuguRLQXbuOWIEYuYAJ+B9cHQkgyIIbiyQU0SOOxYiDFQwEGb+fzre0D53FHnI9
ZC5s6Mh4Y1HyteNk8+5TFjFYNrWi7ZcKjcX4UOPrIFUuhMx96VD5QtfynDC46ry1PHmnLI/x0QC2
WiLjUxygIcGrldKzpQC9gfdAsLP7ma4dn+hsiaAqZhcEXWjDjrmW5pFWL8Ul5y04y17ApDkmtSKJ
9TJN71iGXYgQqAdUL+sMH/55PPG8dVudGgIhQJBeWPrikeEAVL6Pa+TInqKUuNTbfHbyZa9oyjib
xwgkOOVh6iGpKcSdalRrPSnotaOkde4c/1fiSU6fBbqsvHpEBDNtcrt63+X2eos4frR1B5N4gvs1
sLUOm79enzuIVJPC3+KQ5tTBIMJRPk5+mz7VpS+i2D3kae2bt7HjV1EXRFaE9Pf3WQhK+E9dtQ5d
Zg+0pFB3AEK0Wv8AewggmAHegnxC3E8pAKKJ22kLpKuVTLxxPkVlITZEwhx4jAXG960POa5yz7G2
WQyYUfFnXVta9WaO6WDzOsJcegtKqSisCtPXJY7IjJWlCGIma2kqoOF4DCWxmgKHFTUTVHeovv2e
S0dm1D5t3hzgGcsJoq13+ySiIb0AVKRXDd1w1kUauMcfIF4bSboDxOsVzazGjUYf0x2s1uIhoonK
zTXJ5u6G3u2ReTtsifh2G0/msi3/lNbY0MwaVGsqMu9ijiUS00qCdA/nw3q5PRpSFBcSFxk7ZZd8
rpHWxwTNQh7ykLrly2PCtUPoPL+wtGTcdATvb9etrT2qNjDQXfTnSLgrlXb1ymQD4xzDa8Tc/vNH
6NqnoHK0ZLZm2QlTsLDmAbsz20YsIOdZduD7K9YriAXoq2TxVd7V3x6ShWef/zTQiCJQggPF/rA8
4G5Y1Ls68pwW1MPbYBiMA0YSwqvwYwxeR7dElDgSI3suZ809SnNcpDHuTDszmVCC9ZJr/I8I7/G3
sPsqd7BmGo/RUdxloiTjOKZSaGAPU/EXn4a/Ic3bnHcMZ919KhebCV0LzX2k7CxfA8zChuOK+tn7
0RFsW+ni/VUl/L+zcKjbq/gjGZLD9K6+gUy5mwIQOq+LTFpk/Oc7DQnYSjUI7X/MHaADyeZnZCrn
z7NoV4GDRtLxBkSPZDsoH/Pwd+5fcmpRk3VJYaMRCeDNPir0SZq6mZ+W+GNeO77SZLqmw+qF/J/9
3bQtAhxIAhGJmlKuL4367OeAfjoaJhlS+onJKVuXLYM3rwltOxRJcnW743qvVgiYWEKAudj9y1eG
ND8bZLkWrrjcjEQtXtfjatLfsqGQt3P1P1r3I7EregFgXveSBs1pl4AUP8DXIJBOXpBkGMSR27WP
Pwk9qIW+3NKGWkKrT29jD4OExneXxFfN0Vwu/Qf04kfzJD0NzEBOVOpnoMILqB9RuN0vEGKS0vOZ
ywglg3edIiHxPAd46rFAE5u26TQF529MaBdn/9tnorN1dD5sfPaGr/g6qbNxuf6/tfODW6azpSAx
nMwBNeygHtoOkI8qJr/cYUCd4CYAJRdOAwGbl+GH04PLR2u/Wh9OKvO0jutEtM2e1TXhLFa1Vjtp
+wgIX+VhfOwXl4cWgihCbuSKp2pvKWkwf+Odmr4PG/ZPgk+9dOr8QLZ28R7lAUaaoJeh5VrrkewS
oxkBgAQ0V0X5U+0fRwBC770fvIskb14NU+8/2zNodKAhqDePJwUb/0J5pjJhbfjjOic0fzpgpCgF
Zreibx4TLEPHspE8Ob7y7ka8zGV8HJdQcl83WiuGhctTeuM6eZ1SXgLTgmN+p6jbMpdGusOc6Jt5
fh2WPlMo/38gyRkoPvYyMniXhVyX/5mVBeBFr2Ehew0NtEdwMzLNuQ6GMcPtvwpfNlb7sMl/qB7+
GhRZvbo8NEmizTBWxey9JrN7URwoOsbt+DN9kC+at7p1Hf55sdPStThYKXlpq5JqmKUlgyFL6N45
f2wRRpM2H9fqOBQhn73QDOphs/0lZMj09G/5aeyAySsEONpnv9ixh9QcsWhKiiR5TtUq1mhW6tPz
ajW7/cpPsANSUKSDPab150wUk0hmVsvDLddaJCKqCfbPdp3mdLSZRTA6N0qnLWucNQnJk12TojaG
YJjDJ0+2QA1o2DozdnJP600uhSF7wzBdYsjLNn1RxlP+SPyNDGmogqfPYfKUii9dYBRzKVKjjR7Q
oo1Wm0Aklc9qu/QBBQReQ2kvyl91UiypvStogFq3TD7YjJMlEJYO+J1w8P1sHnXYle+POkBX7ncT
x6hMXye+ANQPAtv2HQyip85R85ILOX2rCMtABlu9gMzNiuAx39gn9zo4efXae6YqfS9EyduFIy4I
XtDPF05FZ8WvaS6ZfVDkXOGwlRybLjJOZUyFyLdNWmBSSleYziYOLZkM1S7e/qZAQxB+/L23RqWV
LGEToePlxhoa0gBzTfAHS43/bgisVrhnVV5EB9IIwsQYGv8GDwgS1KW4m+MgaDUm/JBnKuxSFi5q
YaRvyNqWLBTUlj081dxynibrd461epZBArdo36+OGrHUyZ6fdLSJGkYjXfyOMsc2g/k2DdiChqyf
3r6F8Sxogs++Fvo2RXXUsjsJYLhejceTWKKziO8oV7qsjudNPG43g4RpoGVnZ5kXVDSU04RgWCJv
E37CzHIzUT4T6Md08pomgSzSqUtigP8bttXfZrqFCV4O7yx/1cNxG9cxtHUhVboLAPvSoWzqmqzG
kUOMtCV7nEhr5zsEL8QvbYRz3p/Q0NmLH0Ceyis6ORqHIeYns03k4sTK6ygqUlnReoMM0HyVMvWI
MW+9L+t8sV3ZXeGkhRg839Czn99WXXGNZa/SJhG2gzAxdJPM1yxuvSyPZ+9hXJAy6SYQwoGYzI36
wSUBaTe0jvP5+EKk+qfahzPiRL3H7ITvunWyDXmQzVd7luj1CK2fS8P+S7eSCtMbj8Tzgk/6Bufr
qUQwvQOv3TU1JLRq4ofFi5ue3vYwDa1sFxoOtmcxdM4R+mPRBL1GlNNYFoEmt0TxcCPEO1HUuN/3
0GFzi6VvYuzgK+XrFNWcIZpPt6ZzFIzZSTHEN6M9HZsdrX+KfwELAS6ONm0fO+/WB7vmYjv1ExfE
QQY3kOjZBcMILZEQojbC40fgUlYWKo9CrCJPoNXd2xQjCiehS7vfWjtc3ASCDxmhB3/+Yjy5XmV2
3AIUbgcKt0meUbc+6HjpqCGQnR1gWbcYzbM9fTfBPIfkpMF30s8vwzcn7k+Nhda23TeqYJ/y402o
9SnvMJ5WYCSRHs/dI8b8Mw9Tus2E3M8KZiwD3Vv/JL/1EzDeQZqeNcp6VTtWQA4LW7Ohu6oywG7/
35ZSe/NYo+8m5OdArgL2EFr88SICSwsmRHDw22KU5qSaNri5/b/Ma6y325mzBlTbVrFdomTf+Jhq
zhWCorkfVhiR9lTMlwPnEds/5rrsw4CwfQFbMZ5vFKfnwWJkgXeJIWeJVrzkXoFk2auNA+ECRxwD
g/jTAS/Bg1jlmaEefectBfAKlSmAGLG36soKM6T3334SktZ0IB4a+gW1GRO5BWusakEtxAEHqvaF
kBLd3TiCrk2whxs83hZM6rizXs6g//fLUgOcl+4N3dDmQ11n4OsyVwefwHCq/YFdKbJ+eWX4Zuk8
TAeip+nqCCpPyy1EK0iDZIGcg8K4wvnS1xEEr67iFVrbg2fYuC73E126syqFeT+bXUNLCh0svIqq
P9cYz7gFZFrfDtjgjlZdrxGD6/f9a82FMKuHXdIgP+wDWJhUixnqzPaiE/dtFk3CvI+DU+zj290D
CAky9yI+9DgydqnBg2ob/gMLi7jm9Fmtme8Swh21CQlg4Z2r2RbTCI+aV2M+8sutiQ5GtURxaCiH
G7L7tXyWNGewoQyhIZMz/Geu0i7Pv8ORpsI/eSxY9DsBowRmI4HF+Ao0F83Abh5+BU7vSdyd6izw
W1312Ob67nbn7pMY1Sq5R7AjN8Vr1jO5+MgtqBKRIUB/RWH27KSolC0Ll+WIyid8TBsQjG9diCqs
2jK0gDxyJoOykjUN5YcsPLCKjoZdZ0NLKbQdw8sZd6C6v/Zq220Q9SYAImzoht2ML++9ADwCpqG/
uClGHhahnxzcP9sP8KGZrknqpSvfNofobs5s6PkW5smyp+p7y/V+RvmjFE8QTLvMI57YM0NzQtyD
JjBBshfrc931wWq+y5XsuP/iR3TDZKjy3gBrynP+C7CroSY/3+yyynP2nAVi/d/s34j+grCdLO+9
f723GvAIwXe5uWR+dGEQx2nAS1zGCv1BfvapkFSukPQZajy99aKQIZaapztipmvt4W2XoZGGPi/p
3LrHjAhrJX9Zy+Kac7YYfnDDlpfUnTsYsnxvzb4kZoHkDlfIjEeW/UMyePfLT3frsZPxHPAxTP3k
s4D2X4ZLqRGo0/nPLM9oVDk8I1OUnreuUrHGgfbpMNyxDkxCH9lKZASNCYGc0/+5XAKHefs7iOSn
aAx2awSrFhTwth5yyicuboB2rDPODHQWBv9jkQOyTKzSzgafpFuDpS9sxcVj7/bEFbw4tF9xH5KO
pmqsWx0Y0lnqLw9XKo+A30FzckTitLLp/zmDUT4L9JCMMd7OuB5gBpI3ZrYI30InbMLgjGFci8U2
6V1jS1txwKI0p24/4+YXSDjusH7rQ6jSE0utIVZejHaY5sCCoBU9/aWg3gErK79jojxuNhq57xI6
1DCfMcLCZv+/jWXYtD0ZU9z3Bql7kR0hR/BWrc5zUP+yCw4srn09SI0WXojFItbkM0539eu7z5bm
CYkLvpHY2z8YIuUDxm+MobgpkiLfc5u6flaOzuiBuXf052c7Fk0dTs512a3/8n4pvPFxP0SARsF7
QvcJ/TmMf6YPYtqz8at5L182j9PW7A4u5zIP68ddZ59N14vZ8smm2WX+IWhRl2PAWDLW++4r0Xvb
q+Plm80hWeZFr7N4wSFGZ3VrJnh9sohUvehwct52sCT9804N9n7uXOP/rncQ/WgmJ9fgnfMB/CoG
AE96yehU3aPfXb9oEJY4htC04d0BG8h/9yK4bNmIN9VpsZcLkp/B+EmmWXiUOYgFULSLdNEW0Fjh
GzyTvYTOs5Avh3P4U6NB3uhRD5aq4d+EbM3khE3j6ZEgcoFE1W/Sjizhg3HJValvA4Fj1T+8hEIi
Y74Z1PZakAZtY+ElgH7PLBte+JFZ1qYlwjjSfgqbEbAwmRY943Cpmrd3+ulZexQgTVyC6lHCB82Z
5lyuxpXQeOGodvW89T0Y67GLR8IG62b3khIlkxy0ZJOfroVb8FI6Cc6rKodmyFoD6Wo8c5CyRrPZ
L9IG4s/uMGNuixDn8Fl1eg6qfaIDieBDSxSnShiOchgv4encEG5WaetkM8RQrfoGleSzWK4GA4Hg
nFULf6nW5DXcfliUYu3l0/x4ZPw6ti1ReCWGvAbLX9DWn0wNXM7XrpU9NRyJ13VU4/Rn1j6TXgOR
IntALYGTTD0Oylb5tA06j/Ae0JYbTZV9Jpu3fPdLUwUT4oWjzJyK73J0xhtfw5KtIy+aRClkq6VW
yxpQinFteJ6Gtm3YMi4Y9D68yajtDlvZD4W551GMyFpP++h/YkYJMG+7Q4rpaLjZ7cVzet0CY6oK
ptDZurqfRVkkm1bw4zpwZlM2SQeJukX6ZByj+zb7jn02g4TDAs6+C+6sr3TzraPXI/URavPiTkgl
ygcbDcTF7C8mFzChZLU9MBj5jFauVHB6FJ5IuK2yy76gNWsnofAcTwsTNVCknUyErffEjaMoH2d/
b7BZc/yhhzthOfthHZay6sVKhz3q+Q4ORtCNhicc6iXXWJYg085mmpvPPd+IxoW0X6i41wLpx1X2
4V0CZ90585EG01SUAN8fliNCwRV+Q5iOimEI5tThBE067jYMZysef7mPwSwtgN9Z230NWxYMhZbY
RAyXVqtSPtF5fs5YuWzRTBZopHP5iGoGOK6Pe8/pcM8sj6Wb9oTblX0zxIrZPNpbNoTKaTsBX1j1
E9MCzmebuf0GmSFcfr85TiYXFJ0RqBvR5L/rTZngZmc6XgUA4OlGf4/wl3VC3GApdtKYuX5YcGg1
eNBV8NNaAcxAROL+gYzvhYnwzkUqNs+dtpe4QbXfECbFiMm8JRcP2wC9Cc3WeiZY8x/NBNojfWjL
1qLQpxw4ogDU/s+gv/LPOKHWsaptbyRPJweWYvmApkYDv4GN5ux3pR411zKWRxedNaVtbhsA4yF/
mI4f/61TIIObHuJvFkQY1zI0BXTjkEEKiQyDTUFOx+uoLGGJqCMha1p8CBt6eIXiMUBETwCqHLwn
cebr67xTMDGM5qyRAZetjm6O2rmA8AckFFjuXPvSlZSqqLtb2ElbtMI9cmDHKK4fWu83eUWpjk/M
bICBQ8MIQE/gnzwSMPee1JOErmg/hbtD/0agjw3xoK6UJfX0IiBeBuftaglh1bOgLUKeaBmWOn5A
zBNqJGPrWVZaVFF0tEHfKM0hItaLDsR1cVT35YnOYsn2txLufJAtFZYyQlw86buemgmuwDW5E84e
pqZr+R1e3zu8Bdgr+jZ+/CxPdTf0qBQ1CC42eiTmkbhrxWPz43CgdE8e9GOnLMHpsC5I/utV4JnV
lB2Z0qitzzZw3XTfHA4+dzqcZmJml3skMVN+Ao6Cbn+PzHjQhrAVLwsRxl4xSMF41NeemLkzlU0/
km/0e0AJW/gY4cPh5232i4pikYZ8CNq1dHPj7XaGoEiHyvEvJgo4Pp17pwanzEfcsAuGD7ggcRXc
oiMLEZHfbKv29w2L0w6hf+NhD9lXsXxneh4eENbIwBaIa83QVgmH1aSM3rxh6bYPDoyv9aK4Om1I
WYIJWeSjYpyrLcfp4htRmrNtVrzsPanRSuYdqqaHtZ0Yob2qO/PKpvC/Iz/Yd6bFlaw9bRUszhXf
ufzPyLhOW5eZCal7sU/2fUBadRx11nWld2/HBN7LWBdMN10zC8/a1RDvuzfOKCuKVYy3b5WgF81o
vYq+eMnBr5sTgJJ5bLoOSRWR7N7QDkYJEvSjk+cgMOAbTEOUkTHGFINOT3HvJY7mUURgxGg5Apr2
yrEZA1I4nwedIWkOB9ScnJjwiIoL5WR0jf0RXEy/OxCtgnpWQ5jZnLDGuhfaxKxW/5mNC71qn7WN
wcKd7Y3jGwY/ATzmtQmr4deLdr5HacpH621OJ6bmtBSFT1vHHgkif1M8/zkH8DQEiLiRxnWghT4j
8+dd9PHDem8psDs1aTRzesd63HzqpvHruNdkW2I5iFftC5gxPbv5WI63/16CUi6sBaeuoI2ItOeh
IRYm/QcrJ57TVmwTltmVbNGQmr8CrHpPaPthzrKjOYvpYxRXiyOTJUuXRf1lhAqM47fAdJ/5hbui
kE10fMYXtx7QCMq2qPbfqmKCAs34Q5Q9K2KVvtikxZ9DjHGpJaxtHu5Swpg0MYRNkFC+ctkK0q2m
FrwkK88j+rv0qmJhG1Urvn7TLOO8W0Gqehzspsr0C/f+FVa85Bt3fZgDu7XSPXlIvlG1b2iyHlRH
qeHJClCRtvIqv4bF4NXja5v2lXO3h0pcD+W1EtsU2XAilf5uUGjuPUc3EV5Jrk0nPQ0cgAve8nFA
PjVLWrrlnNYxDrnYqlEvpiuTn6MPpDmdpBEGrC9m1IYRSNLw83mKMKDqRbYAKtQ2gBChKXE/TqNW
7auAv+G2I58E/H85rCUB04MBKdDIJbC+UOmNHc9zz1bSW1ALfq+NRIrq4v5b8DCJLVWKciObT8eJ
T/SvhKoOlky0GgvqDXzF37hDTl48IvSu6dZnFn1OL0voBAejdRK/cTtuQSSPbnHffedy/wu9pKN7
OhqYHnGeC1ZMQML1T3tnvJZVl1R/aloSWgU+7rMOeYSTocELh/nmfNGloXnx7yvSEU+yaMveULNz
7uUcC/Xkon1qA+8FfJ42cPAesTxvAOgSVFrVHZJsm+BkA6pxgx1ZZdvAgNV+KwKJTS69L2xUX9y9
JTalk+tCaEfq2NzOf7vMsNxtksEBp/gbsY6/UMY6U4WFFVFZui9Zt6/rUb9MCg/5LYt1au7BsrqI
mTkmk+QBoOfAPQX2vzufmqFF0I8KORgcDZnaKHujCfEzo8RE+C23ffsmTYRn/fv+hMGHqQbSHxls
owwvye9nqEGfRNnuPDSkX/J/1ILCkl7BQDurl7F9fet6XymW4nq7DkwJt0wUSDx85ol8CNVgHr6L
utw4L0qdPzrjAziLLHh2sUqFEGIT9FmV6KoB5QP9khPFGLrImAof8jQTb0QOhe4eOT7EhP4481cj
5D00bzIwBHvldRB9kO84U2IvCbD9s6ML/ThgB9/Tib8C87WUgDrTOpa3YnB919GG3dwA0DhJNd/h
ZZ8SYTw5fp+IIW1X5cHPdYAK9+O+CBSOyDnlGVCJZAICwzhSLEXIDCsoo7xp7lg251HKjV3PtnSi
3xDZ5UJ2+hcFMb9oHK6hevISgkeCvXbZnwEsIlEGVzbZWmKPnyfEEKdTPssKayrWD7B+hWqt+wHH
BG97th5xNhAPBovZHd9f11sS4EE0fn8ymqJU61LMp4fFiz7sA8lg/ZSWuaYZl9L7Iu5jj+4RWlwP
SjHkOo+/yBXL39l+VkpEaYjlTLpNHuXIUdgB3z0pHR4V4a5OQWy4P0l50vMuteegJ/r83zPZBaKu
dRR9EV5anD7G/iJSLn8SaKz0UoBl+cfWvaYe8By1k2RvkO4e5s/nQod/V35csRimg3YZ3rf1Dxc6
eGJqFCXOS05Y1vNRb2hcruiZ2uA5dBdqcgHqRTRP3W9Q4sdkKiiRARr2+DsNNvIpwo8+jSoCNTNq
nOBYP8ON2XfVlSpH1IVwHMdLsiHrJ6uffIJNb7ir2DJDTAqMzWY6qoVyjbSsW1pW8vehPHqXJTU0
gb+/NgK0ZoXeJ/4xCj03v0ka9RlAkz7y10BmRahd9aaUq2pWxOwSH/y2D58iHo+4vdX2JbHecw9Y
6E+14aOS04Zy0vDFftdKgybtRZ5af9Wl6EM7FHAzgskHWO6En8Zyf2MpWxPSDAWln8l7UYzHa5U3
MpJCBcWmWACJusYVfMEkg9JgtosTrx3ydzVTpNUsJUrJ7Jpo9pAO3N+7IGCHFaUR5hGbIR3paNil
707Dq19iKvvw2M9CVDTKUkbTGHVpmN9eZzNclPi8xgo1BE91gitlcpXmXBw5OaItvENlPS//dIOB
tSqtuI6Q1lq3FalB49Jp4geGXI9GAjO4eET0YFzZUFjFJ1y1OGjAXsKk7hPzs5qaJLpTuolb8dMF
ErQ9nvlKkXPdxxnJf+CPZrz61yzqQRfZasFSH55LsPVX+ZHwkki2SnLPOgfT+zbxY2BHyvlbyZda
oyiAyTZ/8E6RlYw6NnP6VTXhP4sjJhLfTDZZIISB0AV9oD3w0pmBQOAIyGoBbRVr0i3wgQkKIHsl
XejZmM4pVTKyPlyMvB24v+sz6sy4Ms5ocmQ6mpciTuZYFglybTdRVVaFAlfIk8UZfq4AVviNAUhb
tssyR2zgaH+/6OTlItGl+6tYg/Rk86+0OztWUbwazR1l+TR5SatTvx8SwEuwHv3ine4tHadRwoZe
rybnCgoJu04C/2lC5jcFqQmX+RTxFJeIftkQ1TEMOWOverLRlvLo/BnXXPIh5fBDC78d7yW53t2J
n50BPOC+yXmPCLfT4CAD9Rqm/hoX7ahuJ5diQXYvOywNVokSGNTfObIXf3DARUjWdgW8rhmfwTX8
11jV/+iF7z2liGTMHj6sRBEdkkPz+QVAJiQr6dMX0+VArOKv2gTt2bd/Yv3fbAK+n/wz2NePjOLA
y/YyaRQ9Kpvk+THnc3S/qMgdgoqkOcfiXa92YaJB2uSd7GD4An7ZVAFNfoaJF6PNPWB92dCBqo/G
rMQAuGpmO/VwELWlMJK2++sXRf2swUfFi2S9gdRZGD9B8tEfNRU24wKbI6xx0oiY9jvjn4w4ij0L
gqitpHW4rUERJQTXGxTd8pKvh/mcoQHoyQmXv3yUHudEkFiZmfoka4+nhiYWqZjVOdbAC+ncBKLi
eRqYXmWMP0X3pVKCfIejg5SOCJKJfwmrEcl0txh2Xt6SWMKJE1LgOj383zMAFJgljeijJUqmnqyx
RW7Oof0Ufu6vjOaM+nTpFCujT8tb8c9wQCmReJuCVommMMwa5Qbfgf+fPOkKuAQj3ffAS0CFrmzB
NOL2WiuWB/DZOiBeLC+L3XpkRDv9jBGkKLYV78iKuLJcT/TxRLIZHwJotF3Cgk1aiFTbh2+F2fDd
ojdqsCthTKAdkS1JWeRqLhQyHgLlz1ddclerhJQZHQzfRqeEdYGdyPHEqMuMKz8SKaU1iGDW7xYa
2ByluWcP54rX5sONdIdHNVfmptWXWRLR5GujdwCUW/MYz6i7cweF+0Wm9Rbfc5Jfu8le0pZvhWmr
Rh90Lta1eteXAz7XhyJ6tvCUe11lPt9p/LHM24fTCWqIsdPGnrUv3xIflzQRzlbmvXHt2ExyvPJZ
Fd7wKqWadjCmmb1isoHfqWi65yIwl6o4uFy8MisLynGEF4cXtXF//6+BptHrGXOlgiMnentoweTX
DKRxA9BhBB4YGLGJwNFyA3fqAj3WDCuHyDs9JH0Fs697fswaY271v+MKt53NusAjkcdiGi0ygyjY
wcq8Veb22JKjtrxC9kho3pTckrm79K+63SwRY38ETptSk55Nt7UWrqiVpJTRlbfJfIhvDyCYIA0h
VD9dheRrq7vYAAVDCxCwQGuUqmekvUiXK5zh2wzSIq5ebeXz57ZRhV1aw6cJdyzTJYpj1EHOisFA
mbwfT1vc5xbOmfPV5QFuUNSnO6ya5ad7k6MW5UmPYVtTH/bqIn+YTxF30WaAF1QyjsnfGKts4yKr
cQ6991f0w43BPSJRXwaw/4p7GAe4cprcaexUQPl9ifGj1wO/WqztkLG+9IofuOdRy0oi4n4rSRug
ukK8DO3shHXeZIjhCiBVzWfQAhqwMG1YBqJ5DCQQlePZ65iGPbLjLt3SWbyjyUAf00fgPugfSlHv
Tf1C58ee42f9aH9YGac5sNIFVJlkG/herFGSV6scFzx0LMK+TRarRXx2nchDRgHy+35tMbJdXFwL
R4qgfAv/lKAz9sC9/gzHeHuP1g6Eh5t5xSxNu9+C4wbUcD5KCd2brNEj9nyRCEeTtzaMhDnlka/+
wHfFmzG+7+BnvUfb0YwDI3vuCDT4u9mz2XSjLSjL12srcGXzepJ3ijvnGzMU9s7cmx+o30HceWDh
2DPoRbCoQl11VjNAuGynqSc5nX7tAlqW+U+Srah/Wp+eCcfEv81EAKtlM1ATsl40aDdW7wPjnd1d
ffx8oJnCqsqmTA92Y7wE1kD2Aw98iGJ95RvDacPa5SZg/NkdamqzKb6EkolbnwZ5rchV75SWhPyC
kU/YI6P3XzCa9MPn392Y4DNR2Sr/1PU+wS2sRAa5gOH4HCrIw7YOoS7en1qBar1OCHZrm6fgXTe+
Pe9QhJUjPrV4bVRQmVUKlNMzyoiQjCUT1a1bQxdMNzXX7SsJ7hyYX91fb0IjbpI3Laxc+aFpVuww
naX+FCjOqZWvgAMci602ZhghLsAZPmiTzTtsPEkNlPsiY4zfSGeQDDnjbu3F0wZ7QNdMmgm8IDYk
RFLk85NF1tFRZ/Dn5mUNTdJx9PlxZkeQ2+rotz1jvqwUvMDXSuchDqCH+EPcadLUvA6Plky47Tvu
knewxcjoQRr+vahdceTlUeFqfzRDVIY8U/qYpMbVMPXAT5bPPJNG9vSgCDrh+B4dlh6wPnr+PilS
eRlSVmrbHrr9X7jT0NwEYaJJ0wi5F82TgILCyf8jfahvetOzGgIS0L72V+qdYV2L2ZNl1NsPACMv
mt7f+v1fHzpGvi/CHi4xQOwuGK3UdMqNVVxKbyG5e6NAa5ct4b4aecQ5HOt3nMTuYAFzT1Nj4/Zh
Cf6vPKNP4qa4/ubxAoaaFcTP7XrIrXVZu7wfkfNV2Mvg4NmpSBjEKTb/2Mqq4slvwipPCvzgA4yu
fTnannT/txb64GoBJupwf6ZYVI0It7gYnqda1sd1TwubPehPqDGCzy1EoxBCSFZGc4csBm0eulfg
IMQtYgx99xS278Rzz2ZPMuwKdZkvtKS5YFXSASftSnk1sSzS4b1TJvUUK0ReIbIBUUfz+J3etWnw
VBPRI3if1LAGmNRCC1zr8HPJRepGtdEl3rU9OWHt1+P7eMYJqO0zVueUx4dJI9ndET3WuhDt4I5r
foPUdPSoSMeXRrWXkVPosoZhlb8t01052eyvPdqK/Jxpral+RYwV95Xo2QJr/KhQptKKPqjfs3XJ
NzVaDHRn3MrZapoooiDaYbtXiNOHEc1pv6+djEy3F2GCFAl4DQUJ/aKlI6J2TvMAx2ZPJKoJbA+G
bRRuLO/QwH2xXmmAjPlzeXDo+HRS0mo2tXWen6UJ05MYugOcAWRaxuZT1G48aB2gvW/RME7xDCcY
tvafbBHlJvqnd7WxfrzLOTFGOFI6xUn06ah5bOVVbKdWQAvPNPFHB3I2Sc7DmMc3gTN8iI8+Tyl6
FHHQ/7VG/Dg8mgO2r3Spdk2KzaBnqtZqLpTsrFAtuazDvEe9ZBI+tsWl4Tzk/WKhP242VttB/Hb4
7N5f6oE2IH1Te5rmrDj7WHvP+R4RRG7TstZGr5z2/nQY7ixH6ObQB8xVb/EjYbll5ZCy7+tSNgZD
1ZD71m9bHrOE1whDANhc7WWBdkKEyDjYOZs+eYNMgcws7vehfjgsW5rR99+HK2GF7N2p33pFa/WT
x1BCYYag6RN73ymNLDDCZH+B7m4uJkvjkHe3UihLkU2/ZyH2Xec7X6CY71kg5HVt12FAOtbXJjNI
NCh09OD4StHcz3OL9ms88IBnDF5v0LikmvGAZx+o5HPB60HF4Xk+vpNFCdLX+W7kifGStSqYes7A
ubTL0k9FcK/+16GiGLnXxdF9T7fPaQxywHMHYJ0I4LThE8QCTeoVbKhP4bDVTtoyPMGw1trDVukv
HygvwIxXjZI20PDCBlHEguZ28wBmoLXRbDYhjFpCSxRbZkRSCHBQrS0C1CxIXOmw3/qDEvoGNmmJ
uQ9rSOkEt9PDuY/9v2hYAm0JiMs4GNc4QVrBOOE+uTrALAuK0uU/WofOqSdh/OvfX8CbRUzoGnXg
k+erreKj+QWBoETYXu72LXkJckgIoY1+TqwfwRCxH5EQFoTTrzg12czDLWkHM8LuBIsiSZvbVxZW
6F9wzxXAtsJZobea/hXqzomy6oGDcyWjnGaA4HW55wZpqWRNUXECt44oCvOaVqbcvZXK68TzgdDb
5uLSEubnhU51W2LA51gCq2KepOVxvgM3C7yRphrKF1xSvSHy38t8g2hOIFkqVPoPV6sXkriaN5w6
6Ni9bIIyJGaauePDLrqI22jUAKtXMC3SySfYs/cdkMRr5KmI+2tozUByi4zxpN7pdH7bC+5eQxoa
XXecuG0PZHBOgC4RrHKMkIvQC1m40bn0cUNzCGGK5xDDO5B9cs2i4k2l4fkuQsKaDI1D2pcm+Zae
O9utNmLnUTbjxwP5mBOomZ0w2d91idY5KBGfktrGpjeJdWScThqpjitSQvYdhyp0JSMZuEGiDtUO
myl8MW0TuZXR07fYcGakymTK49nwCtBr0Aql5ZLEiRbW01Tb7sA02U8I7ZI3ORkTCQbuvkNEbVwI
tYSbIN7Y32hlDdhr+C41msPidAxhIikjLG4KDvVrTLo4AqJ1GMlm6/jIYinQB7vxLb+KSJmojvss
5V2srDyxA4qaD2Zti3WjweOp3qn8UPYKFtg6tnIxQllgI22n9goeclSO2tqe2iURT3lqSCe0veCE
GPP+nUyRa1grxlMcHZHUWZNyDcAKrl3pt2JcWm7w2DNRNLvovn/kDYl2/VxU8JPqPjh05DVpJT4w
LvRKos6ZShOYR9V50lVV+Eele1ddhA+2/9TKElSwUcDFx7aAzSZRdabwHUlMi591xjejsZ1NHUAr
VI03O/pmj9aTMyxFlxqhYF5n9YwrQgESDDPaWmMMR+Bldg5K+tnMS+ouTWUeNzTDTbKg404l0yIQ
hqx8zfUbtG4sknDChspBmbLChq8ED/B6l6ZToN1giogujVHH0hk69qsPzVRMkuPIoBQvQRARcRPQ
smROfXvJrDHDj749hH4GB5AcHdeuTZ8+ZwwKJftr61vgvGv/Bac0iOFcLRY/VZ67waEAyKHAi//s
bM7Ozhl84ypwwPGlaR0EYj1f+jaUkKIHxjGCs4kqsr9X5NXpvDVgi+U+V4JJ7+6fzdlWQEJ/qkMH
mrqwmf7ZA5TpOm8W3y3qozGR4AUryn4WzV2ptgBsxid5v8tl1pXF5HGMCcCBm4eVb5iSflYJhCHE
z1flZXrYVDfOqYoauqlnSfA7Yod+o6vrep8CEEtziHfFA7SZvcjHreR9ScOaeQpYRQLxNPCwr0so
dZHOyOMWMG3/Wk5EpVP8aaWiHx8ENyrcbPTKA1Qq/JgPvj38v54rcR/4GBDwINA3MQjRPDzCWrae
lAOrQ7ndNkUceapQF4S7LeG+LVU6ybMtdN5qkQipACa6V+PPu0qbxcP2t786c6hEObJuCs5s0Y+f
/kGz1jLx8aCmrNks84SEWOs0+bzqB2DPFq3TPPhy2D3st11SxjU1rifC1VPqsBAZ4QyIrXq5GHDW
agKcpONh31+fQoDrvrJQ8ynp6fhleCZgWlSoa7TiNXtuTCbmyjomaNmachyMQVwrkKps/MrO5TKJ
mjbpjiA6L3vkXu+qKetMeDNRwFTNjpv38zEsRWuK55KQUPyC715MpviPeawgUYNDOvUinXw5dG0A
+0W1bdzLjk6QvdpdMgZTh7MPm4+slwaA+M96mgOi3OIU1qMuvedEDfNKkvtasNfEQR5bQZFYkAuY
Q78ETPAhfvZcWP5tnR/+eFnD0mK6pogGxH7uEfbkjb8cXZNF59jPbdsWGLzAbpoloRm5vM29fOIt
Y4giS1EPqpZZAkqDkALoCKzJmDLzi0VLmcebPosFwfAfFsAIy25YPKD/84e8yISX2NwPyHsU7s39
K2FVucLESpKST8Hl3lPVza1c1LkuVguZ+5Q6wT5c0cqhECIp463HpFSmtrDMr8DEbfCyHai8NQbq
KwSPvJEfAwPdhHAt9KGB7uGvKfaY+lQpg0A/BIqk0Mib2E/BcDx4gfsUcNWfbe5BFMwljWlEyWz4
GDEt6N7jW7IYu7J6ICXQkdkuxM8IodbNFpJoyv1ZLYqimlg0PhVzU2aBsdIMiW/zpuNx8D0ieyAR
wPInAMJoVEPsaV8sWZanchQUrZXWqmeCCRGuNGY85KM0MUtyb7Qt00OrEtf0crIH1j578/6O7Hec
49wvMIenhRDCImva4dS+RPLor8aycoZ4W5AGhajDPjk8yw80+hQzz+ydnETAmcoQPa0Csmdy1i0o
1heySA9rob0m6CC4wo9KLSAlFlalLndVvk3VBEgsr9S5ymZfYaqAKSGDu7dCarTFpBjDr/v6NCRt
xj6j1xClsl0e5639RVLkCcf91kJzUW0Szn+2iRSnKXypdmnj52wZ0y/UyCyMT8hA9ylGJPs7swdw
5ZBIdzQiVVP0/sLI2yKWzgfkURm7uyQo17dLGdY3+RmzwEpGxJPEk3b2qYrjFK50fXj94XbHz7X7
skQcyK5T+1/+8VEsoL4R2AfNrDD01UQBT4Lh2JAY5QYuCHUI58qflhlsblnIPf0V5JXs1xXFxiqT
UMNffQSRytDY/VoaM0aHkIZGPoo3xekOJa0hj4eQys0UEOX8bwN2O0uDf7eXa+urRn6YKHadUoeo
LyIHcZM8s02Jz3SDVRyxQkhAIwmgy9xWBdumWAY/l/MdBvvV9xCjIiDA7hnnzjx2sljlHFZVUkOy
795zK6GpltcI7osG0fM8cdaEvPRhHc4jP4LCMJrfURD/+7TUY//nla7trw4bi8MrdfT+QcQdCihX
+PAPS9/SldIRzd4Rbska3xnORo/3wtgMbEkYIoSQR6XCAZIG5MZo94LWI7H8R8cSDv01zq5gV2Oy
K4QiNGLSb4RKxWn16OJ0C+iQZIkr+2CeFKZKz5u3lToJ6GWDkhfRlwaz6fqmE7uPZqYOxHAQjrns
/ONWCGctRBKJBJrRmOhrz5t2+ZnLg9OKkOd0ftmEFcbT5BlJC1//tFI97ljyL6BycDAaIF5z67PA
4Jyxw+p7FGYrHRDkLy3Cp+clKFdkHcjcwGW7wj7NyjjkalvvcFBZ3EJbLfKbk+OtwzEiuePTmN5E
FzMO2DwcTn+CQ7I+gaeT+j3xyGqcEzVlXOMwGvEQyJ/mcdFdVO5Ap6Y7EzKWqfcr4Uem8jzBYvvW
vaqxq9KbgddiJ7BU87LYFR1/0qzqkOM0KFKXI36a72uDKzmnM81HpgmgT5uAm4DhdVz41adPLH29
EYQlmgbxHm3dQUj25KPuh3IXe1WZ1zyBlpji8JvlAaiIBJMb7XxeJmy3AKke72hqECK3xe3c5LTx
Lc+RC14C+NxTNY6gInw8VsEYVgU9ee4zCpWtD4FE0Ic8J2f7VbOBWwpgCskUEmUmZqSEoqpCZwEo
96KT6qH2/f19d9Iz4mfasrNsEpHCtkfAEWhQcIBbF9UiFXhSM5aD6k49pPaEPdDTghmA97TTUbJC
zqSZADOZ3UH4NdWUwPzKT4FjW8LzT+XaiZmVkEUWt/qAJVxmnhJGmYx5CkvUqDJ0lU0s36MNM44q
pkJvW1vLWzG4hNBb/8LlJuCf47d9GNw0yyTBcFogd94NGcvqmSg/fDHdgVbQbkPyOiKt5jNB9g4h
c8X7vhDOUE+/+3V+JC/vLKKAet60F17Ys/TFwJOIyDDzVFgKDUcKPn8GbyJNAvvr583ZOtROis38
eV3mCCUWW3ZoZ5u/+Wc5uBd3fPCj4aBX+yoHvHy9D5EeDqKDKZkh61CEOym4NgU/WQncHUzSNU5R
OguL6s+3fCDLMP8txDqRUu8AskydzmjVZRXGZu6dK1ElCAV7mp/ADXIpFJRBPs6DhqW165JPd61K
AbfXMMKx0F94QBt1SBppsaoZGugEUqEKApv50Nq0q1x69rDEvy1NS9Nnu5E6yCgFEVdQHsMjj4OY
fcJa+mLeAqgs8nCc/Gm8ql3rR30ks/bHlaZh7xyDlXMnkjVhSp4nPaoC3KcT1QDP/kSc5wNDuQtX
hXmeJtaUTs3iCADhTZCaWXERZDTBMMdu8FO6TG9cnVz0/4hRKskS3oZ+7+VIQuDBIEByLOgwDaag
xU+4mjPkPwruZ/orAM9x2U17PpJeSjiduv5wUv48HeBae+/vm5uvnQo6TXjP/1hlgIGNVQHsRNi4
QvYJy9spS2upi7aIrAI3MSU7/gllH+vZNW7kfbvx78VLB3uW2tFQ1Poge3/rJ7IGoajgAbLHthi3
JyTMvOOwY5qbUaq6B/ru/DQCsZiWNc5gpCI0n6Afg6YnyZA1nr2KkihhYTp+b1G4EbEOtGtf6Ynx
yH3GTNRmEU9L3JcqUlG7B69n0U4BfGsBWbwAN7LlvguaHqOSRQfPeH501fnnhmSZxSG4NTP2JmYV
uuU7P0HO8pam3nEPJgPBJaThGU+Zl+ABYZ7FU0Q+rNP0WmHvo4MRc6XOAF4+tEbHQ1fAUld1oj2s
LzDhrHj6LXkU5jXgixcoXs1GH6xitsIPDiJHfEH/DOXLyhkJcyai3NqHvKlAGvl2qqnySOCElcm2
z7Kcq4Am1IvL118GmnKGKaBi9cE8yw4XyIBDQ7599lmCn087NmxrcFPrOxZMiFWdBbuuPzmgyLrw
lrUJJuz6d+Yj8TVo+8GA4PKfj9IxWXpmFM/GjPBckw6CEvxMlCF8ndkeF1mZn9IJVURZJBq5E5jN
PbzrTDv8T2zf7+oUUoIo9fuXSp/UDCpZu1zYTafzl9hImki3FJ0/J6+ff0aKG/Vwnwh+sSSfZ6du
FFYw315a6Lp5bvuf7xZKN0gaXPLXB7mG3rlAXmhMOvzjtZn0mwTppxJqp20UtkPCr2JaI1vUmNhI
gQG8OvNsDWFv9gjfwlsMVEqIIWFLW6sFLki+aJlkCc49bsyGfhkrhOpEHytkVeHDn3kz7wjKELU7
40ZNzIJ5nMYDAN/7LcmPl5O7pKdImiCbN8+TDvZ5FVnMaqJcBcUjaLx0jabq+LDpyy6CfGY7sty4
eP1wnw3rYtAXl2PeqQWuyARIKwRpc2c5UcAf7C7NZADHQeRPPzdLTcZILL/mdRrRqO/pnJsdArwc
HbQJO3iWmkNUccINzgTKglmVzMgPEoITYANP8+8aB2fhZ6u2Tm7Z/JjR6lstbbyOF9cYAKNhQeow
p5wCaGHBhWrOJvv1Y7pQbW7HT2or1j3dWHNBzYRkuTC0uD/STPZqUudStgNKBLTMoUuobVbcRK8T
xX8LVQkpHiKele/UvQb2g6IxEnWv9OXGWvA5BF94F1SLCrq9nLH/wewacr9/68hEZrzL0zoBw6Oa
ALx9gzNW2m4RwQ5QTqc1Y0/3zIwCHnuURXt64szvy8lMdxATUsOA9YSMgpeXRscmKe2mCyKvaTZu
PIV+99SabrmW6cxqgIx3bQw9/BUZ9VeZ5/aIYmpPgbEs8O4xyzRyMZp8jHC1lRcrqCv3bOcOcPrW
tRVD1BucPkaOmVoddEWuMGzY3y/wuK58CdizPOOndvoMsGv2B2EoLHf1TgFlfHhOsNn6LCFZBZjc
sTDd4ivNAfPPvgGRfkPHPnKcaqfagV0p1KyB5tV0LIcUaYJKQ19O+DJqzW40UNIXDQqSJ3t55v2B
8YnzKLpB0uMTXAZcyHnQLJ0GYhq0GZnECFF1VCdb4abZwR7sHsLg0PrCaX4Ivlg22zIo6C3C3Q6I
5jVgJmHJwNwSROFf7kJdBDmFrUzoExkF+6/7G6prt/lKLI5nfnxULGYsWDEKQf6TTkIjeOBFmoED
NwEuaAYjIWhVRp8bkgMDYTFpqmqofIlWXnAIwyRIn8IylHO//KUptLh3m6LnbG8P25acgP4eTxrx
/eT8TeM6W+MhBWLg+EpTzyVZ3Atao7wYQFTm7AZrylLwNMQiU6Z+XpR1F3IDX9GTvc+Bu+wC0Ja7
DCUfnG+VbCjCmnxVsjvSYXCfkIQXPW4d9CZvtHboaMnkI34weWGJ4hWf9vaYVOB7RqjpTNA7LTit
w5erpoM24SSuehUGD+z0LbH0KS+PgNJTvngEzGKO6ceuNUVgH8PK6hVdew9yLnpGhKYDehTTCejv
utDsGFgXfhIQNIr0e6BHK2zGeggAiEWAXssaiz61nFMCiY2BxpNA6QvR9f4EaNhmZzSCEobt1PES
oA8K6HRZ3TI1FXJegSCoSX0RqSh7UF0Sf0dvpERWCyqOYlsq3oS9uvcGoiipR1ZjGHBGKVtxalvr
i74awh/DewaDu3c2dL4OnbTm/yabZiWYEW9+iu4nY7mZ+mO6nre4SKO8pRK+fOyow0dbIxqYnDHu
Rw4nMToSUKXzqcQ12fBjOJjU0gCrULUd/UsFs+9PAkjFkO/rIVDi+4zipHS3ZkuhbXYahuF7qvNI
7TXoA2J5UqtVBsXO44TQi5hPdiZqVFVOqlOWCpQKoXC+YJDabDoOcFZYU+c4yU+ZTLGE1D7IwKse
t0cRgKfy1WiGpjnrXdHcjM2TXjhEMQIONup0CER8vaILPAFaZqWGhBdDFF6KpP/UhYGrBEmgATZt
9FMBScIFSoNu+srUR5R/Z6BYpiYVBrLDekzkbq4Jo7j5CRxNppggCaM9x78gIaU8lQ/r6xbTHzx3
7BByPqoBu7A4jVC/Lcd4kGTlFXzOM4YHzBpSJThFj+WbcNx8kM+SMODk4gAhC7ivI+cPGk9V2708
e0dhOqDkFfVk6eUxNcoH+lKuSK4DCQTb6MMM9n+4i9WJrYy39MJMjbpjXPAuFuKVW0eMCw0WDJOn
7hckyh72LfQNWMc+Ln4Yaq8Ehz1OCHxghMZ8CZCVzMw1pnNCm8O3hJn9T7Gd9d7F4MBqxUPWwyrm
Nu53d6Bc8SRGH9dW6CZZ0V9N8XcH3CaIc3V4/f1qxLUdIIUcc3Os5g3EVrQv04rTh5HfMIOpg9/i
MJRsx6n24eiKFcy+C+zeRb4zR56ueIelx8W5EAKpljkK1hujxVLyEC6rx8K0/iS3+QMCjL2EfQ0t
E4by+/nCMxv2FpefER2cO095XcxTHkkTipgNsyXVrg1Pzn3BUoHnVCs9YzO6y4SpTO+qJP4h9RGI
jzYDFfH9O0H47paJegLJ4NPCC1FISftEanlTPg5Z0lankdPNpMJNeMT1NCTNcuTRpcuLEBqd0zGw
utnXEGXyVWb0yyyKPMFLnd4pkCZTpMjv8J1lIfc8oAuufRIi1Oj/Qb6JrSmBGfdSVqMXHz6OMZFu
oBTWd4N0q1rt280mnBEVhQRTZXSnGfZFPmkX26z7ZzmZYICdLdDcCNtwuHfvIulrthgEuWuaD4Qi
D9nkROBQk4GE0PFPXr3L7IjbX/W+2x8OC1tIHC+HY+NISqVX91kIigGcxl//p2ShC3aROZ560gXw
+MAwDfa3HIvukdk43xAY0JYsCbl1a3ibforpW40CNY34qj+hHD+FZizy/mNe9DN+Hmc96ywSE2Gy
NIwk5UMOHFJmlZiNey4FxZfASy2anx11Ud7VodW5+KyWX7kOKQ654YAd2shY0U9jA0fRcp8kvpxO
J80abCr2CNmGx8jwUw/4gCB5NT5d9kyF+d9RchtCebOOoomFLamSCovuI9UnDApUbo02EpM/SKUe
d8Pfz1KpUlQRe/wImqxTvO/3otQ4rXjMPF8LlXjeHCC+4iKszj064769++VHDcCXjLQXKTvYgeN0
ja/ZyO7rqCOsbEaES/6P9O6OgBO/qbplVKG3CdJ3CBUGCmUUQglE8tj6bRd2pDl0Jf+oBAAaVHUc
YM/oOhoMYnEkh9dGgZ8L97y+y5uXHEwVeME7nzxpOrgmRSrI1CTJy2gA1b++/I46mjsR+ORIB9wt
O7nLY3Bw04LAARiQmmbtGnOkh/bU0/uDMY2hJFtdotB0V+YuKCZL+REA3boeVckb5xfU5F73rtP7
lrL00lGqBXSiwskbIE7JFAmUoWeU9Ycq+vK6XRfGWNVdcuiJsb8lYbcemJUXef6qfYgCsqsGfxaf
wwsfXSoStes/zs9xhf0aRZBjOMH1UalOt4LvTeVpIMvLMP0NPTESc9qhauxq2xLE/0o5vNXZFgZ2
7kNeStftKa5+3NM9PCKgBl90gTedM+doVTjUMRMB5q861Kim+mZyZxspop28vDXkHeygLHoYD0R7
M0W2bW8XAOnRnFbtyX2BdRQzlifZPW6yKjAB9tAlCO3bv889I+AqtN0hRw1Qi7m88TxzxHYYwjOw
M3Qt04hit+GvuC+IMr2EoshWro8Upg/zZBMI/kmuCJeSwsCozzNvJCwaIv6YjSveApVvy10ks1Vb
hz3NIp3FOuTCbTjmk4TLCWV9XtTzRXqJGM6Wg+kmEtwROkcce2C4IBl0g7QMDrisaHHEH3VFeWBO
e6yysOwvDi+VELX6McmalwjM2PD2aQUwu5hqptImtlEauabBpQZ9aH/EdgSJan2mR6+p33F4jB6n
j9E39nSSAOdqBHDmLl+FRoS2VoGsJONvo1XDuf9AHFn0IFPcE8BsIkq7AyeOi2EXnLcVx7JzG8Im
xRT6DHooctKHRzWSRKZRD0Ebja1v69GwoiejekmdnGgSnIMZl0TX94liiZ5BZeqBu9QGDRHGIfow
LIJd9h7b0e8mJqU+T4BGsxhwR0wqRVUkEd8LgVlfx4VayzpZWD49RRgf+QWbqP+EZychuEfEbXNl
l2yrlKlJJJmxt2pBiz96Z/XOV/7CfNdol+hupGDxSGuH4XiEAcwjVyP6j9u5ctQdiKktusczSCVJ
uVm1y/Jjjk11DsNI5bA0lqVL3boDa2Gz/sBaTNLKQRdaucv5AvZlIIz6ofA7ssQitjn5GGoTTQ2Q
UeCKkYIA7XWjGhCtlLqlkQupQBGvjDGyeg6ylERA8OlfSYatEc0BDzgnF1k23H8SgbVAg7SxWBuu
ZpXZJ3NmavLKGRue/gNEELTsd84jYP5lCvWLCNZsI+blhwy2YtNYHeCTBa5SxZPNckwMNgIxni3V
GlS35zlvpXUbU8HNm7jbj/pQoSQB4OjM2rgNtS3bP5lc1GNkXWCtE/0DxmTz/7mOHWfgjrTfxttF
Z6IhRKR+7vedyll/ja8JmnhgIqiiwYA8uTMfVLpcDQCTcGbNafQHeDt1E/Gewv+pkRlupF9+RVuG
yuJVSxY0skzSa5825s4wn/PvsGeyhZM3Mz8skhd3rMBszTG/MBg6dJTsn76ME5JTjVYfnBgdshTU
H97cVeqSwx1sShgXdc/teQJm0fROCIfcYMjw0xKt+mdj6JX2+T2TV74BzLpD4bKAYGU9OnX6g1C4
pgIE8BDyq/s++hys7ai522EQ4lB/4wBhJaSn1OnztbgNB36Mb3I8CX2M26PBug/Uisu9APiPtKXN
iHGyVUtEAxRCs1IKjxJllfCdfo+ZeHQ0wiGuYPGKApnn2oHXLwPvo1Bu/JEY6E4hLhoq9mgp1AFR
52of0jsv+DUpWvgHuakKZuQyFqroXUrmZiymY+XV9nHLR9tAe2k51ALkAP2Hf5i+t3CbvrDIcqAP
+AficPuNUVMA4QA5JedJe/CkEi9HKk2+kDZR92jUxZ+TcO79KUrwC+MGhH0HdfYK/ZMVWGMrUc9o
lAk7XgmKw1F8AZ9uDtai2rnBMvARKDZRw4H68qdFuI0vQCUVqjzHiJhO5EQlcBOwWxr7D6Dq/t/6
bqZflSoVFgxssbgUgGr6ipFW9qWLqpJdFUjj5dAEUo+ZB4HictdCpyJmbDwPP2wmmNCA6C51IZtJ
yp7kqbYuPBWAoSJBv/RC1ae/SAfUDpvlnlws1XIhX/Dgf5IufeqAa1fNyFUTMeNRZZvO+5lLFB8E
EKG8pUeT0eEHb4dHfP/iuWnzP+dd2ETt2OlDx80Hd/Xjf40DxZMXmG0M1EDhal2ubVC6qsW3VuSd
eoDvE8zSLC1eyABFeAJbd22fMs+x4wVQx/ocjAlF2xqx68rPM6JLJmdPdiaJAo+0casEuYMAn4up
H1Sg84nQfJBtkqKnuNVkDSBq9j0JnqttLMl7UKT/cQ6NFjTDDF9ca/99JH2qszXSg+Jr6UzQfXts
7snkT5LBvMwjlmgc5qTtzPZmUO0PsRh010BNPgbEXhpQGthdUEQ/JaumPYhtz8MWQvJxLRlqpMtg
fOJvr8T4ufmH1lk3PhZDyCoCaB32Nwa8w4xklXCaglATBWYSoyGwnuIfTZi3CbfXEwg4ykpBm0tI
8g9Ah88NmmsPGqDz4xirIG7N3Bpn6B6DBTmEQf+kQ2sY0HpoXR3jRnAEAUzIAVgc+XxIJiVEQuEA
tJ2NRiFrgLoHhrBjRCYBg8k4b+yeD1hqqPSKJUCaed55I2R4froDwMmzoqYumba6GSAhZNsggAJn
+y5E0/rySH+s2ITnA2ewNHLHU0PQ2C3humyczxUU9M28taAfIlWmU+KyoiPcAuE5jR/kurBCMWUD
WTxSOHZ/rgAhoKqMhy2LJ0kBD9+m2v8DdggYNw04e0yvZ8T1DHEanCqpACCOjZQFtDwyXPl1/mY7
Fe6U7LMFPwst8RvKrtITwnDDuGjpMm/8FIw+psKH0NH5zBPBeTDDVR2+rc/efvkCT1lTJGiqLn5J
iJhwE0mNMaZajEEtbb9A2+jwtqcLfnHt7w2wBrUcAkJ5hPe/m88F7kjr1nXZWei2ElicBbunIDt9
gEk6dIBiwpCVenjsRuOEFSDauQ3Dq7XlmJxKZQkpjggI6AmXkvcdcVwPA277oC7ERJ36FZyTITaN
QhLugWM4IZEjqkuezoXbflpseKfQsIZ9vGFMZw+xeiZuzRfOBeGfNFX2VnD7TOXGE/M5H2RmLhzR
eBo1NaZ3gkLB/pzF1y7Gs2ujBJFsRTS8WmVYIQ6XavGBovcgvgZpxZVLfANZ81Vf7ZcmAGsWwcZ4
FbpC4uqudMR1DJAP2V4Y0K3c/vI6TxF7QTBCWtw8tnpP7lSG6Kv1no7vR+j4Zcdrm8FULhADuptQ
mt74UKeLpxKxEGb7Ti/lf+uF0k2C2+NMHyW+GTdp3ARm89wgAON8+Ddc6UPsskAc8ysAGQtgzI/u
E/KEaWSCPG9omCSL0tpiUwTYjNEyTFTR4A2lIyahiK6LLcKa1yEDRxBIbGxVJ3yAyg++SphilT5/
R+2FaMh4Vb6JUBMh8WTbmAteaeEm6fAxyVS87uHb3IPyxGXjLGJluKok9y3CVcBut8kVgkxIiW2r
DdISQikA+HZSrjB59/BSJMPcjLoVAOmSvSH/+xHpzN2eVgyNj0m6u+CQa1QNO+vOVJFX/UbYtVyo
8h1T+BjI9rXhW6WRwNEByn5ltviqn9YJ68wzNge4o578WWV/XkROLCmiKHCT9guIMcd5M/WxoPzu
rT28d8z3owDvj2sRK69quz+MSJqTW53RRD3QK+VuNYS0IGSxxB1S10CkW0Zv73LO15o0JfQvEFgD
m8QOctEfIGj9GZ61s4ps1rRvJKZ4TY4WOPnehHW4/hmNuQz+ozq3+tIH5jSznbUg1CdTA3QRcc6p
VimWs+1UGk+6mtoIpziWfgkuNVnQOWYl3o6QGqZdk1tjb5oo8Rf6JE+sDQ5nymQGi8us5CyUMJsS
wRS5HY6j5JU/Za5WpzjOFohwSKT4gIJUK0g6RrvbhyrJgGQ70jRn1tF6nDl6L5rifbN2Quc/h+G8
a2eHD5PuPTNnBMUEU65hFOojThk62D0fgi1KjYznJNCRId8nOLZEO9vYCR0nzH/nyUnx5yRIoUV+
Njz42UCTkE/nwwBIyEcuxRScDlWPD+ZfrxXzp/Gb6NCFgsColhBm53+BUOR5wJunrQiVuG/uNwGT
mnVTcFX0C9BsjW14SkfcD4kImeyLM2bCXwyn9QNCYLg53xo3m7V4UdAlyQ3Is2KbvvlFfNHHCsjM
gfu4CYFeAjni/kReuMiPd+h7QOSVDxXWHNWFDhpQnDiBNvI7GZkysDpFylpI6B8JaKsTONa2VAuG
Lw5xM/BRrJCGWvD1N5y4yeTN3QwYx8bp3VCqGgdCXWVySM5TNNeXftq2I5psZ3QiDyYya0qj2aLn
s+9A0DWJo7DP2myX3K9pvmHpRX/M6YSRLzqBajo4XSmJYxb+eyDVZRcmKs8M/LlWCgleK8+E8WUA
ObXn//K0c4xAQDgLAFE9eNns352NGdWEwQ1R1l6wX3sXCmg2LG+HOhnuoTrjTsX/CnqSbf64TxDn
rIF71w8IFQhgfLV10puMGwn6aODmf8C8o2u9IMIRzBNRDqB8bt+T1qHsZHCM8f/0CXHp7mdYMqph
0k3c9JuRJt6sJlIMGn/hoyMytfiu2Ih5pLGlTx9Y9QyRRtsLhYVY8rHcxUFevFrPYdEumDntPrEQ
ksSj6iMuPRnIH0PQut57PAiOulBAo/Ft2bHSFZ9m+d7Kzs9ftyfyN4ymUZVcYwZgEksmeathx0SY
ToJ8VNJcvC4GP322q9YokVvkw4JEU+oifg2x9oTxkPHSmWO+EHeF/I09EEBp0+w6vX0NKdSIhqXJ
sobQNN4vAC3J72jeGCuJJC2T8/JWzoZNrHL2a0lg+LlV6Nz3raMVxpDaetPVrFdrkbOomCRcI/Dt
oLG9qvtpoqTOnl/CEURzHnvQGM8QqO/YgcjsLm9RoeCddzqpf9ZAYzAGlOvCHvwq4Q5zO96qTF/0
koa1cVt3kLma2qXPKc4+UJ96Ebox/2gsq2KWIdKkOsxFkMRM1C60wYFNCUYvJ9k9fctCh44nVPYF
RUIBqd5PnNLv2NhbNckeKd0lg3/uWaEVFzJGmVi/XWHhXAZb95FL29zMGzHlBo9bxlI93K/+QtQ4
D2yTwlQEDKefoQOn5MiNoNljDch2KVKv2KunAFhAfgxNHaD2fqC6hb8zIlvWpX4k1eAanPHNR0gq
W+g4X/fJKOCPe8iqJC2IsMn3BeFufZ0z+7uW9urSrGob0pFhjnDvsOHOjlQWfaID/3hSYL8vD2dC
adFDC72Xeqbkka2EJMCLvIVGXBw2JOFhtz0uQg9hz3AVzrhRMTZMudoLKkKS1aQBhTrxc0hspu2v
whNYHJcSQ3uzuQUhxaqvl1ZLvx1LYCjFSJW1MIwh1trgZiK9p99lfjzMR4ssdtluXPK0tmObMwjf
r8rCEPb6d4xQws3jgsAHbtNq3CHSo7QvbgnBErjedb4xHgcEnYTOXku0cK8XjUHLwtqGuBmfj2eS
TD6pWeYdP1v+Gqpo0P057qklXLhJAw8mtNGxMYTRN0IP4yj6i2KhsZNYy5pOWKfL6JFIfrjBqGUI
1H0hO6EeaxfMORzsGC3TBLlB21L32+q5+fOkmAVKTPf1/DEGAnd2mSiBmjIHAC50ErF4e8kWmS0D
rz7irefZK+nXzsnyQq/IFQ1fa9znKMvRB/tFJmFjtc6ZKzwCdCQ2R6DfavFbnsYnED32r4by75lG
LiwwEiHcT1LTEJmiymJw03xpwOnLNuwWfwHVwmTcVivKb5tlMSgYNI9F2F5Rgie6B0Fl9TdybmUE
sF7DuFQWGk8ygeRJUgZSXjtBii77dVQq06UWTjBOY0MqwZ4tFsT3+5zdWUJZ4q8sWBkoUNkc0TTO
r8COo3m+y7Y+5ABPpEmINJXh1tBQt2AcFbScKB07oLzSxt8VC5ZAPh3VmLjax6AGeal/fTqMUvn7
UHzHIRNvnVePp7ffjHioD9kNh0YojQF/KMnG+KHhKkc3u4j5mpQ7d1pxjIvaNq1YKsQjdORiklx3
ZStO0UL/tCfpjUpAgOAPIRqxqaofFrtqaVzUSkZ2QWkFVRLiPNIZU+Etn1WPI7KhSS18F3VYrvQV
6T/L4lG0MSoPoLk+gnnAAdz/uRApfOVpsSvQp+XfPEB94qLn8tNf33EbUEEukmciiVhtsesc6IQS
1+BPxelJRC/JAkAhbh1zWJCeSaytDOGuPuUb9ahC+++AzGesxYO6t2zHF6zcWtEAoKRbMjeIaxKD
bHetiV9WSb+O/0s638g7O1TMOv/b2TuKD0gjSW70Y4oUaWynbrTVbNtUsSKSrhXKODt4tuoQFCyI
/Xv8MUczyRd7wosUAaa+y2n8jxd2RsMLsF5XcV8hl8MKVfebGGcKXbaQh6ONVP37GPEUHArrH+D7
wqSDtxiBmVaxEZ4F2QrdLKOfnJor5ipJ2rmiveNmS678/oWlQKo2KrXhQY4cDglVM/mUJ2OAnaj+
o10ObcQifrw07x9ianup6PA4TwejSgFnpY70z4CGsWo+Phi9+6LMssx9AVbplWaMqLpp7Tl/wd/C
i4j2Evlpw4/fW0jywVt/CpVbPyru+1C5Ub+TQBh2Xc/IfLt2AjPimggrVw/RKhLH9A9USMzuDC2n
6I91xZEkIws+rVc3XJo+3nW9PVTq8mZTrrJf8Cylh/zMenAAB3XGAcPqx0ITo17tZqwCB2Mc5MvL
8MYjWY6OuHFt2XwS7f2TVnbpFjxvhN4m6o1ORTTXErcxAv9RNrHcV9JaykNfobaqOzyU2g3RbhkZ
KHjia4+R+7zfFyA1S1jKggu0ymwY4+iOSTumwXoijwQhbnIUdaJQ1n9StG4jGnTM7tqnR8zGVVdy
oHB6n9rPVIVlpvdLeMxcUVqAUC56Hb4pUDXHME+3jFSrXWtXLr9p/Cw68t+ww+edwOaDqiQ3haYj
cqm0ILkYg3RCwizpn6JNoWPEsow3d1+f9mFcrnq4/wgwS5yy++vdIW9TcWM3LIt2fSpMIhSeDcBz
E7QRcnbQ5DVr2nBui7YiqQCJwGTmyqkH8F7JWPv0D7awzJW5Gx8N2rEfDCKpM8tRdGZ1joQnpQTv
oVsUt/Sa723mepjbqSZZc2rmbwQKpAr5seaRWJu9E/fPRKCU7hCM9Eg4FDbi37OzcgUBvgMbxRyy
MEftuTC/gKVZ44A+N4zbkhkrA0rd7vcPDqkNx7jSnLSHeapfgMmUPjdIYDi3XPz/67Rep7TZnBje
9SiIiMcUsFkiNCVHW+Dv3FAnud9Xk5SeBowF4hg+c8whq2Kkz0nHrOa/9smlyMkPcXMi+rfNc41k
pq2ghtpWkqo2Sbbq4mLrZTLP2X0TsUOUJe3e5YpYGp84KtuhL01wmQ203cnXAvTvaCCj83VnuGef
K+BEz1o9L5Exzd/916uvsXoyJZgY9A1MNzztpnmkXqwd83uy3Y80xCXOAnMsJbIEZzAfacfdU9Yv
+hJ1fz9meaSUZgjroVSXxDdm5bp41qy+VADqVQYdcSU6o050AyMDBCjVjHRyLaRejrY+GxXPLnNq
fMymK8g0+XzJaQvbmeAR7CH+9Atg2Z2lQbs54dvh6bzDmmGg0lbCvR2nGAfXN4M100lhZ1mohUt0
+IacMdvB2SqgRTp4OsOJkxHBbmbu6kE/AQ4JSD4KWeKnkUlfhJlcMCSQf2TNfFeYYlBHFHr+UYqs
TYRrUJy0GTD60zUTk2lKsybJRsgqxCldU2/6izsfPazH51OluI5rNDIKRnBqL3u/9tRz3DmdCk1a
1dBmO/A9adBouXCwPq/mNPitXLw0N/IEBSA9gvLQHqSnjcS666MjbxsFYhR8yh0nPUzdp9O5nnBu
rY8NZqJ0dJRYDAue+xWensX5s3o6I3eK8aP4M4Jylqwq9ZeeusFMfemy1ruhMn+MVboj2fAclVc3
LGu4ZoYiEjNtIronMJ0qGdQO9gnueV+HVrd0PEO4dEI8+x+7mRdqVpfOauCxLCSKVxyCTjOQLjXE
9La7+LR3CI3Xj0PjklGYrH1qur+4/u8uGgUQT1W4AQBaAgoh1iOBzl3w+Rv/OTaRPM0Av6MR6ana
GdSFyD4nuu8uO0Hisuhxsy1Gi84azK5l0jm1wzYOXFeII3JBi4TNr2nCVVLOofltsMYxKs/RlCv9
rCtGOWgSbnHj6xho2sU+iJvFmkZQ86sjlfwsUbyyj5mU5UxxiBQ8WhvKG+CxfMY4pN85gNYL8dRT
N62Ijc4o7v3h92SVSRKIxfKdekQxHkxla+/5daXet0ehzsG54+ZHYRAUsI9YYH54Jcv/gus3evJ+
HHIPWgAUAAFrd+mvQDr/z6UqaWX4IW2Qv3GAMv5sOd7nNdu3rZD71S24XKnhpfkBq6TK/ikU6+zv
enyc9O5v5H+Pt1wfII2THhiYua3336RoXS5KzXRD8gqd/bkHlXW46FO1NwzHS5JJ/ZeMwSAiL2pP
Ovj20wyW3bL17cz1zVzh1cfcCVbRZ9fBFg1U3OjsCzvEQGZm+fx4B8himXvYA8VZFnDrG8eJEiBn
4Qn9CV0QozTacvukwv3IuCoF+TKuvMm0/ro32D2bNJjJSr68CvSHQvgXWiY1AmWvgoDZe3OJfGW1
IZNmN8aWtOTEVa3QyajCjvuXBq2KYR1L9XKJwZMr3mgK/XPVF5WpcOLo2hbSZnxIodYN1GzF0xSQ
oock/rtvM1cqSc2OQype6mGwyDDc6WLy4wiEXLfbAsCU7oEX4JbTQi6oF8SQtTOGs4a4bDpkaRGQ
DMDmjMDiEWHEGUdJ1myQSuO6AYRyNA5rZvYT/edNAnLTY8h3cGAfqdU6gFCDWy/9bXbGOExIs2rP
p7YZR//1AeiwfW2Unp5eUd4TU+v5qkLmy4h+lOURSGJEzhXPwWQAjkcD/hEKImCBkzQhhrbStyYr
aPZeATrkLnq8oQanlssS3TXBkrZokyoYjVnO16BevXK2BGAgLrvDKtS7jsuk3ToinnihhNgx1lM7
4SIl2YVSQZZeI3wM29WzaxS63RPoaTfa9eh4A0OpJnfGZIvYB8FBivqUIOdYlp+PKb4m9dNtM2eX
+jzd/aVhB9VtkoT5hUg/zyQ/HKEMATpRrK3Xy8T2kQC2T6WPPL7Hbt2FZJ4IhO7shhAp+Fp+bmKa
35aUPRcZr6xBANUnL3ABhFfr87cR4wLrYRIZ9QauxexriTIKfUq1t6rP5S/lggiA8lCvvas9Bx/m
fi2x8eNp+ZkWr4OVK08YiWytuqHBMObMl5ub/Ms3/x9j67c8OFOylakJuPtiYJinmGe3oBilGJqN
+eC4rt5iGEJ1yDpnMF5o3K6PTsJGR6yKkpUdlnYF4RLqjqS1oMlfbAJyP+XxGElZUczE9xBtQtEn
a9FYJsyS2uxF2oPJDvA4N02PzYo2XIhvQIs/hx6K1eemFYLebMAfwD7mOnTVblbByWyIOU2Kpe2X
JgWARSphx2h3SMjpY8SPyvWYF6KtZogkOsSwJmW+0FtM+YxTcCwpk2wpdq1IVGQ63Yh53aVoLS1W
f5OGGmTfZuA4JLPi2Z77pY/qsYJ6r6zOydtiojeJo2kTFsLKGwsIcaF0Qnejmyr1ffxBeh0szAUM
fv7bkKhZ+BWkwZZv0dHq5QxYNiy/jQxoH/oEONq+naiCwnasN5nddjVGxPRnyDJwnzsOwy0dfaFp
8l8jIYlbr1267XTZ+bvRLbk1Y2bq1ofOTyfLwZPvXPvvXFmhWNZHKzTDwNQYIoy6XTATzoDuHwNU
NZRVA4RmNQJ65KlE0oAmnK6srWT1hfXd3H9xOLooyVZVg0oi+xVVRAEVnedJof00S1p0XQuI125H
LuCRp7iEIfW64QjGLoPaAoZ9Nc2+rs6vyDGV9I4u6DQvnenlNKhGqa/F0ZQ6uoWBUxxlcLfz97lg
L5N/R6jep693Vcsb7FosNGG/9gnOCKeXg1RrxoSpqU1Y+GT+3dSWu4NgbxUncgmi3J3e25eQbkBb
WTaDNzbL7y+uwctMp3rlNVXDXjwxrDEJFOSpmpM8btNYS3kS32DPeBAqZfxlaoHl+R81hdn2RejV
41yzbC1Le2fSKp7I5AJxI0nxJKMOHUfEqyLU2U7vjB9Y0wIEbauXM7kgMKlHzSBW4ZoC68wIaSsk
VkRG8bzrVxW52IP1zJXp4p8sxvg/AU1Yh4lZznT+vb5BV107S8PLu/+N2x+G6I62V7g7daeen0pk
YI8BVOmOgqj+zLQ/4cYCyzH6oBMJkzmniaT8uMKEWGaS/2BMaOUjzTt+7N9lM7nLMcfPkLwfMeJb
AEkSvnmKpCwW69TlvXwdFvPXv7KnSF8TN7Xf6IO71W5fBbxRTyYGy2SAfRRBD/7IMfR4FrUNI5GO
0fE8CZWAlUgVYBRLT71E/mP5ByJLgH4d2OO1jgopRwqA32NROlCag1zmUPw4JP1/NwPrycZpiq0p
ucI6zP2vcZuE76tV6h2Pz9S6ouqtQH5NZKrveuEq5rKljLlAn5Q0pI/oeHio0ET98cqbJlIYVX0e
6r+c6q3ULSI48kOzvaxV30Bg5GF1sxXOAm/26sjcIbP4yTKZjG4AEsK1KFj4N+YTBk2phAKMNoSS
S0x/zFZy29ZPztEmTFT0GyekUnlQltJir2gos2574UkJSkbNHAzUhDvzs6HWXKnyE5KwELgF34p9
CLC+sQP5cXtji5wUw+56WZOo2S1cq7xZmdACu2egr3dpoMRPph0fHTWHtJaYBL0ewBc4W+9RvRB5
WJPOeEBdVfcY0icQK5No3Q3gSZvv0+E+Rr/SLi/qsazYTwHrPFzpEHG+UwwlNsLtcVE9I977JLdM
9SJhtQjrb/MUiiiXBRnypRYCKMB/3jtuTRSImglu6a3nv2FtcSLWAtnMqmR6ZEPGETX626fT61D/
vAnGvJJj2EKiZXvlsK9VUbp14SvD59+DKNGYmhjzPd656NM4wN53fsZczJzSHJSOu0FVcE78wCWy
On/RzeZ8ZdvwDxLJ0id9tGXHjajQ36rghYeB/jqzmf/x2azVG+fV81HSSv/8kR/8VfnrH3nkrfOz
QXjroI8pBb7g5m6TgiZV6bkTYWaEIFMnvf65lIcmpIJHcJ3K2a51B/QepVLMpD4bwEEpthfAIBjr
At6afYZj0B9CHQjBKiHx13rKQvZ92cCoGlDnGXl1ekoA0Yzfven+tv3q4B4vk+Y0eRazz2JU/8jJ
0rQpqtfDuwU/9DVCB9+sWqcMKsRzL4S3QEWiDFCMSGFSfMAXspPhXTYBxk/UdENFqNVcCfNX4Vz9
IUFP6hmsGZdNE8eHuZIctNfDXKKeO567l8BEg802PymiIUX29YM/VNxrH2U+1BUlrrzE/IuD2V9X
8YcYhHTpb3pHH8dy9v0qDV4a830TkdG7juaLr7oo7G/RrqQ2bYYYCxVDOfEUnbkAyCgEQntNCD2L
o6atdriDailAf0wsriLHvKSe3l84x5IT+ftpxOTejZo3UBm/2THM56p536CHobGnG1PTr2BprhrF
ahjRyekc44stCMmCq0hyOfsfLLXTX1pOOWSr9hEkys0uZIU0U78g6CubMJkmfRcrBdozeYLPXqrE
9kCxo8oYheS+FQcJBIDEnju0EkT9OpFyKkUVmjN/WregQdT+vuE7Q/C0miBR/blLR5rQ2x8JpGca
pm7LsC9yn/lHopBvHtiKrr9Bdt87judwNOHsakfWCdntSDBHzMNoAbILvf7GTsrb+KBFWLM7sW7c
ycCNdLq51Ru1k100vxvNLMKy5+wZJu0BGQ7fl3EdlUVN1omEJKAEUo4IRGFdSyYtkben8ugc2wBX
3x95lsrb5l1wWMKnFgEnV4v59Nnyk8GJMq1nlsAeC4ddPrfZc8VLtRkjhvoQRJPcQi1L3jwueCxr
A+iyIaBNcJh/mymK0UBr/LCjf2ozuBBmUGdKz0OpaLR+cbLwoiCoK67QV8dJ3iEYn7o5LKAbhhj9
I7LyMDaEWmLrN6r+66O2FEddL0PaNQByrshznZ6p/tbWzrDg9LpEqXopnmQWL30BYHULfFLLV0Av
7desMWlCPSahKtCjPGGNMhROqTvFNF1FbMeJIz9gig9jAEt0cJIRY4tb3Znrz+6Ibv6Z/MLLtUHs
PScbOHuH81iqYZdHdGNpCAclMIjRXq3ywADOJC12YjU93fJ17EAvYNI8uLiNRcP0gQ6d1ZSZiNif
GHMBkfRt+BNfsI3Gn+kLgwaSRAHmuY/Looh2L3u95V11uMCwTIbAU/0vzuy6kTWD/9cWEFz068Le
rvA5ho/D6yvs4OIbPcm3dWs/q7ReHXnKMEGudHxkm3tkA5twz5IjUejUhVcJqRIGim99QTZeofKo
8s8MGrIpUk9EkVb8JRWLmsk45kw8f9CcrUAlXvWxtsy3fsMHAS0uEYOU6aa7zfjwwD8L05I3Xr9p
RHRHSvzgtkElHhy7pdyRT0UFrWbOFbKDjouXlTpxMpOuLQDeYXoqBhH1/SHbCLKEc69pxkD71JBk
8NJzDWm/z92FMPE9XlfwsGAYlEvZ47dAhe6UF8MGYHirxqz3V6fqkFejFJdcWWaIHgbA5mAWMwFf
5AQ2L2H/vlwfHW7sz7VJAooSf4z+0rYhvNlz8vmrm+6fk6tsc39goAyq2NJHfgDjVBuuelZpY7u/
V6u1DTGyFzhF00j5zrOXGRLhKofeiG6LIsGTFXKaBCqYRHouCHWeDunlDOIXL3Cv++b9lqTHItkN
9CDP0S7BHUx+ZoW4RzeBz6kj7ycIzG82YllHVWWYlB8/GwjSz+Termezo0Q+/yn1bmxdOcOS59f2
RyrO6WNhzVxdGAGmxMxHTKRlBO1PF9t5mLUbsOSxf2IbLSPrb4iLlEYrvYcmF9XOTSD4I63fzcV0
ry5m/hitvswwwYL71tMb952YFqBpgMpMorD5U2c3rDMJcr7k1JkTo5jrW6BNOXOUIOB+xJ3XWtQy
apAin2LpWnfp42wwMmj15hHL5uQbpBWH5/FNBHi0F9f2UzXAHhEBxUnm4WAVguqw6WKuHfdgTJrv
6a2dHxemk+Uv1KjRUStGQq5xJwgbWLsGJjACCUXScQKXCGdfuGrKF7jSaIS0kzloaAB+K0Rav0VK
AkaFO1h9Bfqqi2iUK8ZSRtWA4/wKpMoR1YpvxrkqfE/DqCzZgF5Ue3lvV0Ei3oBHegKVAGjFt8V/
HSUhPTeUAsvxkCtJ7NL+er8S0zB9/e0TfCITW5gEdqmsqGlHSQ0YrcmdbelbaCBjl4reL8mfKWHg
OWVveBa6YU7NAzrrd2SAi+oIOanvTYVOoOupZj6VUWl5LhmiCLc+dKCSnvuLNHBPBE0WzUSa9BCU
JYOQ64Fc7ipUe5O5VVCJHWHlyjob3Oq0AKiZoqWCZ2W4Hq7Op9XXtWrNRbVpGhAXWYAKDREbEfvw
gxZdGeLoNCL4AVGlPD7p+qre3NduuzDeUctDDJ9mvFGKlYWmvYa/lYabU56TVVjZTpEgOrg/zQeb
joChzf0ZRmUIrc+7SyDxi1GLeXHZkb0IRsOcP7YVBPrd5fNJ+jzb/uCikvNTi2h8F/a9EXCEYDs3
DA+ZVUBaG3MXmuTyPpuIF7/Rac/xI+AmrRJFAYXh2zUkCwQbGzMZyi9IG9qJw1OYih7CPKnX9/sw
v+7xrVjiI8qL7PRjTKccu4H1o73rnrF0aJ+looGO4SUzxZaFEj/2vZfWcgvdWebb66xfsNi2PYOy
Jx4rARVZ6HOlSpif0uwGDys3oEIpNrCbSGiHkk9TRL3RseK60ni8MOh7z0mQxFk4dUUJyQsonLsS
VRhZqUdqi0S7RMfpJOfZNf8V0lQc6NBpxHDywHjrdHdzN0iovXKHCCTWyxDKudcQqIevolOoYa6a
Ym5iQS2aPKGiD1sQDM4ezy2AQmQLSQB/My2ryagu/Qmx4wNkzPfmM3jeVuiOYAfvA5gpOSQsI0BP
j1Oxlse5TLrq/4LKVp7R7B/lqXKsSf5n1xcqQDkQSDxshi7MKY8fc48hLNqNiLztxWinjDkjnEok
ppmw68c3zyfBt98CUyKLaiK1vVzs9sktvZ97k+1wgZ2QQ9uzDQKGLrYd2pwtHuKhQqQTyU//UxFN
37uR+SqlKIa5iLAwx+ggxm22w1XwEejxREeNsBLfNHlNYsbOzjiz4+qPk6DFJD12oDugFmjqDG/S
tNqeUKNOgS248PnedX57YYteS5f5VoKB3m2r6BOkKEnqZhCIaBn3xpE5FycDxO5nLbPjfmItCbkn
9Fo6rkE5Nz18Ke2Twu/ERW5oWLgGPo+XB8VCrCJioMik8nmA2SXpy/+4bm4WVD/spMCHQYzL2YeD
iA89JS2v2oN3+l6BxSer7RUSOtPdyDdwemmi3a2jdGjfObHWE0xH5eZYGuMnEMz0ifH8fKW45Y64
cg57aDlbWbyzMSqoBU5jYG01Eb9vbqQmVtDKhTCGGyblYK3/sqxmk50QV8bmiz7hpwznuhjX5eGS
53VycrLmfNx41DFN13LCSbtcK1VnhiBD122q7eb+MybWev0y0mJpOMU+bahemq2Vce3dkSlJTUpp
RVdvoL/rSmp8YcFQyqVQ2EjXHxk3pBEMMQgnX0QEZ3d95AJ4WnASCn1GD6LQmaRUFzQT/LTZXHt4
2VlFE32U6kXwNLHjMP3aLXawt1MeKI4slWyXJmMa6ZmbYnuUeg3S9a0ko43LI2Bqr9Tf3jKeGPoP
qMDY+ZvvwtVGJplAAS3plzQwZStNCaBEpHvic7E+gl2I0Y08wRNhrV+G+cNHt3zF52htaXe8ghvy
SbXqMvsogENN+CVrM+3Qtrlf8gG+SKhr8P0VANpBl/4txdKgDfm+N/ytKjEBsXB2xaUx7uPvULa4
I82G1mmsnBC6D/1ZyTwv7tuLofa1/vHOwB7DslmAbghUtzmGfQJSwSJLtn4KULrYn+EH4oca/ty6
1AH+iRPO1qHDF7IpLcUtf0nwI2FYyi8VlBTNjKSJlmbwx78oJNNwxfSjaaEgGq4u0un6PeLt++Kd
otA8cmWuShP52DpiwWKfWT6hd1krPNGiDhgV1B4P2rYCJzt/XuGTESZDIfijW6nttspp9cRYuO/O
6hY/BrMXBKyx8oJnU4GAUzoEI3hRxvJl6+yiVE5RYsfy+o8sNSz0L4ozKhGySoCL3AWp+MMJMd2i
e/v+d3tJ1hIWY/aFndtKScWKAjVeMr1rc6vxM9pGNJs/57OxVMWvHFVWr6bvDQXzYqQfNYUuoiAq
UTeXnrp81yfCgTjrX+Orw4wygSFQCYYjiWGs7Dme5eo1F1g66ztKzJ5LpPzLDkn0jQGAinrB2aV7
m5Nhzli3y4EwT1tmifDYYHL6YZskm2wd7PGNIiYWOMUvqUX7VpVDoI7UVCh0Cl4pk0e15o0c3Njc
PPD33FmT5cyxxNa/8myPhs0ONWV/8VOl/4So2NpspnbAgdG6FVSdcTB/duc7yDHbYtQ/ulQmMUrY
HdDjTd5gfmHN+1gVI130FOVWPIzvxruxb2Duwu/5XoojX8+LmgLIgoWxELvP2Snfxk49MWFUm1LL
VEXISSqw7yP0g/owmupq9pQjhQFmVC659BA/I4dlUEg1BvCB7iFIufsVkzzsRl/VlWdgd8CqiV5N
Bef5UmWw+sowbcqAAT4xX/i1vEOcZtcHuxBN65AusceEcavMHxLtcYOH+UduXNKj98PNQ5N6SQIa
xjjYaOwyk0yeAkaRDGL/voHQIlJroDvI9MQHsDaUi3UB5v4aGvW/NzLOTH8CDb68r7okaRqB93uN
pj1+ir93tsRr5Eo8iQGX/F8/zyEQwBOq/SQK3PAa0WkHxHifATYwGb8sYTwwEREl4ZXJwtPIVCIB
2g9sB/5bmcF+jhqkWAlDbM0IE255ToLHYPE/hKu4yZajZyEQhlgl7EPfyNLX5LPJXB5ua7B+4TaN
ZN0J6Htdfc6la7tVlHjpbQXm54qusODSG86ynzbzhfFtpCHkmqKhsNzTl+YY6JQ3g5DsHj2wjfG0
s7fQBR7Ug6v0yCYKdL90kvQJRZ5jA6Q2bwtnIlI40qEMMRE0qbkK2bQ4+DqyASvUgsNX8LHxJAm0
roZLHj493xh2x9W6DGJ/bkidg/ZssVWc4RtquxwjrQR01Z16RSnnlQLYC5sV1NnOJ/74VgNLmx1C
sPvuC4zEg2zXrHoT9KtJWe9WfMSiRsW/7H4MR+ISDQjiXVtUJPFRpwWxkLhUwNzr3XxOuTc3fGZy
odPEKcvnA0csBD/dVGX5tZBpTtsLeS8ojZLdtdOrx+p+LQmnUeZtL1817uBRruzYuE8nrqlx1+aL
rBJzVBG8aMH21lAELbSQeyB7/P8xO7Pluq4MDDUuCY84d3bvngATH2i054EcS+vrrfqcKE58QTXP
wYfMl4VueS7DBftZpFto/v64v4Caz6iDuUKHjA/3qtZ7ZPw+QqlZqNnscdm1RPnZSIj2rqcq/uqk
xIYlCJZBdtzVyeB2IDnLNWcW5Ei1V4SuWyICcLO40IaWKzPnFSY+hNaO20djz8EfPlz8O9kn3g91
H69SV2nj0G8A2pDux/P+7W+c72jz0GWmE0aeuWnwxw+wVQ73tarWzcrhtXB1P+zmk4lV4aIQXD66
o4zXvaYNXPI1i5emXcG0Y72XRkT/9jwsZ8cM5jbC9pVoOkMItEZ+QpwP51gb7fmYZ4quXX2p3r3h
9MycwK1s1UygZFRBtx+MOcQZtIqrBbe8nJikba8ePZXuKXEH3X+TQNC53VZRH4wfIia9gCnZGyVH
nm+9MuUmYrJ3XP5wnxni5q4UM3B41wO8QFZf1NAbiVmaawbl1oMaqJAtC5WbjuyU52IxIne7tMtu
gfjOQe/gl2horQXWvgaOSQBr+JShqkALw/H9C1/5Pc5wlbHO5S8vwZCMG38BgGzz7SJjR/x+02UN
zSwNUC7TQD1ADHViyAslNTnJVuD512BHpLbuL2QYimSu02HFHTbt1hQfCjz2U40mFEZuW4s9g+bi
fH7VFlpa//Tt/y+XcWP+o8wJlcecb9xhJly7h5NOaiciAHwf6MrlxUBaV7TucQQ1Wj5iI4SS7ThL
iXNb4ZnPIxox3A86jF9dTAlzEMZKhlgXJqUEwwGco5q88+ybjpBcvHotWFLG9F5F62fgxwk+Q5fP
tpcQCL9oThuERC2+P2SxIRnto1oaaSzVePEUTdjuCbgvUTtsBCPb3dfAGB+bchkHRkQodjp6D44j
hZswDCbHiOBvS7QQLBo/s9aEJHUc05YQnY+jeSgBkQFAzxRIPeAqLy4H02kFVsOUPTw/+QkfKswE
dB0gxPDGLt0XSsdfj86ihZj2SPLWMXnkrfZXGl//1Gllt3Emjlk4xw6AaQpVBRz2b5pEzjwYzZ8E
hDfqTa/n66k3Egkch2cxEEIy7z+51376wpwuulmMfjCDG0iMxvl+6WZ7Hl2TX6S4wCv/TarEwrFB
+u/Xr7IHyYZDwsEqso5xl2RMUJ7T09LXG7pFXhIN0U/eobfKQtlHnL3HtDtCH3VWynl7Ikllgmku
BPSZ0PHzpbfhZmYLru9JUpl9JdUp/zTelYHYvr0MDyaQIGS1mGVirXLWKdrT0wqSGMhDYGNG53ja
m6q0ayt0fPJtVB9sWIqfI9+B8LHkaZjv/gH2i8nDQgBxHz3FsaRn6zmEizb2aUndZuFUjpBHYNA5
wjpQhu9Sd9gRlt3inlCyPyktZdDXuaFlpoO3fi4DIL/weCd+EP0bYITTpPayYKqKuoY2C9BM+kgr
TEJbUWfm8RKqctVmlOOrVbXWTgMUoHY+WWnDi0GM7gcBppmsSKtBG6bxoyOK1yHab6cxXqSL6kzK
m5keHvt/uHWH5mjF0Enx/gJ2JAsjyaWHf5mfxWB287GVkP0DdHUBhmAAM2m6jQECtl4Dck6O0cQ+
MetgrXx1lh7ZllOJDz1YN6nqJ8bpu2ykJJ3xeRgnH24e5VzmyBODeBBGsDsEWq06H50gZI4TL1WI
4vVlPPjTR3n3DwiirGq4ZFEZr6E4Qv28ltKAZDPAFq9sBoYbRzwJA26Ro9kb5ZSbRIt2hoO0CaF9
JbkperdDbHKkx67L9gxWC+VbuKk0SXsEXy2Dw0R+A8vHZTS0iF4yk2NpYCqkYCLCM86zooPk83D0
M1IbaxGdcFMIDrs1WoOAQ+Ai/ojfIVBNDiorh52NFx0RMUyJHA3/ZgyhQ5dagLsiE2a3JYMlbI1o
+oh2P8TNFubiw7Xszd7b3xqSZtWEtPoRIFLCcB4zvqW8zjAfqneYAqbyr0SVF1xLyUYVh0RKpCjY
aMFi5xGAAVhh/SOJ19BqxvUD7P7dZEWvms6jmWFYIdvES7wjBw0h+afUV2gYdViA5HjaErZTHRlP
cq+aidUFF1rDVEjz50PGifsO/0CUwGNu8hlp9OL1AZeRW7tkOOIY70ubbxKpDuhR5hfw0FFEnBkz
ChMUM/kk/Cd9dV6Ftwoh0PuOvve5RDhMoYT4OereqvEyfiuf97N3XiKaBbq/4FsqJ/FmyWOIJl4b
c8xnqbncXPc0oVZ4JCBfotfF/Ww08Tv08EHQc3fMO2WlmpEFj42DvM251tzyFbJNujZckx+vQ7S+
59Ur4bGSDVB1gHDc1PU02f6zyNTpJXtOeV1aQmZxmBTPZjlUmtRQul/YHGJADcdDLd9onTkF5Cau
O5I92EKobWCx71+gM2yVzI6i5/dUCZc0pQBIRKvHaFrQWm52SeYnSjyroPp2jDxEB+3dLxXM1Y77
2LoUUJAxnjckpoWvjukoP22sEfMsr2Ge2opkCPvy12XbU5MdG9QysBHnbTtUm6Rh0ksHLAcMBp0h
pyGzHx3N4+7H4EjQu1t0nIWfs9LNAP2NLUi4DYP4qjh57Dr8KHyj+10BQOzXW4IzlzbTAB1vGZpR
wblbtvmSMdbUF+vhWbgfWM8ghrKepy4DHZ4DiWLILdTUecGPvu7G0gWVJATPhotmqjZuA8yJlL7b
gRv+LfSsd4lweIjalfAkJ7vdZU4AlGCZiUJFQEoZ6B73a9dJTlasZsbId9oMoEoPKcSpYnq6rgrZ
5V6Nqi4CEZYD0aWwec60WCbkN86dpuSG1toFAOTqHMkSysiaX2h53rEXRTk5YugNaKl0kvJjuUCE
bu/forzI9Vwzx5k++g4Uuxpz9K0WR5Qr18gF0ycn7kqihGup/+Okl3VNSmd2GROh6/P3sSCIyOfA
eBgKYY5mKK95a9YDy5N2/Dh8yRa2o5ZjymCZDtN7k/8SEpYMTqdURK79S3nfKKRDppiJvw3h79Am
RwJhiWTjzviGcvlqR4xXUGfOk0qdEarSagE8qqECCxValOozDZEaTjZk0TxCsmIMOaRtEst9NViV
j073je8d24auuqRZbnKYoLTvHtT5c5DiO48JlBieZD9oLjqosa8Wpjp3wXkSxa0Uu24wyDxESsN2
6mEwVFtYFIKBxQ0z0VN0Twf0cF132M56MElO1dfa6DhMmKoq23A36VHHChCBVuV+Bi+XDsPB0PYw
cieIMI66e0CD5P0jFFi7mvfXIbA+Fs2FvmJ/vWYkmtX7UB0p6WDpjjqQVxtS3hqu09Ur12sXRuiH
oMAV5sJouyfqX6eErUQfbrA7B26/E58AjvzhYs4V/S/ENyOJrsilvOa6q9bOhCBDJM4CKfFP4ilO
bN1xJW0L+6TVw7PxnTMDmuoIXP2IdG7t5p5+VapFBjsa1toUuwS5AEQP/McVdSwRigdKj3KYwhkf
k6iq4eDR+ezARcNKbQum/EElNJGZunVgzWgR2j3vudLDjpg7yczsiVnS3ejV9qTQX77P82kUtc5w
7v9jOo0dhHWQlEWoOg/Gmu2zRH/mEhfM38HIrsexAWO6gG6CggbdpNj+r1qQOvkvrir9d29eq+hu
iOXTt5bz/7jf43v18VNw6oYplCSMPhRom1YUMdwKsWhqxUmx9/QVwBmfnCYi8O1yDD5bd4Y1kpUe
xIXb7YmkcDY/iUv2vzOtBPGuj2BGmUCNRSBjBT/p3wzVLVx31yq8xXBfZytJHdcYrTnrw+u967QP
QTZ/EISvgEDXKWZPrFsflkKiQGIWM11dPYsdMvbsYO9kFqh/xI+Sn6l8PDXhWKPGGFGmApLbqX7H
kaj/VQlLum5F+2YiN8ARK9H0yOLtc2A1ryfqJQJuhVY6zRmiAtN4j6Tkh8t/S6IGaS8PiFUSj0mC
sHIVh3BYKeOF8/iEHDv/6WD4dFRTiSUtZyOrYe/4pmK+Y5fbqKZsbYmXGqm4/L1Z2jebVVaHdOxX
/j4MQLUA5tOLoIytvcQFqCjNgDcdhhE3H1OeUJav55vsrgKHrwWBUWO+O3gci+ZyVDB+3b65Mc5t
44cQQTzvxhlwfdvgRMx3ZXZc7zF0o4C5NzAZKC5CJP0fvU5H+21s6bgoH9aZ3L1u3adBdL9uHChf
VTC6ndJtA+Zrv3bDtInfA+kRzZGKA2ePXjJeMMDntjQupDPQ/cPej5Zk96EjMXD3VgmRg5s5rmqb
ebnLmr/CAEiYZWb20m5lsthABiVQ5ZqzezXYkREdiH+SWywHMQqdaEerWc9AuGZmGDB4BlgkLieQ
RJvW9s9LFTzpj3r+jp+2XijFujD3doEKwCXlIE4I8uS01XYsI4arhhy57GkMyv20FOZOSDnL8emm
BiMsOeG84nCQFzs4p4AkeqR7y7u7XVThUENnuy1cUynNEM7LCanACFinFLNB3NKkGEx84jZJOFL6
gA35IhBt+qdThkaxR34v3C06xSvsWEnVnAB5cDBTW73cPAnwGZA2Ytl1gbo8MNl4AvGMACx4eZiQ
ZTReBqvBChhyEZAaPi3UUI1zwtM7Yqh6Ch5KllhcP5g3Py5Iwa5AArEO0yQgtWXHhKf2owA6YsHn
V7hzoRLLUVwD/RuuvbyYm6HRmbUIvrOHQPSoAjwsLMasybIgKpbTDqbXpOgLaRL5hOo9nbfEvxpt
q0Apujp9UAjSGPM4OuQH38YBQnqplgTpcUP3s0L/rUT47PiLSqoLaccR/XvDv+V9R263Li8tq3gC
m5wQMNGf8XnFaxUtYLenFm3iJdYbullXmTcaHqSZtaaMndCzK3q381P/fNdDZxP792IQNor3HAtD
Eiw4cy1CXpkGWhST6aYUbMcRD311v1OXxxvC4TW7F8LIU3S/zoEqVyKVoGts7QHSUMDXiC4RWF8o
zunnAOQOE1ZCbYS3oH6VbaSVLvHFZfVMGShmEjUejxYjAzCWdIEQ1HbelZb4HIpB/GEpCRLvKS7J
sQSAZ4T5rO9IA7G2j53H0Hxon+AhJrRAX/4oTupNTvh9OpLxA0JZmbh6F1MVIPi/AutiReiK+Mlg
zZxPbMklzZC59OhrL40L9feHpN2ZMlNjlN/BQywMLOi5ryLgR9kEv0IY67Encmb7oG0KDlmxjds7
gJaRgN0/pMH0UWwWs0pQgLeXHbazW25CkFmyRIfB60oxkjBld2sa6yQTbkA380LGdYDRxrAY1fN9
OeB+m8SLyvzmqDPJr3MbgHvvGbTQxfTJ854ryWjQwHx0u/14Bu4pYq6LwVP+yche5bowmWqAms2k
8Hk3DJfTJyUAAxK2X2+XS536RaSx4YO389OAUW9j42pcg7FkGAmbKpMWkUfeMQb6Aft+N8D2w2pv
L4h+g4ZseT4O8Ws2myUm8S50FBSAdXWrf8LNX+GbUXodw5aJB8E1Ipe5ms9ClubBBRorOORF4BaX
aSSD8uQeX9RsXlI+8v+QfVbscyUvWUUHTgDwYDG2yvQmo27eitzncoGaTjRwBYkv3Cz6cBfL5h4c
Xop2oTbAuaIwu8MJa9ML1ZMaYlWMNAHiZwDSsSk6OWNdWwgWK0d9Jxs0oEE74nfXI60ygcwpVUh6
jI6mwxM2f3rTx6d8VLDjZvq64AVexHWliW1oJ1C+zqjmFvwr67q2987cdZaSAXbL50j/N8qav6+F
FaGv07zfUkcoardtAstaOji6qaHEYVTTySaWTVpWsieE5HDj/JSwoPndwT6alV5t0alkcYDozmis
yiCcYHBII1WV0c9u1nL2L5yRo5egX+N2d4hvprGXJzT+Ea2diQnbi0X5MszDIjwEm/GV9PaDVNfN
j5j1nrDX57Tsl4jZ47IkGTJIpuAfcVB6o+GnvMyN2roGARJOzyYT6dS57VUbOpj3ApYBKfYJwQ9j
kUarTQ24Mdcn4ZvAg2rdQyGXbDNvBwibwxdJqTnC6ZACWwnXZW8PyXdn5i3Q+jEVT7SKfBclw4Wm
Jjv3/gvC+UgwOTnJHagjFHJvqOTIwxy2TCceDUG7pTSp80M74P71rY871MkqXukVrx5hv9lvqz5w
qLMYGudj3cPVUg7gKBklp2M8eYqTD+Xz1XC59c9FW+lcT8JVkD25sJgrLqZgGufvFruYkneHbae4
nGzxQKoxTJsUG1DujH6EaI01V7PiUDWveFcF/AKUmMCdVdZY2+6NG+Q8Is2RThVodF9yejUk8+OE
4QL5U0i2XtlNdmkPlSAahDkr5tnAfns3pAMaroo+HdqYyZ/MZhXuYpXsovfRqnxnQciaJU+KwtFx
CaYKozzYZtawrhK18+C+zKxY7RsVRq2d/iQl0RWAofvHQTyhuQ8w/oEochtBoW5OUMlLuMfBoieR
obEr8Uu2jn83D0QeelPSKBRX4ftNaU+cvCEdmLeHePxwhfF0hzr2XOlbw8YtHRIZNSM6IwPfIf/k
WIaDrV9o5YGHDNaq3Z+MfVAMcS5vYvuJY6dTKI4AKpHP3L/dDYL/hOITO5A3IATsD5M3QchyiQeA
LE2rCQoHEsdEYlalDlJt0j/gNvOVRHDYiXRDI955o1V0uWFcgcznx5WM68/VyEJzAqM3B8RaeCDi
ZVFINdK7nHSasWQQ+wJnqWuI3jcuv5APl0HFpGtPdD35556egIFXoMZU5UGRaABH+qiqYPa3dmNs
HNpYrGBF61v6qmkN+47b/Yb06s0RWo5Mtuh20V5vyma3167scu1p3nbIEFEwvkoz0u3Rpg/t7HFx
DHWPU4nlM9NllIN/slgFUKH3+3iCtFL9OmyaRov9jDJ4Mj+cf2O+7bP7aFI2Kwj0X8SrtkIu8bBu
2DpLgV7dGNh65E3H0fWewG6ihBZbt9xWuiwApmXu1NAMezEVsPiAeWCYw3c2T9Az9XMAgFhI3lmY
8IAn7mL3NE1tq9ToYV5yGpFr9Jx3LWf4N0FSH4dA48H18NofTlzuRcW5zH0cztQAEtYBsGGyKUjT
hQ9D4ehcv8wDeAYtTmuIIKqvyi1HS5r67Y8e+vY5ioOiTSrMVKmW4+dU8pbhcc5aKzrfI3O3CWJ8
mmejMA7O1RgFCuG5DoyDBv0qf4TfpAv2Q8V5w96T6cYQWz2uqftm0+wVCC79aKa0EqahWbqlTPP5
fUMCBNMBYRvS7/C+E1yFnr4KOsHdklG6DRRFj5i8qx3ANZ4Vtk8ViMmIwPfXhckSGYo7ltxflXTD
Rt7i2d5MxjNrfWzZlji0T/8y9cZOa9mfELnMJzeNI6Z26tSEKHOkd/pQP9J2L6Lv6+huIvFLU8ty
oNowAsb8t6CluygeP46nhCyjUKnzOKqP+8vyUnUgsJCJzyQ5v0Sw4zRXRDjW/8n1NgAvivbFcvh6
yKLH73b8ImnOgRWhGZVOGcMiHf5J323KVJQP5PaINWK980PUWohl1JF4dOmS14rD7xfKP8fo8fUF
9gH1u5mIR4vG2fEJiW5i1y7D6XqaA5jFkIyr8+8H5CySpunumXAT6PJF7XLjvzMA+Shf0W+l8Lh+
utY/sQ6HixcmkEhM0SSZ/Y3NTBaa66QAGtoCZ1Qy+61QueRo4/CL09SLPD9Q2GA6KcmOg7G1s6VM
9JM9Mcpwl87aLHSacVaYvjIycqRA5OGTFMWZmQcjp1WVIZ+Y7cGEFekYkZZ5yD36u8Cx5mz3y/Zj
uYOQSek3eST0kaAU8Y67JoTpxx4VXy2b3CgO/WeFaDWJSwfwA7HqPRH19pjqolcu/AzbYchWuorg
3fRjs4JP2fDOJzRyed3sFDsVrwrE1laGlxmP4Ar+oGQCtaud2ixFVN/P7kMFpqreJjvBM0O6GBgl
qnwChym7m9mJGLMiyKtZkpA9gxcYIiZy2RyGokEzJzOQGSrHl3TGddI+BEeTL++FkRP3TX3TzcDi
2ax0RDVg2RUoOZV6kHeMzBPWZhPbItrwbmrEPuLSg4IiA9Z9K9xSugOvb+EHCbDTMzsK+maN2X9A
WtBKEyKRbQys4rS+LtKWPq119JlPPEn8fy3w2/O9mckV8C6UZDmf8gkb/tDILMj8EFKv+PrYAds4
tYkikqleFl6bvESCBUjCgJewwh6P6ZrWtjZjk55vcb8Mfuvtnwo/xhByRPkGl2UZRvxWHaH/8/5d
QDstI4sSVgOz3Uoetc5WMxNzvUNrt2hTq1b7tn/rNy/3WaCx/JDX00TBcz0L3xtlsNgPshZY8clC
oxIZG2TE1Y4acz6LuNU9IzgTsE72ipa8/cctVIkbBpBxufbcOZBR2SvHvIMGJbfrXFbQY5qfoXc2
1M4fv74oglXnvk65ILDCsGTzYlnfGDHmvODGTK3HAUj83/vIyCgds7LYtuGxkCGbJaL3VO3y3kUT
1qlqwQsX/IWYyJ3bpNuKBgd2LnzvSTeJ7KOfgv3MPs5DA/s5BLkLKpjYsBsQ9MFfCW7mYiBa8t77
0ai4ZRjANWVA7mRwpFrdHTPLRWZT9zzxJJFJg3nr2u7Q9zLTBPM1MxTMSfcp8M26YdEOcGvGeB8B
6NdzQrxMZv0dz4/XjGDID0vKJBkLrhjEsDevqVEIiBv768MdiR9vj5NF3HADeZDRc9hH02yZDzjQ
d14SgpBtnjACGpgA7C09gcYqhSvNspB9Bzlf/Nh0LGXMgXfW2mBhiHBCs+0vxi2x1SJXMaR7+shh
IpSEZl8QoTRYI1qOf8KGaxKz0daE+ZVakM64LQwrCYjiRK3MVGqNkDY4D3V+VfbL51lrPcbyvIvm
mjPcYcUlWpBsoX/d3CDpfvx4JYILc1evLmgzw887o5tsdX205EghMmADLGav5IcUMcOkaPTVVRck
hSi7MqAfZIuN9ql5fde11eJ3kuXbYCHdyPDcWo4CgUE8EbJ119Fa8x2ffmyrdUasKw/fEb3lvnD2
5r38aHurV1s5peGLr28YuNsycJhFIb+QU3W1HBboho0oCGiJnlpDzk3RtuqPH6r5ICUQf1mPpKeK
qjtwQw9XebhuFdfj8Byf6m601VWNaV4f1s7R5ePvp+2hVFAohHGcE/cGwsKYU6BTCD5JNZjWRube
ka2CE3SzMzT1042oYbPCozN01zDkOKDAAf4ynlHunX+oF74d5GFWdcFkBC3C/i498hLCpSrefpRR
/kbRPOds5inFSby0x6XAYBeX+ZZYHpZKlqv8o0gRTX+jOeC1E3g2vBV4nV8/1GKSI2LZ0bQXA8Om
w4Y0zvLKaFjenNVwSgpdOxYvwLJaBiAL7w7wqztGSxJo+EfP7dlNT+lB4p6FoV5F8YASxpGX1FTL
Occ6y3LM6y7H9jYbeAEVKdpEzVL1ZkdtXlZkNpCxsQeJRDGfelO8c500gp8kEmn/Lz0ip+qI22Fo
tmMq7sek9I3TujUg8HQxelkII1+Q1mY6RC2Fa/vYNL6y/j8MykGkA6tknhewK2QcYbSrq3XfG9br
mWwtl+/XVYpl1hIgOIXwRA6UpAdVPqJtPnfYdibeOjKwlvmC2u6CNz7b2S0TjUCmaUSSJDbA4ut4
PU0msiSC58yRiJJE9JSvx4Uwtp/6lPYMdavxKpwqDxL8uZhS8vntSjcWBHp/RKH03BjRTt+yPcJr
0h4E0FneMYg54TDYkJCG5RypLwLBhiZXK26PXefl8vJ+LprKgMFPD7X9ktMfniWWsetDXSiT5ASu
NXly22AWRNbj7cSvKb4Z6v0uuZq3KytdHVXYAyewKKjm4gvG6nAbnytNeQHM+wzAZmimpFB8Q6VX
TSoVT7IlTFSaJ5vS/TN4e3l4XLND0ttUMXKmpkzCxZdDJ0Wwl7jtxtwwA3xbpKbgDn+uoU9SxKf1
iovN+fx98QUFU3EUw1wht9chOuvVhDOoYf5HV7v1QZjXPIiOSshxiM9dhjvpl8SxLQBZ6m1cvg+w
rjaSjd51HHYSSuBmXg7qxEeUnODoOKMdRNdwXc3BtKLb5LY8e9u7mEdvJwqkNFVe2OAToITM9ADt
9M7T3OuxcehAJUxhXIa57Pw3d/T9CtLoeK8yhEraqcSdjax6lqYqJEZIjbU3RtzWUuSdBvufblR8
OiDh2SuWg/FqjCq98o4mTQLOeFIkOo+tp6xeGEqVZgUE6iSzc65dzB1u6isvz8tt6a8wu6uP8KEw
UeIELYa1LvWlxZeuS/eCKoCSysKMg6ta1rfiUpJgsXgSHuW/wbhVQ2ALG6pnhfhTE2CXpbIGWnDw
74VS5qTZzSyGVP0rOEw3QB4cRWUOOcGydCWu/JqhZY3rl2O31yArodVSlz/TBPd7LKC7PKn+HAkU
LeduZka2jXloaIX/3j9zVqXS0kEXIMG6eWxM/3wIhGLHzvdJoNT5lV2NPZSTWqFs+bFM8eYC17+6
xpupGdyk/DAKUiuQurb+M64lfKg3QHQo0ovIVWuOQnI7XeXy+1wy+rGjBRepQ5omTsOdFl8OdQnA
h3XBP1jCcIGBKJ6SF4X3wZhx8RvRmrdTAndDiPg3DouHlTdmXScKYyeTrUQA9EM9GpEB8o7fddOj
8M+L+U9pPe1+2LduYaySKWYNzE42GGo4GpxRxBiyztWh9LCXYTsx+F5MRws2b4uzLLqoQkL2MUvG
t2Sm0aWq5nCv7lbJ/hOG12m13prpA19gjK6I01SFJM8lpyKfcFb9rtne4H+YY1pACxV9/oNp5T8s
rRCxdxNezd/gmTbfLhvDEGVrlONs+vGA5lS/RjpRycK9MMnAuh/D2A3YHeYVpAbh1na3XTgz6nSp
eSS+5mO5yD6j5UOxehT16AEtfdewpMMaEAah2hE0NiZcwk1R8X8XsFoRU8JC7j2pdg6EbOXvJCk3
nUEGFr762o8afdqGe9fJUKsB5LjdabQChfwKYDi8feerF8volp6toSmYHjPEx1nypwmozxbJF6Wd
/Wp9UIsclPRpH36MFnMlKAXXTE7xLBUCzP8kWdZb48ImzPzEN+TAFwq/npztDSdtMobju9aJM+RB
loXsaD2ArcvIdzVezZGzxPzwqGzPl+EqCdcQXpGgA+ZboKL1NPUI/510W8xDpQ8h12VMdjhC6AKi
pc2cyYJ/G3qkL+fLx+L7HuvSaXrPjXynSItcg0qMXRESg4eg818wrseWJohYfJDLhz0S3lknizg5
Gjhg1EzflpPa5CRiX9S6g3hvgFAGn7InLL9KGqTEjs/EF1nE0PGQyRBMNC0jIRUw+YmyJi4Dt2sA
43eGvJtqcXAt63xBNkIkd0OKZ570fBJiv2J1eMx2GJgwLZNf4FC1cCTxKdN+jzb34vzSLM+3p0va
9qLy/Qjl4tMHx5elAHQu0gVanfgB0th3sy3k1WppKRQ3HFLdQld/dant3u3ZyT6yBKJiExEzYhwP
xIYqt5R/hcZbeF866a/Q5HMBCKRPWPS7MtDzJCzDsbVVpA268vDO2MQ6nbV7eL5LgbyMEC8mLaPl
TE9532sl7ZNUQPP2SikLqugJta5YAB9HOWaqICmtEfqXryOJ78HPGYjd0jSq7YE60xQgWmAvzBg/
+8rYVp+caQGbVE8PwO6ye187b8gTXX+E0b3G8KlNeXxBAPAmJfF6s9Mt/nzKw8wSEZY2gsET9IWa
9+ogHFLmEGpMtFcdXsmdbLVJJTo+Zfj16jEwlv4nREF4Tu+Pq4tuxsXZcWgPuDd5memXDXehAEbT
QmFoMxito+R/CiaxdJAFf5rlkWxqbnfHNw3Dr+Gjb6QUlHMU8ljKryJLSn9uPyb5Q8abZ40QIoc2
uG+Vnjwvny4SXMM7GMDXDOyWmoWDs9WN43FRuRkgPDvNS6cTjPsridZ1NUJo58lmA8AZIf5rrQMX
xcfaKQPtcpo0hRG0PGMmVexqgN67E/QVQzVCLS0UXiFKdTb2ewM8mSBEMqv1pn22oDq5w7F/MTYp
k5GqH1s5Ld7ZCy8STMXXGvWJs2Q6kUT+C4lxWkFaca4jJlWPoJP/2/fjLIl3PgKToAne3gpwNHRA
KA2DC/K2EEIqvn1BWdOZUjISPXNuq/el9DcENuIvcJL87vE4iRwk02tmYG2KHB0XMVuijXW4FY3c
w7NU11D0Fm0Cgg2jhUf1Vo2FK3V7IKjzP5ry+bOc1LciwFvEJroGstznPyrRGYmqX2ef/8iM9goP
vRTHEds6f98dcOpLWMH0QKS2eFeijcTrB2uz7WcSjh5ii4SVpQ4wscCRbjJlXMAAzI4yXwIuUHIv
ecIayF8dZTo4X6tn2IvBqJlgmjSVvBlU9P73F2P4yXP6gmA254sEgWh8coZo6WY9TJhhWX1CF3Ar
ayUWaUMhSrBUI1KfSAgySSblLZ4KxUE5cYPZ/GduBtFv5VKvPxuFuPt8D2FoGCyaNqOg4g5EeALH
ur8ORGMo0AH1kbpb+SRS3KPVVkB4ylzBTNBKLt6DpuTYYrYIs9VGO/GOLQHWLFgPBYr7mJALc5cG
UFw5QxTk2BGBusKw9+SrZ5b++duxs9mGHmmtE7mIDuSFU4VSEbj9bR6qXlJH/6BDo6MA/38HZkzz
ZbK3Rqk65kGisIHOpCRmPhuetqdSthD+iXttTFTwqM7AzF8sH3Ox7Jho+7UoTthsfso8jDaUx0MD
Ro5xoDJtmrfouRQuh30kQ9T50JXEpuVHcjnKmoYJcxmcNyAAfeX2SaDHnOjTE/bl0aZPVeGXmfBr
ygvB4vDl7SVUgDRwKyVRDiBzk9d/LwruzrZhAwj0VmTY1Tax4wbLegDBrFLqNSfsGWATVF848Xd7
3uhkVzPKw/SH7GO7QLaeWI7Y5i6RAyPcPVU54VPLdXrzTw5KARTg+uYyu/vbdo1N4SrmSvOCZKkp
yxdqV29ROPkvp6YVPJgJdtVGiRcY0qvq4j6oTj0gXOOO4Waj/D5UJklXnFoXrfzHD2s+oeXGr0Us
s/uvlzPsFoP0j3/bD1aGqCEudLjXP7xNqN8ot4Ndt0QISzQ45vuDHXMWAC7zogbZ77gXvoDdkYpy
eqMmeCJlfi9rb8+bpVExJxnWPedCD0mcsT/jFW3rvfjDtqIZBujVWHAjgPDDytl0z1mQyMvY1eqH
u7Is0ZVm+yQloGofj5O5dsq4dhPzMOY8BIoZIyHCk+KGRTNuyraoWlEmgQ3IlhHDIw8BExDzw+o3
7OvCwelK/36JSKoJSSkONvIG/87+1HZrkpCn6MsdS9bQaTBgnjLjKpDPeW8tG1SBLRTb7MEHA3Zw
6qPdPjvLRNL+/6heMuy0qCJj8RsvJML7FJoEUbaQuFn2hQ6lMRvCzmciQ54VQ7ceDGYXrFaZB/rH
oi/5UchmyCaHR9jPiaOZ+ZgSmphhHI24XFtbWvwkz8v5SMTl1wx2SuyDYHCyyMO4s0B60I0M60gn
9LxmyCDrG3dLuI5Z7N+ajuKbLsEGUf6ybtsRStj1ugLUsZMjZtuN6WeG/Dag7dB33u7J8Vdd/lOQ
nsLkeTBYCzFTJ9NK8njEkvUjPCZgAMuYziYhwr7/bEhwr//xvw1KGcBhuVIcYwiQID0zJG/wcMS8
q3iRQ7iW7VC+s3+jAN8nih3jprau/4S05hTXYqv1tmFGOlqm+Dhzb4CSlGmEnay74c3EsiSBBNYp
i64mXNjcamdAxLlQql059STgveqL+4YRBSXM5UNHATRn8G+b1HK8vlqIWyQRP409i3PHXBXxY5q8
fFa5LShxPTyqqRhUJ4mq05Pu3S/gSr8R+yJOXKqv88TUoua7sDPwfR8WEuEnUmlStzJOfGNGx+jO
KS2EIT5vEgXlzwB5mtVsMcfjAcgxfnogkMVpApVc3mg04CcCvFEAhwUzdO3gjwtlPutaQtLJ5g01
F0FE/N+YjGChv7wTDqf1/D+GdgugsaA/cRAMtQe+/ISgas6d9JehtwZ+LQa8EQfRy7SyXs+zTOOH
4qUUeEf6tOw3aHFmWejyr26QSk2sOEs2rjD6RdI7OZWDexw8/S0G3I3Fez4tNCvY1uXlOjfWjcrj
AKhpntvWlNE3G6bEIZ2Lr5CDRFTTWgkf2RfKOLQ8SAlr1Op/mT3Rg61ZrkX19ZFoof4LX6t9cN0W
M6uAyYMRr83ApnK//a2fO1pb19wjy1XbUz/OVIP5GZpUm+Lcw7SS/fnxHcX+Dg831MCSF6KP+lHJ
9A8o7JgGg577JleT9m4FRJU7VavFAM7sRHBaD5gEEvF62gfKNzMp3lcu71Ew4SKHJL6OOswu+mdZ
uaZ6Wq406nwykrduy8FD6hfMXrBKhafi2rKvzmA/7zMcMUE88VZdCRPrgezn3ZjED4DbbQxfDd1M
Hua+u04E99+8ZIJKh9Q2VgeoMG3uqN5F98biRijZ/3Ogi6yyRDz9iHj4qUcs2NyDAuIdbxRY4L0K
xSmSYFolBc/M/QKRKYNoSkxVzM6fZb5yn/mPBrxP80btWP9312uchtR9uL24dk6j1pUDaW1F/kVL
lS9v2Urkt3ri6Xu0Fudte1CkmdAgvzB7XdGR8Uz25/7x4hSu4pYoRFgh54vXt1wV/852+3yHe1Ot
0N5T+LCtbtbCOfFbDlKuihD0cD+y5pOtZ4bEBDljZZtIkBCf/gEhWKiKlTdF8wuvLDpQPnswHa5+
gv2Aa/+nqy29n3Ut7L8LR2X/x00UOzeXEbaPgYd1c64aJ3YNl7aA4/Lc7iv3n1UsGmGKLwvJjCQf
2cgVlJyYdt3jw0bti0ZF7J+RbJj3YOdCvjJC3rT+nQTcwcJVuzk1ue2aV8UQl4vnoHi2XBAlEaSP
SMVFGlXLMNTua6/pj8prphPy7hwrV1nECXTiHYmZaNxahK3ohBPBVsPvrEHDFhM0uvcvn1YKU2HG
1OfrcwZSpuA7LjeN1GN0YQZlET7DcUPjHJwusc5Ywqiifrt75Q+5BNMuDCXqCvsoja8GJb9zQNQk
U15N9ZsajJNLrYykRCIPaC767quF+nGDkYr3ikmBIsnzhj5B/JZ9OzvKwVOvNqgHPMcoYWKdVGbY
35XQjq2ltqMR7iKrNiw5j51uOuGAapeA1i5vXGOX5RAClkJVfTkMmG+XMeG/b5uYILj6EUQHpoWQ
3sfyc6J6rvoAC4cK/KsS74ud1Us96aD/bXRP1Vt5hiDxF7ygMDJT1J3JyEhpM/3YaXM9Bi7n0gBZ
cjR2bP8HWyadcQsf+cun8x1mYS23N8EtSunYzCM+h+ryZ28AcGuf/V72yt1ui//NWPLyKINhOLcX
kuL3yI1lJrYjbP1heFWwYUv07uI+fKKda4fN9qvCGd78aqR/zjpgX7qWgU2nR2g5raQ89n9HOSn/
+dCq9dYv+EU51nqvJRYEg0b0vNUn0e172QM8aBH75fN2NYiUjboS4Ba5wrJHAAJP2GlemTxUvAyu
WPUfQ300GOgWAJw7QCrDRnNbhGylhE2dQcCUCLcH4Iak8PMbdVkzv4Z60TAG3Yw6HISyiVsIjJDo
HX/weaGMcauGqBEQk4duqqBIY3eOo6+WgeYxa+b5Tz+ZOpW20I/FbyKmb1nx6NXw5fyL40Q6JBpi
7JdoCQvxmINGVPZLFoNfURA33gMOafMJdyoKPLTOZ6+lI2wHrVqM8/7lSFtaO62heQ1bHiA3sulX
eTqOXxqafe0Kep5mG3U7TLVgl4etijuuJcITxjKb8W7cv1tSbO1wCgEP+bAJ9halXdO67EKhLUlZ
IrIyMbYdhrLGy38APa0p1wyuA6ac+m7HcFOfC8JHnMSYrocDfkRn0l986EI7KH/U5Aa7InDolE+O
CpmvMcuUWqIzw723JsIuZ7cZeywTHscW9GB0ldvnyq+JQ5a3ivH/un/H2lrlRhAtvw9X1xV2n262
44+0V8wdOIX1zfhokb46OVRN6aDGTjlJhQbXQIYiReJoi1deP9i0BbKUJSc8P4Gdwku30PI9BDWX
aDaecl1TdvGxkzXGWkq33TH6sWUJiH/K0PehtQe58Y0FAELrXq24ttAIucs0C+8gyWYF8NvdDDHO
yZDTXpuwR/Cv0TjFqgEUaUUq14Hh03q65bPDzSijS+byC6pz36TT0J2wlWoJ6kbJCq7y2U/sidJD
NmweFHrTWjMY7BpjkWdIGPL+/3P5dH2y09OwS1yDQrpW5SmKu+1AlgHaK2lontRyXWvzu5Il+DHh
mV+ar/dSaoawg4tSbL7BlqXv93b9qJ+veZo0qvtzzVRMRnXOb9CEyGjqneven6Mxvurr+geYFNsg
VE0AGQpV6sfe0Jm0PIYPBzoy+ObQaz/LZesS6yUwgur1URBCHgOa38jLjpNbCQHOlUeueDh0o8A5
8DLAumk36lm+d8gER4EMRemBO4T/fbDCILyuN7T4+ypalAAKIA1wZIcvqDrZXBPO7xg1+CDAyfRC
bfTPFmTs5nqifVIHWHzpCW0ps2RipSx4TCZzJwuoN0euTZnGMkATD/Lyx3fW8wZeWdQ+ntBrCkP4
MhboYEzNn5AEVDPUekTQeEZmfQKFCGEUOauh3uEzCG4Dv/Kb9/UrJWSrTRQ/26qwkKiyWyKSpHh0
AqmALdmlsQpw6OrtMlNbtOCL2cbRPmySEcqH3luM0z/Q/dZR6w2i1lmh1r8VnF3azbYRozD3mUXq
pA5t0CubO9lHZTHXvDL1LZcyfA2M84t2jCjY1Ks+iVOLujcWOzn5pcHXUD2jPflHdUv22swan8uP
66nECvEV+eIv1q7YjB9LlxQFMXJLuOPb5EVDCFo1QI1bsoXnXdliREMm3wIaajYZ/BKlUt5VvmZq
XVkrsJrCnsOeIxf7bfkO8iwcJ9Iv/Wx0cCvCo0xzr4ls4zfDaj5iEI6fiOjCD7/hva2ajNypeXC9
Nl+2E5Wa3cGwjwdnFWN0p6HuqlDC5Oa5kYfup9m/ndwDQd+0t/gaXyaftaLhfJ2Qu4T3myNNLDeQ
/W8c1cSQzWYSpm40CK53+f29QRq6y6FbCka9g3/tSdSCTXJAkT5g7oK6df/z6sE4BiZ29XGeu3hz
mtO75BzTTj6sR0hpsQz48pFxFtrXUtJWh9zJx45dg0xn42uAz+oj0/Y+Pgy1LJzb86JeIGE70GAM
0YEhr79yMyqC2gM37PZIOKi+4DFvpiGLStQ1RsYKEku2ovticOSawVlei3P/tRm4xHmJt1OLvKuN
tRQ4JBDtmX+d3jFkKyfGyimutMa/CI1jVFAfI0eRr4Jh4XYJyjJ6EcXxea+5UqxZBcyIWCS+xUxw
Qc5IohuU55Cee0Zi30LAmbYLUAyKrbQGIfqCssHaad2N/ZCIe6zC7y88vVqo1274YZciT2LwFXQr
dKLNLrwXDQzoLuIhe7tQXUo9hgJ46a54UnjoHJJOcqioOw2dwg6KrSOvtWdEW+QkgoSQKG2kSvbx
shNDO2xVVFB0/ctzyxn1GWmzCwbvn+/m4unVrpYh0ne5MY3ElDWxsxfa4wDulaBVywg5vrJPb/qz
7/nT8muydk1AkK78XuGxUUBm+dizDwAMvsmmHYycac3u2UbDXLXMj/b9l743GLOChwsqQyXgoTTd
Tc9H4lUYjp8i0cVbAKTRr1V6YcryXCCodvzAohnBtabZwuYd4KWzjKY2EeooJybHhLv7sMPK4OY1
BOtNm7gpXblykugmx0rJqGcPB+91fvf1zS0cewFwa5ddg6qqYHtvhHNY9y1p2/ECAK0wafrCQl1k
Y7wGHmKbzwKI3RA31e99NPKLanOmWHn6wdxrBM31H+DYr6HKHhWElrT3B7paDSkQbiPu5uCmAKX5
yw1GfzoQBotB8k0dJycOifGnYvLlz6dev5phs+Ihxbnzj+E4eeUstFziMWcntQPDfnvGkPeOQZUP
RbxqkI+ntrKD6OWNpuPWOmnzZtHO3rgcdp5Nbiy90rOPBg1mhmwFDLDsJGx2226la3Hc34S8txG9
r2Hk2nkcUZKEoX7AWpoX/adbAd9/edhjG9qBm2X5DVQWthQqYPhzwMd285NTceMfJIa9Zr/phMlW
B6cQqsO1ODfYztnE23AaDEiXsSDBrv7g5uVEg3VNIxBAMTTxqkUB1enWzTB9i7jcvEPhzBcFikZ1
M8N2+/4vCaD1mrseOXd6K2COAN6TkBDQcWjI1Tr+2fqcvzDnkOdZHQxCgmzPcRQKKKW4wayX3BYj
as3fR5moM9kf2ztkiKc87ZPjgsYgd8T4tAOap/qdbiFNoO3J1B58MJl38jqpPnqdlcuL1spSpwLJ
TAOx9QMXPJ6rakXUJCnAxRpE7sSZZVpRo6+lu1hMDU1X3YC/Jm0v1OAMCaN68b5KF62M6oLbp4vj
BZq7FQjCDwcR8zjwKQuRyUXlLRSbUWbugUH/Evv+JqGPK4LLMbIu1y4/uA2cb/EYiKq3h+6zlbuf
ZHcn39ESTZpjP21vmF2r/+dXyFzpnkTWS8cMbCvtWCJ0upO+aBQUMHbYWW0okIDfUlOR8XhWrIfa
qkUZABKsnBnN6kY/XMGjTvWqieIiXe03o1Us5gk2Id0LNRT1fwOeYRyQDcyxxJWHl0A+Uk4Agylx
55QDQS/+Irx6N2/+jJqHdRRf9+TBeA+WbXlDCPEwWDfDHhH6oIS2fHkDjsL742KvbmQLK0du2hGA
ccy66+k1O6HkRnQR/dUxg+3lUPwd4z6XQtuQzfeaH1bKyKjomJ+ZN0Kgm+gdJmF3QJa57/gAmH7J
sMZKrMgSO9h34t17s20+eiFwUjEMVtUdf83QzNl/eXROTAgd9TmjbOICY5S70uG2gII7L9+um+rD
i3t9KP7UPba3nuFfNABVS6hAqhdyqlpDysvJnJrMew/FAsPXIRcuihOeVi6R5Pp2BXB81u7Og//3
Ym125T6jFWKWTBzoGB3NeIUoVjA3Ej3FIrhFA2EDiIrT71QQy/XPSjGjmaGtjM7KGBflzaTCs5UU
cpYqAhnNWAXEo1EyD/++QNS3jRWv8Nq7kHyGR9QHb6EFHA9uXoVxdeBGYf4NRdhMOql97OrYuDNH
hHBozsrYvhjsLITgqcKMkTDaRRC2RcviVEO5EhSM5V1UY6QMErTLYtzDiKaPYRD0RUcTP09huNUR
W42BHTl9O2pxPBSFKaxI7CWcqCQ6SEatNM8cd0sWJn3SOzOpX3KIqhPZFzmdZde0bh0dU3S8XNws
++bbYMwCJ83S68gX0MvrnfGm3fKvdLT+FQrA+yDQChzblK4Nzjo1yREPansVdZ7PfLFRRlxTuWAp
NYXKjHq5bP1k1ERQWiEdFmNGlLL8g2XPQP2eqo3TNoi1oiLBoeiN/D3KgMKLEYzL2Vw7wyhFZ/F7
vqJMXEOoIgqHPEcFl95xWF5VVQohDeGMRxul27zAwvstpcKN8kEOMw0ysh4ZysYpW2pPh3bscW/0
neVGONTPr4Es6Yuk3UrK18FLTrDFuM8cWUQgIolXiT9xBRGfdtaCp/ZrVXBG2IxUCkBZHp9+Iaw2
XbjLgYni6PsgScREiEoFKE06PAIStyjM579jJBGzBRhdnmQ3hrMuFPfWczxHmEWlzE6swvGIeblx
2NvUcC8bU174akFRcuDB77sDDLCuMQ/TXqG6fv3LZkld90LjWqza8LkilwnSE9EABnfqjFUtzc+T
jAn1ViooQjVaRbe7NJ5dI4uzovOv9UndOo7SAB8CkM+MhyZh2IM9nH15rtXzqC1T0CSfdbWcr95/
MgKrJ2OVJ7v27YlQgDpvIj7YaxrAxy3Alcr5wKbVWLUuQBJ7gcAYCrzJkwbbfNM2zsCXXnUIsneK
Cgbs4sbEWbwnyResqN0mA9Qr/rscnJ9CCaGZq/NNE5FkP9p+hqqKYPkrb3FirhMFyOg2X/3zPkyo
vtEWLYNFjV16pajuLm9QXyBfbbhByvOQ14amU+G9Z9xYUi+o4av3ejz0XJ5NB5iicHY0OUlnhMUC
uStaS2CwHoHwzg9IgjBGPiJ1T1oMah1c67GHhkWpBg1DJ+eaW9LwAmc0E9Fn029moxuvSniw7Imv
ewjsVUd6l0laa9gTgrKSjF9Sqa8vYcsXI/kfDCGRrUSMh6Aa7tIjK/tj4xzqBJOyFUJQK68zwYzy
34+awyiCwPGayGFgyjNIN6bK5Cx2XuvNqLikQbsMjPxczdIImlPrO/jfqVIrX7Dg3mhXbwv4A4Qq
sLc+/9IhlXiS+kI2N3uI526yefIJpF51cTv/G7aYcMCwLwSPi4OV+EwObEQftPmCZrOszkVqLIKG
67O0jtYvfK0ir8mu+P2T/Q+32kMPF7QipMt3cDh95iX3qjkTKdvCwYU89X2NBVZkUYTBHwYEM+Qf
IkdAWZhr9o0Yi8v5Ul1/cWOv5xk0O1/55vGq3bhhhpNoYcqEsSZPVlw0tEhJlkDSmiu1sgPQaoAC
uKz5Qz9tcArl9mNA9vHliWiOAp9DKtgoZduByqT9iiFYMoHZeBmp9QnVJM7xYAMcp/0s7vtTLTl+
yHL4v9ssn1Q286rgM38gNMiMybo4H6FOgj3l4kR54iuVT3njQ00W6x9LlnGxyWRbVNMY8emayjBM
3DvEd29q3KeqvfVtx/a+DsfWGLu6BFQC7gjQ2xNA8PO7/Kz3/xzld93sK7XtaDGZ+O5BxjBFtYYp
UkDWMnwT4At2eVMxiMYSQx6HkhFF24ghwFIwVkySPfXeEOab04bmdO3v8BXry7RWwo0PXlVe3my/
UG9l33keEDUVukwy/tH/bwj1QvM/N4vO5k13zSbu0a4FZwWCELrf7vxkc30p9V7PHBQuioruWk8H
+pZUN0LcofBGw8LlFMFFEg96v3GhIXgROViqoYN81A9T7zktjn4Ncl+dSJOsSVf7YXprcpa33g2A
8sK6rc7rPJztHFl3W2QnFG5P/5mW0c5YTgo0zylKnJexysXMdf4OJBOd8K1lvDXVoWk4MKUg9pMj
ZMIgCQZW7tuC79Jijjfpi+/t1slx3x+s+RcB1dzlUzfRU4JuaW8rzqAxLDCJZP1pIK/UD831R4A0
uNAqSERi61pPOumxXRnk4Go8tg74Zc2+/i7m66B+R2N0omRYvTddqNuPexsOZf5ePwbkN3I/jt7H
RlFBeIoqxrPHHDOwbiR10+efTkWFb9PjB7spFmprenHZzrKRAQEp2qZX8qqq52EvkqfnivmS03C5
8SY/XjpNnCf6UaUqVhiC7fKuP4zi8U0h8cAYDbfYJQgvPfUQIVEq/k8BtWVJggo8/+c398ZJkwBh
d8BJ95C7ld+xcuaHCSforrUj0ZHQ3IkJSnGoDbLO1cb13jZiG53yq5uK7JG/HLvtrsmz8eJHb3W/
TyiNK7arb6ma4JjEKGGbp/7+ghqy3AARvYbGjMyDFigrdnoY6fSB6dMgdonJYSrGEKpNAgz9xey0
4E0+B9L3taYvf+mktAEQOrGEc2RSZGXWmBWGG5Dc7Zb3gTOqgvM2xIxXI56gRcqCU6ziT+1qRxQw
4lY9lPPuqGI8Dokkx0z/jYx0UE9/dhw9A1NLqf/0qEp2Pjt1erPmCtol7kfzSPifmoVrIhTB9wUt
nmzNHuE6RGSetLIl1neFlhFNxILHEXdh2MJDQBisdLPwq21BO2Vv4E0TGhOrEV7SU6wq2HJLQspd
oc/0qAmmErIxzTDiC2kJvX202stqrHEaAkmTYTO/8NNNP27BT3n1fhxStrP9ZYJcNoL39uypRGby
V7dxCSoxJVPo5wV2isdK8c+soYWAWbuzvAHswLhjVnNYx2mALww8vo6LXduDhwZPM5+z7x8kkHfZ
0BSYQjsAIwDfWJphinMroI98wEjltwZ+xIGNhOOUvLu86KFimaiIU5UcpJCJFB00w9BjUxsObHQI
bDAkA2hHYrD2Z1CXp2QrV4/RCWoIDUJ5fOrYjs5Y/GpzoAoyZL5E4jy5vQouCjQPHNoJPF2vP9Ko
g23D2KLds5s+ngowtK8ULSnEZqrrfpo251KH2gPGee0hGTJeyqdXULHrWU8d5jpNaCzufZWNoOje
IdHs7fDYvIhmr4p330e7soa3kf1tK276dWq+TXIa1RwmIPE3WTHjyfh9rb9nWTqbc7G0x7f0fUOd
h5AtTkpaXDoXGxM9uuUliTjqiizsZA9raaehicvNBObCrWexACmjoAbZkJnpyTM55hVAi2cUpt8H
uSuB45Dow2JNgd6mRFkFnNM9RDGx1v1phG5ahIBdi9KP0hi+oloQx4jDV9fzZZoTlhvsJ/pEeWu5
Q+CAc/0fFqsB1SuZxPCCtt3TwBuLfT+A1tVp1QBGoyenPbLyui0mJjOYRdCxm/SY/8FVH2F8md7Z
P+fQih7L3zUhM400JOmW53BYx4nrTM52WVRXrIR3gT5SaFnxvfJpwDEaRGKu4qxyvgtWQzaEgIhu
0NSAr5CtacZB7oF+StzrhRTAZzK0zSpnjFGdTeNewfFwNT7l9QuMtkrB1i2rsQv1Ie8ecjyoaoMJ
rE6KRBbT0Vf4rxx2c83gheBa8n5MQv1utQra5mTaBdnzw7m8jFALIqHUcO/38L80Vqy16fB+7vdj
mcqjaSj38RWBO1J2HaNt2erRZLdl2RMr7NTMQWBVJkYcNN/++qrJ0cXcBKhvIaYoRj0uj+acKil/
QP3pUyRm5MDVBRYyUs6AcY0zCbuhxj8jXg/d19bjkkxz2ZR/U/jh7BTnA9NGoVtr9zszM/kzhK5u
uFNYMiOzo/gjwLYjUdyn30TX7JCmHeASbxVmp4GummgAzKmPTM+DLfRhgrae4KCYrjUVcYndaK9z
n9r2ALPa8XlM6Qc2qKm3BDqvI+YQPnBRDeJaB1E1sMs0aREi0Uiw8JrvKEq3IzcrW3E6FgP8Ux7T
BDdAUxOYyPg2fhBxOjQuBsOh4u6SuMfN+NxwDivFxe5w4PYgSUtpath9evLUCC02kVEOZXD97kuh
YCt0Gyy8L8oVY1B3bn+ewIPkexFlBxzqISxKOPYZyEDZKDSY/S+aKdNU+VFiCbrkG1NbjFSYzHEN
xqkG6hWSHgSbR5i0zuzWg4R4BVypVlXjc6aG7e6rIEm/4oSS8yq4FAfPuizyxctjOhINXlBoR8he
oGNbPYDSlR7QpvTJ0UTNkmMWeZ8z8e1Y+qJPWScaLbfjQeRZcXcJf8Vs0+QmC/q2BZYfxrbBWqpX
vPXQ92W/oHE0ktcqZf1FL16nv+hmFhk8rodQqumEFmMJYxT0EtdwpNFfdS7ST1s9tsyNC4kfSYHG
iPOL3SAWpAf6a4qoA/32HXHk/f13F+Hqt7A4nZuao0a54gZ5A/3GQqYb4ReAH94biFTLr3RN85ZE
ffe1oakPwYU0LwKFVHrC3oPj3hMkHwSeVD7nfkcFoP4hWt8+/sxw3kr3FeNjrgU40QmnM+fv6rrJ
/exI1c28fGDcsfcqdtxRNNc4rxX5cD+YLRir+nAGnENYwX6r3wEJRhcNgumqm39Z8c6uI1QUEBqJ
mk5CKBRYaKcYqqDDIuXsSR4OlVxCRIyCuzyzH8a7924SyvGiMAG5YOPSOcIU6rSDnTbATTbLXtdg
/RgElewgpWjo3SNOL/twmpK3PAU2Hya8Odjt0kQxjGc+Dy51DG2lnCLdQIhG/z9vGMegKlyDDgWp
YZ+fPUcOjaaxwKII8nxEvmKvrAOeBPOzdomSkmCg+dGDoV8X5gPgZDj4L8xTfUC6vuMq10nwX1Vp
UBIkiV846OCa8S9szBnR6u+9CzRNKWqVbf8CT270waLcQ8FLwqqdxjXyx+47ChKs5c+V5u8u5oO8
AunGTCXbPhYMWF5b5fiPcV5cDnpfhyjCRtHJEEmyNY4naDEfavapIjKncudDeR6kYB6vUbocqAzV
tsHLCZpSRnlq9oiC85U+klydZzOag+0azKj0aT+/WcCmB2tS1WKdBSYa4cP9oVXwjbaUagZQFZcj
l+lP1OHMw4iWQsNrsC2hS+f1BfnyufZj917KOedJQQx2YebD20N2PIxq9FowY3flhXAFe6A9Jute
7eAfGxtAMRIEu8EKCdfxFg7QwN9Eg3yXa7WdGW4/vjtX3eFMuONdO6JaVqWz7ahsDxSTPw1p4hTh
gHFrD0WTvtR1H977UtckfPtg7yBhvTH2980js862XcJte7jENVIXYezU3kuw+WyHOpoQlIBjjzl/
cV+jFeYA9FOwPIiLcvJ6zfXxG6u7nhdzBhGrs/IGQZiLrvoZi0z8GmvG6zZxVCxUbSHwNGGOw0jT
vUC5M86IE8qqobL1lvSASsQgdyJAIjSTX7aUY3oyExXzfA8mKjfFRL50Os3suI8Hbb2RnGrYy4y9
3TlJeskxDqKzp+WZO7qbZCNY3GsllxUFT34O30N9QqO5hkGD3+KS1CtKuVr4Tv3E9L2SDCCXllVg
yr18BPHEHT4SUJOoHKsvE5TlLhcooaXJG2qDjKexw0Oz+vpx0nR090xDmILvKYMv7A080/wgdaxg
g2y0YY+36VSYo7lqYa+iUtizG78MQAJsZhA43fooBCTJxQzehVSG3+c/GkBXIa2wPQIpUt4AOvYu
qf9sqMMOFJyYLbTuo9ZuTm5eJqD94LWguOo5wulIk+rVjQS1df0aMebTItETO7STDa8kuuINB4K9
Me5pCH09YtydzKVlNwikLoDpiBjTauytKDtLaOKQ2p0hTEa1KuByRtuJHxgvYMDm/d5hRHDIOjB7
Q80+Xsh1iBKJfhO5O9kyxiCsf6Gx7oEtAHJlsYXuD52fygAAFeluTKtMp/gpUOARkXchNRVmbQHM
uVFWPjBvzP2QmCqUcRgDFGp2hjv6EsruKm91o2SjZlSaOzERor3Oe8PTS+6cG9/Sd+3KX0oC1uN+
VQFiA0bdnjW2ugriX6RLkGVoKW61AzTl2g2X6+nWB/UtMwAtzgrr4m4mGAMlPmakRp+6IJyT+Xiq
DUSUQ70C4NEAYmPysDoAD5f7KgZaXE/tTpEpQkzO+CV2cTKGGNIeubwn6iFU5dc4a0hPnKZE6wA5
axmsokX1HAwVwCScmSjxgfeD6bsnbj2L+0pweB7d+IW/ufsM4A0ZRwi7UnpdMEzqpzWuAoasDxMo
iHtcltpnv+HF10Yh/YNiWwnMqJgME90SqwTQGkCJAxFBK35lcPwD9Ys+q23LeoXFjspG+wSMPmri
W3LQu+C4+uhvToVb5TrQE8ov1SR1oybTqlxU9gRMoEIY0Od+1gBiFXaiWvnl6hUxeXI6GWLRK0cf
Rx/GpHyChu4zBJ2LazYPgvuQffflveDjxCvkCa7pCxgyvm7P4FU9/k/g1uDwsPtLzSw/zXI6NMU7
x4F8AUMljk2v86fp72WnoC5/aJJ/CvQnQ7TGm4aXtvpl7FwSsB31WxU80vAhhDqIV/DECLEUpqnf
dt1nuLsDkTxPlTPmQM2DhdJtQ8Kwx5p83nr+gh6QnwrGqY+a8oKHW2Shu+DEN9acoj/K38qSAHHF
LEkqOkRTnD6+MTiik459mMfcqInxzqBMNfY20PSh+BfXL2esrK4SDcpR9n6M3fHdNBUh+gSndMg0
pPwcRM3/ooTUjpQ+k3eQG+Ocr/vGK7RKYfsrwYaQc60+Br/OsA8J8/BnfAFJqwa57xx+B/2L3dP6
MCyTYqgsWRuAEb0krPk6/suwRHVLIqprAb/5CnTxGLCFej+eeJjt4jFFhOWobN6CO92tnvvBaOjS
bMfi49QPEVrhWBNm62Wa3amkxKn9hmiio6n3hO7+mbO8nMdRBzjG5aYQjwnEeZsseRInExtuRsa6
LulDBph/enY/Y9WnFFQ9hTfX0bUhv7b6egtJy2SfSDXrsSc028dNEuclakAGz9KWKf7DI+bMy7wo
QNR8PDxj/W6aRv48Jam+8DZZRGUerh1fOMmhkL9T4y2vnIiUUaXMzO5hRvdIvCCBxgXQ/SZhIbZl
7hWtMSjCx1VubUcHREBcrrNV5v9SFiyFbaRiPrES5VNKn0moZWtabEhUylQnZQPtr45PQbQz+NWO
2JW72y4BjShgZOwBBOq0XVFci/ckBkp1VCcZgvAZl8gvhYdwI6/Cn/gNl2ZI0QVyAKK9XejzTKUm
sKA9qef6VIg3tZcEUcG3JEPyaN24c/NLN1r2jFaCvPWxHrZRRro4MQGU/mYrOcvKpuWPkGWC20BM
OR+F1CPksEw5sQQZSf6Mz5c9inVPpRoZ3svBAx8osaXVmI9W4ardRkMEx8rWda3LIWEzMaZQgCF6
af8Gzx93KYCRxQaIz0Ew5jQ89KWbJj+Vw1YJ/xdt70krbbRPCwE6PzGBghCMW+06gq4f6HSpQy3u
DLWVze9a3hA4moAbgTsgYAnQNkUXIEHyxeWgbROQ5gV9SS5iR6eQfQOyw7qVbqoyi/U4simsYC3n
TxgqZJicQ3tgbIZ6xH9PhQXXx+0UIbEOhBQYYQfJK8abRZV7VK8sf7nFJw2wICMcQ8iBVDabPdfC
/S55cLQ2e/6VKxtwhYciN3sb5qtZbaOYdmgTkgwAgHi4K3Escbwg5Qh+wdhOl4y/CQLXmaLQUv1u
gJWe5MuImuxrMptPFjRjBk2nf7R1o1r+lX8c5K+6Ikqg22pWMesjigV0Zt7+Psfs9Xeay/OZwfzo
p0uSB5SEFbEXWdK8TG4WsE01WzGoj1N3laKFVKw2FcKBUNVPeAL95V8KfJ7t5QTqXFr0e67WgPan
M0l9APIFihLj52PGH9iNq765BGgIkjK2+1lo7ulQVd9awqCNvqyhKswfTDwOEH2kkiJ5G4MsKoUv
2qQP5XkaF22syTPYnxdwagbNS2U8ImOkgB4jHed5TmKEP6gWaHZZjPijpiiEB6r0sSZTARLVixly
0nhouhM0nlEHOO90BiGKRtTpqEGptAZ/sdntiL/AqVNhAb+9ipQJRXo3FjOAYyahqjmcI/QmByZQ
tVL2FrO36FvkpYPruDWJp8JxaDZHdQryZ/a36AWUAwUS1+o8aH3hgmdmVuwupjuTbOE3ruDxR+4d
/vobV8XQ10pvwLAQCO7x+8CNfwq++lWvAQUmpPbzGrKcO/qTTsalD4ulFn5zV9s/jG0kZy3wIWI5
qxifcpciESnWoS4ODBtIm9Ozzbya+W1/l6KRLD7T6UpfpQFGO69n8crzO8605I8Tw6VR8AdHsDoa
HtQZtkltlsHmI8rXVwgrokzFCfx0u+CsGbLHGLietsPAt9uU0Zpp7V3PBAF+Lo5uz/t5C6P3nkBX
zYttKKboD+zFWY+/Cp6M/M4zcS0m5ON3KgT8hEvw999JwzqQxSHLoXX5p2oQDdrWohCQCwUO6xRL
Veku6rkNpmHr1eEGaUFy5ceoGhkb//A248JRRegEOdKGytLMtW5YZ2ou/zJJK9VGoV7J6hpSpXyr
QSFXTAVeLi/c+EqzydNyPe6ogDEv0FXMGNjxC+dHwmPQ/jWGNpyYETgKBCE8olmTVzzLhSq0B3QL
s9Pg9SgdXGgnkF8d6MIe2I6s0pz+dFg212EDdSeGZ7zt0IV2qUuPHZQ0TuFIwJO3tiTY8HD/bBhn
9L6TEfB6e5wNS7VXkIQuAXDKOJ3dbdM+XQGPRxmjLQM5Hc4+j73m7BcW9vS7XR+e8X3o5yShT0tS
ckPkaqaq8M98KFsjJylrmpbUfYpiCyGZzpId6oKTU+ge0kRbBjWwFSHPq/x+Fh3c+qfuRkFi/kiZ
9bgmEer1ynbr6QiFrw+ItiqirZtwmoxV5xcg6YXAyGkeSCKmXuWMzs6wH3ivyDd/mxKy1JcWhcNa
9Gg1x0KPV0UJw+1/ys5bfp4cifqEQm/JoRalgfB/iQnYCZWYoyzoJVz+UcKzHDyvJxDqEmRfJLp6
fj4gWx2JlP/yfPCxLI8EoFaHArMPmlO6mRchkhN8dj7C6VSS4OXyvNa+4puE06A9d1YtJQk6nPfI
1Ch7sYHaIwV8n6ipArAMcI7tLFTkIfMYpUNcd0VRRnd/db9QXjz1bKdiizEtFvQnMt7P3rbz15Nz
6ZX1z4rByhdgqDPuPoJkqBBTlVia8k5CeziquQbmKIPAzas8L8dnx4PhxvwisNykNwl9XOMbIep8
ncLZ/zzqZ+EgYIFb2EPLuRetVchZNFVZPmb5/zXNkqbUEAQEg246t1Vtz/Q5CeD5M5wTOQK/9vba
GjhEksnbDTj+5PQ3M/a340nIZuQKAnb1UkvY7KMOJrI5fEh488ECLPDEFHstY0JnhYo90udZM6cb
LnrqRko44FAM9bwZxbh3tKftqaNJ9qEJUgsvWcnvzDZ6tnYOYw3JydDTHMxz6Qk9vsShlN6JWn9P
XpmiIhISsHCIQkcrLjx0avtyD5KoXtrmjaXKH4Nl8mv91iGMn3+SUfmrjde15jKyALP+EBB8ZwlM
E5zM16pmU2gANIrCVe8IrqNSsoQaQlroj64aH8mlpBzXpiQoumm/EFXcBtoIh2HheiTypWYbu3VJ
tv4haBw3xWBJ5//AClQv7O9kaKUrFfW1k/oQb7busGOqrdP8ZMFhkx2tTvAiung/o68haOD2R0Mu
34sUIKXa1UF68ZTLqIJ2Ljkvu9GgBM6df5duSS/5aD2Rh/yMfMDVp0YR3WKozWPplkYPnFTp+8d6
Sb97xQsFFBAe19b6micRgwq2cLzVP4A86WCOMdym32FHRAVDrYMVGJ+Xq8aGM6U8b9lwurH5K7Lk
poosGI0mU8bNML2RBuKekU/1Z3iLoGs+tRxMxWJxEHGtuD73d3Yjcik/sQ+Ow206DuQ3EK5vHpgU
Alc4aZFOXEPQaqtYyKK13IZu3VM+doC0DcKLXlYoHF0nCUx6g4tiT1idmGHE5YJ64iYue19Bp8K/
/h5Mn4syrFye3rdSNrvX2wBZh2RhhRGwRauY7Q3SyHbr5LsBDZvKGO+L3Y+uWx4ADCgrll378RTZ
6DJ46TtDi2qgKATxd5dyRzzMzw4QrXSjyqOrECmYvHKhMoCVrpadrGApSQRS0L2qgDhWbEWPkcxv
FK2z2hIxDt8G0eCQc0YwL3/QK98nSLNKSHBlBqD48QoDPKkvjNL8hVLL3HsdevK0HsIgqAPBmL8F
5IysRG+Fe76v7fKdjRNsM9U3WQ2I5tjzBTMTYM1UcDO+hs2h14FXk1KTaXECE9nmiX/gkT0VYurg
1SVDmgK59oXBeYOp5cHscnn/PBPAg0EEG5ow79WpeypAc4y+AVivwEdsXSR3RdBBmLeA4RShAS8W
CUGzk0vf4qJwqt1lWIZK9LtSQq6qiHpAncscfWG4z7VdMwIudqTaFk2XHIbt3EajJn6DzfkhUqHG
fcKSi5ZRD7qtY1blqcJDjmukmyIhfcp8Rsi4d3erWila0IhjoJq9hLrlHk/9APQqWGfi/SUYeJCd
0GGtn6ginvZwWl7lfBZs2xY2Pr3Ay+tZsNKyJXYwes8U/ktwxQKb+SdLZIGomG+oyAUGz4bQWG1l
MN6I6U/dLDRtLtsLjC18IBQ6md0mH0z4SUt1V8KUQSwZ8GNlUhjpR83qpZBKKq2Xb3fpSxwhREA7
2h95mU4iUBC1lxloNLYawV7ZFUwh1UhCK/6cyezkyT8e7HjRI1w7CuuPxtdi4WWHimrcOYomLSyN
Ciqgnnr9uDPyMvVSl6XDy+jAmSDYQ7G1A4502Q8CxXs+eA7vHget6XGKv1ACNg4Se4y8xRl+Qiv8
gUZiY1uVuId6NlTAaMWYtRM51Ayl3X1nI+ibci5HCP469pM8w64VtNjvp8I+igW4mGsHdfftdDr9
1+niUY+dnDGfZ52E5y4dZ3ep/54ok4queMfoN6aHoRshp/GLExNBhZVK98igvtpR+BlZvhngynOm
zJUYZ3CqFm3TSwrCFPbFECwtNMgxNTd1p1o4I0WJOaQZZEZu+i8IqQRKwJrtx0cw0Zi8qJJ5cuE5
9rW/D7P2DQfeTOo1FwtBByq3LLZ6nj+FDzsTZL/548goHi3WPh1u3BNWZgaiebtvDl2AGZGrzmCH
VYxyjCkP2Q1N0J0RqSnEly7LXOU/AxeQD51k08/qNHxcXdvsAl6DhKhZDI1ZLX0Mv64ayI80hXtc
87ynvK3VXXTgo1k+dsB0rdO1c0k2XfRvMYayDAxWzjzTGf8ZoP1QLH77k5YqMuESOUfk8f/a+Grc
1LZ1YLUZdGSdMGD/CdTTTdHRntX6TpvCiemthr46K5k8YDeIYtvJh0rjzwQJfPTI1t7s0y8sBGct
xTt9aBTZyXxeOOjgvn9ROIDxoYTeQlTDYwW+LAJ4ztSE8mTpmR6dPYdtZWyrM8t4lqqOb9VUxOuj
dwaPCQhezPMixacC+AfmHkjvccBNeHu2DOQuQxjFrV+eovpHOAh6sE8t1FToyCVFq0UR8YtJgA4M
EK50YtCb2H4+96EwAoV5okaQbP+FIU/8MwOYuB4PbUaTW743e4+D1VtUs5yr5+4ubgcE1I5XcTfp
kpmTEgOP7CN/Zh3nvfMZM2+t2Gqf2/hWtUxotqmZydvx0ipvDF6fEBJ1xC5aPmlNEfsGDvCvmnGU
6vv7AjHRT5h2O8vpjK3FS+v1HBCwjlmzV5/BUsXrJMLQF+3/gMp5nyfoMjRZqnHM3+7zfDkrQpic
FY8SpXDTAFpelyVqt4af/2noJSZXlsokPSDtIUsmaCwu30FtNq3BplMLyJQfdy/tj3Y/MKwDUFIL
pWO1fK6zVhsaP5oUqT8m1MzFGgbj/PhDnrbIV2qa3XAIoYmvw/XSGv97NvbLOTMxJLrQ6tVZ1qMu
4DThGWGjUoyCy5lOM0xyFP7nEOmYeRcBMrq21Fr19UY4zEn1rfBBGOBn0FG5r+eKLVHKRLAAT+Kt
2y6HAFc/HsNJmRxsxeLzl0CSMCo7V91OB2yIIuopsh927fFFMQv2QqZtwCaAf/azZ+z13/UDRZta
Zsy842c9VVrvC2i8/fG0ier5GO3ZuJlZY6frEfru/4iGUHGuByICF/Ktdw6fOL7csZFL5JKS8Vhw
ZNzVEbvnZSJwDBbqFXseOTmjntEEP3DCdFLr4IkESNdTwUAFn/zs+qvuDzP09+uBmcCR7/nWWFv6
lsy8OXWVgDyxn12Tj/a84951JTntSo9Zz/NHMWOFBPf8l2i01EQ+bFksuvC8QvAklaQEOtpgeCQx
3y3ERVh2HaB5Ir8NhMxEdm8zjBFKkkJVz834CiUdvMluG93nlsMq4kFHWC3VPHlGCvSxXVkwVPYN
SxU29v2CbFxdxSjrctxiIWvaZG9g6mTzXlWaEK+VX3wy89ACSr2ypZ1OTUsb/uRLpICEWJIDk7cE
6Sg8+kTnyuk1sAVfZN1QFOc24JW2oFYDwGHU4AwVDsdsCN1CNXQJ0x0nRywDMAdi2WpS0tuUMW12
KRO6tJPwNvbX/PU/ADZtGtj9t90ZMVakX+OZEg8ALFEb1kLRb0/2RPQ302qQWBX+WmgSm0lkflgx
SO3YSPg5pSpFAIoyk0UfnOkthy0IkUY7iaD++AiPWWSZh8+rButq1CLOknTYVeqqXBPFkXAu50lb
549B5YETJWVjpFIYsB0BNgu2d3DNGelsPxTH7oiLrexowOtxo81A/lZKhb2U91zEnIVzq9rGidyk
1wAsOUxHfW+YFxXcgLKq3Z6IlRyDXomnPbRTTkDDSRikwPwiz3mw+c642BrXJW+m0asrtR4WUyN2
8smpPljxcOnekJaz2CtHKCfvHZMgx7R59v048Y0DtkXCAiO9MzoZMfXfce0BcRP3SiI7GESpQ9nD
pmyvSB6qKzMrSWJBDcmSsOWG+cXA3NDQtGk5W/h+cNcOuJvUmAMyUkaTRb9WWztYTwBPbGyli8dI
6VzqiB6zXDtkKCiphD1Do5cPqZs5R1xG3FUZeEV0cOCZdnJjSEOU353Lavy1ybE+SscoMHCOjG4y
YMxoPLzJjDyS0IGIWNfHBFgT3mHbpuliThnkLuNXKlHIO0YdsWrBYPh4u+PxmZ18eGNyENNH3beh
825PWI6V8CPOtDZl7rfe/+4XpA47q3TCESLyG7t/RubemnTa676RqgWQhfBjv3tI6Xc/yf7fK1VE
vezSHdIRIaGWhT0omqH2o5zwJHQN5XTjS3ar5E+zMJapANfIEKMUb3QRyOVSHV0/VdpUipR5q1wZ
hfjjDeZTQ49WY72VslmOGSNpVogGmeYouC9tNlxPt20NlcDoJib3qvuweo+FuoqnScO7PzlCT//U
3GGVZKT6l6jK9LqvmYSoFwJfoo4p4Qe+1zNSB8T/6TbfWmp0E0AXmbFdgMAiPW8B4VCa+3UjFqTJ
4PW87fseKY6C/9+TUhmGq6bdiRwn3DvviOQQUcX1n84zwLoXjWblEwjRmgd95BiOyjyn87AW23BL
v78aFsEMXM8kCVcn0lXzB2t1scYCRfbP5dtxPg2CJoK0uyk0Dm9dRsxjlZodgCpOtk7N8U6GI/co
b8ToRsWaP6UiviSzvCTJNweDdqXyDF9e1sIB3CAL/CzyCD5FffIBL3pnPb5Ccs9VnMO7PtNA5EJB
4irLM95+U7fmD/dq3Ar5Wxl6K8bjnnRFzQ1kIMFig61mMLelaizKUp8YzM9JRj6oXdx3BkjmIqC+
P1Rc3IOUcFPkQ0QncTkNNYkNTwM/I38tPXqrsAJKFvNZXVpYCzHVrr8zwoukPYlWd/f9Nf+KDh/o
z12X02uCFpFMAUxTI+uWqNhhJgN3rBPzdyqFk+d4A6M1YWOaSFayi6+2K3Cnos9KbcWhPIV/uTkc
2udCprWUe4q9RKxoA5ndEbpYz9DN0AGpb6KM0V+W0azEsSA+WWfrZ6v2Waqo2r9qNuVOtske0ORp
MsAmhZwfNz34qtGc1AuqJLxkTA3TwNZ9rHzo4quaZnpiFD5zcw+jE8QrF7rnoly8nsaxDnV0SZ8J
VS55w4wU7BZui/34RfIqbMmAaCI8SKNFn5G0y4jYnExS7k3pYJsqghGxU0uzrMpYoayHgIPNR9V0
vqEYh9YMm9HMdVVh2gh5zjRy3XkrN1sbsHvOVbhskOpiicWP3ui5Rpi2DpysmrTDjiusJuMVcATh
/1yuD5nCwSzTwD5K60oWNkTsRIxxzU2dJOGKG/5Hoko1r2fvV2wa8kj6C91ye5aAzluNNm/sHQI7
il32jj5r1iiU4DZWH+aJJq2Y81rFTNdVk8sTMGjgWoGuTGTmdXFXTDwZREvEC8aVCjools77cVmK
zya1fMXT/9J4AwJ+Cn7+P1m52/4uX6tgt9dZIM7XscAWC47TmotOjzJJPtRdA9gYzLpxrljqDpJy
R/hBV5R9ofKV3GBkzKuHrgkNRwqh1yaM0vVpampUNtHSAK01WSRLrw+0m9zsma9z8AXqqBJO33yv
FR70vs4X4Xucl9rGv/ukQ5V7gAPYYPSFDruwtRND4S0LNoj3NmU9XsSC+/qT1j/CKjWIm/bWeDM8
y04JyMybpyfBPz5G0pCYJyeP8PAThM4oVZnCWeqg7QoE+tIE+menaDDbb2r1+6BeMWz8OnluvNym
Cvor/r5oUTPuXyYvNMwTRGnkq0MCgiUgTud8ireNDbpzmVCMInrIjLPEMLYhk+b4Pv+8yrftqmrF
YpjpLfT9blZzwizgILaHjdy+AV6nQnwmgaFenTEhxvAGOO0NFtM1UKvQuzuXdNiks2egtmXfQdkT
WwAnKEDIaAQKU7OCBXX7wAjn1/3tgSkX4rsrGkFJOvcWJWHi+EYzUg+svsy0wuUx3LQlsjYorWV+
gOwYkJVglyU4R0vgiBpwHvnBE2x9ed6CCDAIOzUnuwHgF12Z+h82vtZgG224taoC087LBX6YibR7
LRLBl3cGyo8b2H1Ac0iF0i/J070g3unVKwbIGU5E+u179hPbs2TVhZ6U7/1xDDkdf/w4PPytaTFd
lb5/uabGJ+MwpfiFG1sHv1HZCnhjY56n9gIAqRnp3Z5PBqTdG3MyJJqHdUdwJnCSBpryzspA5u7b
fZZ9ay4VXbVUKEPj0gD6I62BxjEFpYoMXLHRQn77eFtXD1wbVziYUXcsPvuqHh/famNeV0r4Haox
lMP5ELTwxfcG8OK+EUpTwWcb6QpqFyT6yirLh3Br+ICo+vD4VDDJP5PG+8qJD0P4NdiVi6D7mT3e
zHBrEBcRVqjmLK+GuXUamjJWrp03w8PKapIqOo0jDW08NX+n203FZvfakQmD6HtALg57qLMmLjKY
F16mydFdgJ09R1i9opzPZE8HL6MPuJxHbN2fqJsfCA1NLxfAATeuDpoOSNEwzR3MjdrWPSVN9Arm
XZcwdk61akPogamtzR/7KED5iUuIyRqDBEK2kuj5JQrLynrYLzq2DLj5pDs+lb7w+kXK0OIbmVe3
9jlFWg+bpLTG4Bm50F0aToN9XaXq+Ptc85F2akcXJHnTufARc4NAMhs7X7e9IdL1SMV68PeILJCj
8IImvn5GU41menbzglxV3Oov0xCIFjI6pLHk/DUbICGubEarg9sKWjXf3sFYEBl7hWd5YikT7E4I
LxlAPSU0nq+7tjZZuQE2QYNO8vIU2FYR4M9yRRpuhnBCnwUOWmuWlYCOa9B+I1wPj8nBM+ydo0Z4
nyYRL/pwqEKay9Yg70v0aWinCbvEWYxbp18LUO24/9H/G9O6lfqrETyaxvtp4pgcu4cUCD6aYjFB
jav3ZxbztEhjbZJNSYEPV+nIF0WF5rDG/yPr9NiVo0CFUuA8J0xjwPfp2RkwsAZbPkuH+RZ3ddwr
66Peo9L9AChGpVqYK3FFVmkdRSOfdx7rluVdifQuugqDJY6w3sS6ZgVxjM5X4IhNud+MWwLwAkld
K9YJ+e20IM2QnrNwIRxU4DbYOGofqzUzpZNxWnvCeyRZCu7Ie2vnkf3ul3c8wvM6pSWUv0cP/tiQ
ToylhHbk1WFE66bE6KPUz40wMN8NXS1eiNlaLXnMaJH6I/NQUKUbnWFRt8D/kbt5XlSR3Lo0EorX
w0OaBE2RcVJAMH9cEaEIBLb6p/xEOAxntr6jZHmiXZAihg0S7+k1KCrdJpK82FJ73p3bOzsvY2AF
Y0TkuN5r5sLUhCbHHMWCr7Oer7ca0BJGdUd1D35vzNv/0xea4vhZZ4RoUlsf86jkFiBlg40FMdJC
OYE7FzybqODbOkONMsog3wCdZsTIrH9AM3RoFQJGwHKbbsI+14UwtFKbKrfhR4YuDlRnJQUSKbXL
/FwWkKf+nPMJTpuaI1xTYx/jESzO/HDPZ3hQMYbg//f0Zsa3f+9OzjkxQwLw2js/5cqAs8cWhxYK
msfERaTF/WtsXvlDbFRwLeGpNSfpote0iGgGDbJkzGH5c+tHo9aQLaXGRyyrFMh1fFw3N4kTQs5H
jEP0P+funyXiAau/0qRp66MzHSLwMpfYgFIyhnMmkM9Apq/DIryjP3BgVcZ379ZwCCZTLjjnb0+/
Gsu5Q2KJPIxJ5t1KJ7vWLP/mKcgghyXWmfExUH8qUXTXrF3mPujUVXYgCJIqRNDHcylx9r8Y3kNO
zOfKtaQmttpqcXmhDg59aQSxZCpVlsF4tlUuLqp0bszRrHxSGOAPdUDkO/yrVvaq96tutbmVz4pw
NLU1jIbrT14LTq8v8ElKOXs4+5mIGk1b20SlyuUJBhG28G5wKuOFege61ONlwUFpIRxefryxG3Xr
k4BrGh96ncq8rXk5Amjc0qsfrI/p54+9IUgYt0Ws0UEd6QvT/tPAS+HxYIT89ozDC9ABMEGVYGBW
Ot/eNlsQWaFgnI7MWFLqpLgElQK7aVSlML7idpHhVbvhW7QT4jFPrd6lauYr9uG8YFkyKrHJs/AD
6MZt5fYnZ0R1gUzjbTCDRblTALrfrhqGhJfN+ZVx0uxCvv3HDPZMZGbkmQBagngmSf98ooTe17H1
PHndhpMRPBv5zYqYJ3rpxJE5wMJBms6TtWx4inZy2l5GEYfaytOcaFvcEEilsBSfqblSbsW263hd
/vgAUIfIXImYxdo6n174WxMS2AY779ba6l3oolRqfz2ohfDYCVGM01oGbC5/VXVmAm5v7Z0IVMEP
fEqE0MMvzDuk1HV5yqkVfcHOPsXT7e2ss4/6B0/eSTaYehfqDw3KkgiafL+KbpXFFgqSBKbv6Vwb
QA4xhZ2RFZbc6d0JyIoTsEO7WQ07y5G60lY7wgWxomUFU+2BNKTo/WFUbZO5o82v+4NBMOIr491e
V88CaerV1LhcYplrwl71DiL6gOINHaBk9pUfEXmeAB6+DT8qT/6CTCmRdBeqVlhY9gCr8tRwV31A
NCUebmwJ14wrHJUlXYS4f+HFt2kvTHEbZW7IEi3lSHdIUCOapbdsPyjyFMdWTrWw06IO4oGrxfyC
xhHqWO3cUjXr0eLRfX8G8m4PxIPlL9zDeUQkj5c+Nxxz7FPPo2z33D/LvFFZ8zqxUXnxw3x/u3TR
2mND6ph4e+zL3+Yk9+aH3ZD/pgYVh6Hdpsp/9ywpPARdH9rP8T82Ec/rmMrbW1UAU7HLBDNvrB31
pFGsEMb+h5kLg4NN7Syn2cBZWpW+zJM1cZtB36rJwMlgo5jgqBJWTtCFNLyxOsSZztZwyydM6Dz8
89pmCYL3zeTSAP00smtaIzEJM2hTJsUgf6qhPfk9JYexeZrBr8TFYlCCpyJS+NleZbDaOdOQHzxR
S/j1/p7wdKGC5hkp9JttCvLBdyy6pqi+BWV1hA2Y/blod2EMzJU0az6e9y8Urn7P7PPYhBsl3IdC
iscr+uqH3OgqRi6c+wtov2q9POTimjuzbdrKpe6RotKZ2+xZ6GlBjNGg8UjK6wU5Co2afYBaeY47
vai9EU6C92gSDfsSojKUsMtI3HwB038IyUluFCwEN4M0Emzw28GdwINM/Pq8GGhfTT+me+SyGyAa
CFTDIAe7+XqNVNhnK8hX+H5m75Q0dVzpT8WboSHmPZFx/DUtIHJEw5XeZpxYX0h738IG4eDNd1ux
T2EBacRuJK50YZul2y1KmkyGtN33ZGfFKXAjaWx3ptRuMAglecdFKh1I1ruwzD6MD9MpmFW6qjtC
UjkugwsC/SPDFYxOvUuLUM5qgoOdq78mrVvTp4Jp0mrPyPNuf0+Ix1JlrH0bXdyxLHvfQiy0ocjt
6kb7V0xG2G74uohSafQGonuhvnq0UKbIUs71qMlIqJCvlpe471lp9f5p6f6nL2De+txClFgjvF8h
1Lk7kod8uKy+iK5mXxUEIW9cgbInGHPpxGWtny9Sp2b5qLWohq/21+04jtrSwL9lANhoxo0qDkO8
tVHZ6279zaJfJTaPRJa9ZY1lrVQ42VSRDf9Q53+R5ag0XKaX0sNNf1nqVn1B2vPTYvh5c+DMhjJc
f0wIKj/4tJ+WNMvsv6osP0f2hvkGKudsomeE3hNP3jI/RiqVjwStrWEDxb2oYaT8dN8ol+7vPyOh
h5Kg1kW0qWj96gglNMcD4IwC4lmMCuSbgFvKkkYiN9kdNBA6FO0maUb96rICB+QGI8W+zCfKA3XX
xyYmn6LKajqrlHHpQ03gyPP1/R+vUK94ieEQWTAsOxxjrhBaUUzwyf9kRehSJ1peuIs8V/bw+npz
mUNHGRAYa7w4RezMLmXYO8kzcHwWnyzt0XA0YALK8pPn3OfXlOCT/v+8dAKbanWRnGP7iS/EZajs
e85iALOqGyjr0ES3CgP7nPnW6FjHweUsqrbSh+cOmftk4ahzbokHY6X6WT2KV4xQX+JxAH1g0DYU
/Welsa4OqMwEBbOsxesm5fJ62HX6A/H70g0h/JZFWUshHsICAipUjKolMTUGGGF1PhqIUZ5X667B
Eb7+2Z1dXWB9cbC9JaERo3hjbHE8R6wAVoMHSfi5jgeVKqHDNYeNP3lLtX8USbzHtlHl87ulhLDP
mWbIjcJ6S/V5xubMGtVNvB3EAs1jm3RfhODXo9GaLhg0xlhoAQ8y/MAERqOupBymKFk3tRc/IfqH
O7Dffrv4Wvwq+Ax41ON7uorqibtIuyeImtuZLFNZfKtNpNaCycekjDhZWgCkkD5wl1tpvcZLZH0g
jzxaq2DUvbeeLAtcIJ5t5AxNR4mCeMOLP1fUUFo7JIR/ctjAxvw4zfxnUqQgqtwjPY8dnTtaUwF5
ICHVufV54Ek0JMvJ97hXIxRCSjGVVqgdWulYqHjNsYBKZMOHOwUIkKk2YWbfDn6l2uELL8V+DB5H
Mr3XBsujvpWxvjZv4Fk65DH+1Li5nxmQsQmD2hVhFSHfhZOzef/rFhVyE1VWBewl2lKxGdvU4j09
M3mgangWq+e8ZkC1s2YmhrRVr7yNVjbbIpfCSlFg4zxs8QQ64NeNG7fapGzG3SG7CAgYAoyJQWjf
uv3x7O8NHl49+tdy/w2NS/L8Du1WrIesgpWWCP1n72iE6097avECAaOQC5YGfq0I7p9c/b8XrDKn
KmZkEJAmFBfVgWwDcb/KRatTX/pbCqUeWeVSXybt5Uo0EuNRs8QCtUNIFxUbTaD9TaiuV62VPYRX
ZlybVtEcOHBfLbMccEIgQCCISjK931xNaojlUxTngfoFa5doblhO8ITTay+uJPJKg8z745yaZ54I
+QJDDQtDws566RZCY2ToeBpCPSpOwhKHeUuN0lQKifg7R49BAoMV8g1yp4S1ivdyqD4PwqxfHpBV
AlgEG26zUKY8OJNqivGUlD4SWEP+I+j4h1wrPBwbd1D+wnt1QqZe6UpvcaGVRtRvWnetKPW2y+e6
5uR3B2+d3Ru+5/P558iYUfz3XN2Zw0mPuEHqBd3CSXebLHvqp+J1WdYqU2KBOJZgzdtbpwlT9XX8
OFb9Tqce8wCmXcCyaVISlafKwy82zpsOfQhQRbW5Yq2atzJ1FZKUtM8HckEstKQUaAeKT6QqMfcZ
p2ZVDFX+Xzgp3rAqiGJ7Cyr5TfXTf0vYT5soWmLkm/wmnnmd7Xg7R7z1jhlpcsSxg5GNSq7wSo07
zSy3cCjhV/ghS8SS1mtQXIUVLfnzEyzFVt9D5Dwmm/ncqHrNzU3CA1Yi757LySkHcPeaZA2BgGoZ
4fUDMqg/jkvAhN9Q/e31an17B1s2eLxr+OVmj2uOUieEHZCfJjNqGMfDlqX0jb2lNX7iduDpoTih
Hn/w4RoSy/XNfSt3b8toayIluvoaR+Cx5rJhoVtJ+jajo7S4kKCZfCZWIw3JjHw/y/xNeWAW1qOy
pHc1JoV4G/TPp9EdXmaW0lZDHvqCgJv97KqzjV2Ac0ijvs2yq9vQgL9nxJonqDCjPV9iH0HJpN93
NueziLocmGyTIERkUGCUQWx/8XCtr8s946q6t77A2L2c8au2PhHjHS6eNX15slMSWYioy/opolde
DCOdZ1SKYqgC40P0V/2lmqbbgcAtYouq1jJnCKmhlmTc2A5lORLl5YQO+DvRhf7TEhlLNiT2/7D3
FQ1jOmxhMXn6N2rlk1oBJQkJb2Lpm/oWZ7v/2L/Uj36BKJcsIcq3ISx6FZRZ/c9GrBBov6aJLoWy
QsLSx2bi8+XOKYIt9sfbfu8pAmtjyxqjr0GTiV/yNm3uVbVjUadpnRvMs6+rMd03/+4Nfy2ml7bQ
PsfQNgJf08YTyHUGsRwosN+bvdM3SJqStz9j2qPeA9EIm/Tz0fwdn+tkVIB+rLbuQ9wG871M2HSA
VcK+9xrGmtXpHuCa/cDzwmNUO4Q8zfxm2ujqmtCp5Pb9iFUW6ocmdhhqQfbuOlJVyHCOyTfiunQI
/00pKJ9pJVzyQkczm9mil6AvjH2lt0FiUf80aSk6P5NroIFPXMdTe9bjWun5ZhIYbmHGcV4/go5R
exb3tG/+Nlt9K72h+eKlswvMKJvHVDlayLvQb9WmQ1lHA8i9g+1ItM/ihaArX4iz/POtufeexHpj
3FIzUH7IwtS13YsNDUIqz/SAsydMIgNhn1roPD4WgiRrfDYFWBJphmdCCy4YHzn47LhWA1veZgsK
TkeUtvJV3QCz/cXT6Lhs/GDqEP7j6y+86zWznJKKqphRqTeg1+1WyP/wmmieAqelCimaK0gYd6qF
quEhGw4Abx2rx8gbftnkAjl4+VpMcvJGhewpWCqZ16P1GHRxpqpDzFexpSL4my7kxzA6cNkLgJPu
uARw0MQeYqqIbOYS36An8tF9Cypa2O6Tk6kX4o1z4eBvssYwKz86pBG0RI3VUaTuOnL6rM3ZSjc1
j7Qv5rZWiRaGd1ZspOboMCSuSEz/9v79uurrS0h1hiWFyH1kcHZpohtApjzKCxwb8em0h2mWspc1
tMAr8cfMLieXt4f6sxR8SLYvXW6LaYt5R9zEM+wB3Chfj519e/M6xrrRYme+j7H0N0zxILJs9ZxP
r/gAaQf9G3Y4j2HLY7IjMwFj/g+1l1XWZmHQIIeT8dF/JP4fyat3EkLpb/HhS+nBX9JJ25zPrRdr
jG/AD5q7Oey1WuYCSA4iZSVaDqxjmQTEE3jYzTNpl1n2PqlZ4sJ2+MiE6u9R7VdynpIljOTD4cKV
XVSIIGSXJbjLV11GiZLfX/IRSYUYo2iGJ1XStWkk6icUtQ6fHr5vDfkeYwhJKasV7C9flMhNFZZA
DG3sTxrYgGbFG5PkmJ7SzIzL13wLqdoyDYZv31rMwOb4xSmOWHTJhLu0iQdBnzYuxSCjYMphSwci
9i1Pnl7ulpx6NHSqabKBrfobGdbkEO53/FHkY9gkRS5gDWBRlbvXzk7STTH/N6nXAGLEQjqH0ARN
g1FYP3Wge3ClwbapaXlhRnhPcYsS5Gf4GO8Esv2vy0ilCu3VyllVe3nJHjJBSebgbq5RKW0Dd7hr
PcyxBQ46m4wMWzBL++LJ7uziIm9dSd3EBOnTrRqwP1WjniMqdSQ46k2BWpgRVjFZKKFRqxoChazW
PI4KzgJeQlc9R2T1ZYeplIXWW/crN5JhSTwMsIIM1ScWGhPmeC+tYRpMS20nFxfth93IoaANdSf7
m3S3C0OJi6Qrm8EW1Xtr+Ren7RcYhQlvGN1j5/UJsHfhvZy9QQcbgK0Cf+0eQXwxJCmlPx7eT9rI
ope9EKYvQ+NZn4bmndsqdJnRrkGS5fnlMzdEkKTIfuMijnKZm7qaAQUrobV1llUAcSfFZm45AK1a
2bDigf7+UguwZ1CShIy5HLIfuz/E9CcaSpRanMtuL6ODGJrlxDbAe6pgBONUolfMzKLkVF+zkwYz
CgWDHAYXEipTnoic8wydBj8DoJj8pPS0I4dX2AuX0sMdBMMUuz9fIjX7jkivuOzkiKNxEmx1gGDl
v8iPxdZy9Go6cJTt9pzrK2t6OOq+BuyUks0uCItpbfevtD34lPrtaXGpPzoW8lKuRr6HKk63rTB/
73onK/nAOaZnDbiLyo1hmm7cAjv826d0fy21TW3182U4+W+5XaRt2A+fghVOYJa7iOfGDBQl/mGc
eXdHaYFRFx9Rlw23J1vvTcib1vDaVXKx1O9t+aD7VrIitJ/JF/mBmmy/SEdt/86jDEKqsxpm7ZBJ
zg+ApASGuyhF8JCh6DYoO4IiOAvPSh1N1ig6hJLna4nuf08TZJDr0BcBeCVgYWgxqBjvWJVrQvH3
C2NqhXXmrC5zvMTMLytVyBNWseX5P1R+9+QZXR7xfe/BVPjEy37oRjfNMpNpRqt3IY0ILumXflmZ
AXEYH4MaJP1+VBNYIjATJtFtEbnOiohiHk+MwPG2GVeedzRPW+JpfSBWMpyLA9sB7vI9SRgjOpNl
SKzN37ciei6w+POBafaGcUv3baRS4rTHz7RSVfNLTsNsG+VJ6MRgaxVlrT5EzANdVh5hF4kam4hk
JkC94tHkjrP+rhY6TstDzy4LlVuixhyFwI4jj78RBMkz+FuLtdSy3jKI8YAyKADalqQryIMXp2A0
fSjfIX+9dysN8RiD4NyedSkKEUTP5u/EgIBZvSiqwXt7klbyLvh6deRzlx4ZigGcl9gMxz59C/jq
6px2eYoRoADDmm36wWZM44ALT6rEr22mxV9TNyySDbjC3LcIr8ZsnPmGLRJ3F3WrK0VqYFx+m6XK
VuZfPgBSDafis2I3zIx940ERzRvWF4in2b9ShPWSdPNcJ5bxWGuRFmgNMTvmAEf23kSQ14TEk9Oq
6ko6hqNnOTKivNP7FtbGanymgVN6jEzQjAr5bvH4o+EKEvJmVHy2kUfmi0lDm73A9jZyDbZRKZmD
3ycn4knblXiVXdixMLCUhNtGKYjLFRnNYKgWqgr3Izy4iuvay/V+Ya9CSyR17BB1Udg0i2p3s9X1
9mTdC97OA1MfmZOuaMG9/b3bQl2vT+AhbmSAEXH9GEeg0lWy9CHf48pGMZEPjyKofX5k34mtoUbl
TY45U6GPGwtQ5EoKAY1dimSFOT5cIcBFrApXGIquQ6IKLUMjSS9iNJWoezEuT5YAZOUzyMNSa2ez
ph8rw6tIuK7TeGkTi1WYT9vMtTtCwyfdAVmfU8LShsDaTXaslMaM3OI6+cPTRZPO5lH//Sy1dj4k
QRavW3iYlRUEqDGzdcU+9/WE+hba7JKXyt4ToWiMqX+q7QChv6w6GWkPCFqEx+E7U3D53KyKlneu
Ep5xiGUpL1rRdawe9BpuSIvAFavwDlhMZJfQCUXxIflYKGOzMaWBnZhYJ+6o6QesvRQyGme0NTy8
/4p0z+/svPi/T8K78eHl4QGtxeIeSx5qEprbMQYyQHh+pBhBYGAIH/OACtLyqkwPjNFQo600G7Dw
hNOgyTXqL4vtIHXD1RqSzIBmqjGaAmZsgoAn4XyItg9p87ymf6FAWHhEHBQXUhgqcnlA6EaEgfYp
CUS9L4nr/3az+gOwK27LwU8L+yOFJMTIXyRGtR28/W/EfGhp3bJRzwqg92+N2VgTuQLU26Xuedr0
RDrMYXBxXqqHWIpYody4qTsx8ApwrMkUmIGHmUyidt9NmW0DT/5c//QgxrAlfpGC6GolGYixaEZK
Bf5BsFtmy4rek52T11+85KM/YBoAUuvT4Ti2AjOhIYnveu8tVcQ9ciDKesWBjZaFFnOCrambOC/x
KaOCd+uom4PY+QBLzF4IO2GujhQGpKqIuup0se2OC0EHVpOaedcUJ5AJD+MrMTrOtNLMzceFNXJf
Pss8NM6JfGCwP7pwLS6HFBOBEgvacMD+aewXVqOP4KU5J9ohCOJo+tUTAmYCq3dVRGzBj5hDyskz
hp1mWdnKSF1vkvJtyA3tWMGlmAKZCGlwHjeEHXVLjYHW9gFGQO9E8frpaD1atG2pJTzUqFXxnhpk
OpGE+EMWeoh5HfKllVJ5AdWX8ZNn4XWc7udcPRSTm1fxK7vZqLBrC931QQ7tplZvNGB9vlMHX0h6
kOew+vd4WQZ7mn5fgUbqZZVxb5e5w6rmkDcTNT6yskrry5fVtkkOaxv5G9KO9MEx2s6C+QpC1zgx
9Wbmvi9wroUwsfKNqwrAvWh96xc5Od8N18HuJmmzm5HnBkaeRTP8AbwMbk4ZUPKVMgWMOhJ+63K6
VOELm1TPeorp5K0oxssA0LByaREFRZxwQa2uig53b0D1n8uNw4/tPqSqlZIToD8AXPx5AHl88UG5
mcX12/iLqbO5h1JYIytHk1IivmdNKtS24QXuFK4KgmVVp6WsUsbV0u6zjQi/MeUd0qFs5g9EaYuA
Pa3x8pyXFVjcOT1GCwIPHKuWDQWh/3j2W3nmCkRmUaMGGAHCI1yBOnq23SQovxqj32XZkNZqM/yX
jiJwbjIa3zYiWg7//hl1MnZ8jFBBfrzVPZZg2DYDwKBBAk7RyLMByRlzkKFO2BvUIYeOvJjyUqKn
CDLACTbpWs0ROHqYXB8kdc2y8aVheVy5TAz4qeOlGdtvgqZEKStP1ODkn9dtSU4sg3qfFcQcwdnl
Si9SNc7Nl6xdDZta1E4mcegYv9XKias30kUqttl9JQqnqCk13HMd0e4dh4vMybpPO/GH1Sr71iTZ
7A8LeOQfreXGF4T815iJ5Fzn1+CBR5WdNuud4hTJtQWU1yBB02ErJUj48TKU9KNaK3BfbqWEq0Rw
FjXMdpknvXigkAdG7k6t4fOLcxkhhJGSzU1HQnwhaZ1YuTwenKDWUjQp1OsECWfUFqqZrfOfAzBw
amQOJW9rAu98MAJ5/pZXv2J7/LO3pF6T0kmO+cL0PSZZkVcvP5g3NB2Fo8XdcqfCqzKFZp+jJo2W
CYMksHurKI4bA4Cfmit5puavqo18hyqxOMk3p5QYQoxbdADYTFcgaSAuBQtAC7wHIQJOjCF7jdxJ
FKXVQi6D2Si+d0n1v6Thv3VrdR9fglBOFOjpLufm2LOiwQ/Lj8aGr4QhYTPeby/NUU4AQ7afKgFV
1xpC283uS+ITHjDOYmF7pdSFc2Aqfn8zK+E1Dv1FDLnSZxfwZImXsJhYosa1H0tjMh5jRcDBFE7o
qA2dIQQcfDcECKQIPLlglt5aNLhOU8zXagiPat6EnxCqDJBbWWlklgwdQpUGJWOZ0ruQ3weMtKcJ
3QIGwQFiLumLjP0ZSrj3sh05n8N8zr3rfQIpjm0Ytyrz88ZkijLjCaV63Fynj4szwn94bHNSBaYc
4WjTGzwWGgJu2g+Buc0zU5R+eXRyBZDE/Ort2SDJsSJp3CXVmTE2g8oNeU9aQYmhnYRuH+1vDLKi
wemlKYcxlHuYnsklr++4qN/oDQYZrx/MF4sIXKqnOmcCT7TDNFPDEOxOcE63NZOtAwzVI9ulUnRX
0xVdkaNiWi83PT13hHDi0l/e09L+tn8aGvSetwO+kuXHxgQzNYwceaWUTC/tRzl9OwS0ITYTVDOy
bLJ64MNmvxQL2qJS/OQ9FpSjTxmFdDU/XU8sMIHUCWuos0tpbIl1QuP/fgfryFV/Ogd/kVEq3m9b
/7Hw6Be2uFMVIasHrIwB+JPtKde/ttkRI6ejcuIKLEugUCnn+AzjRiJEJWK/6pN6vD8QoWxbyBsp
wqic3ifaAVFDaUdEOfLC1+Wng5AdLNecX20DaO+TlwjZYLwk6LUg9wG42yql8Of8/VD6HwHfo75/
c3KTB5NclQNHP8c1BIOR1aOi9noztDKR8g6JH1I2WPdzM1NJJOSu5F3S4xJIJRya9dyifw8wq8OH
xGWNPUHFzZ9/Xul+RO9GSkLuar/5AQ3Byd1gijdIe9dxiV/71g8idxDsZsZaZJm0Bpbdkrl0rijR
ZdBN8C2VmSXcrb5GbcLQNkHHyKAvODa4Z633j14s/YBKpsOjcYuIFgZjn/nEI+fl0hYm/Yo4z4Qn
0NzxPgcOoDQ9roXbwNS2O5ReHP3/DzaZAmTplnwgGeQyWUuRI/frBh/4yK0rEBbzWEC1PXGzEvCR
RgtJI5l+VafIwgEHmc2ubJpmm8CTS4U8kpaKXasclw6eRnmaATXeKYtZbfbIpwUjMqJaxNcu/ohj
cv64f9i/3/zqhgJZDYAR8tXLWOAEhDlPEjjb3qqRsX16JiPsoFQPXxEP3L+ww6BWcVuI0Fc01B+w
/joOs8WkXRp0BdMQXaRuKFltQbnobdoGnP/UMhyqtUXp4FnyIp5D6sxug/3zShEcxe6YhHuwhyQ3
wjFKdNWThIvoHBk4Sj0urQmKF7E4CVU13XOhwn1Pm4F/ZJQxidJnrI75pKdvpEpL9ZgX/EsxBVy0
Up5dFLQzYGSr1OC8Q26NTbuy5fOXX0PUSUiUThY93eC5ZK3CLORfpJ6iZ+IAAGfJ+sENfnUS6+QU
XADfd3WjfazkOoVHUxva78pJo6ehtIckUUkmHznp3FWQhR3UzwuEfdb5C5F2sufSD3g6JNzLOcxk
2gQZYbR17xybT4Qgk6moRqGzGSO23uNku6nQVMW3XuM5L3YH7rPyfayY/8+PfrDZEOImH4F7oXJB
Hjy9IuOKD1iy0tgfTkp40wFgj8J9Ax+2FKZD1hL0JfmLScMiUOPNI7hnvKhIHWRFeF7tDi+XCPLK
CZaWzl/JABe1qLy3/rzwMcdjngQZdduxCpsJ8cX/Ws9gitTnptE4doDCX0mMBjGk4639Zl1+WOxz
KPh5+Vozu/EzZ2CetJdQChEhl+O8mx/6I5+KuTpYbXJGCzlSG6zD8Yc2I4yrdUmSqKyL7H2iw+Am
Jf4qeo8Wzs3B3osntwgNvo/54n9/6pdzRkNVEZUHh3caKVjBN2V6E7tbWawj5JG8zoh2Je2X+nyl
n/tli+Ka+buhw/EjlegSvlMe4tklqRDQuXDBbLpfLl6ko6OtNWboQGPbhvRGz9azZF83It1limuG
dCIuc5Inbt6YoVEiQMrj3Bh+oZLozQgvSOBrSYxKbip6jUePigyQRvapgrnUE4tfB9GcAVmsJSN6
fk8Dp0ESbNWwPYHEz5EN8YTBEJKdkQBFW3ZEIz0GZMp5JIg51b67B6uDzhjOkifqmKykBdkoJOZg
K08n1fpEBqe+hlWInxaW8TGKoHGuchESKIOoKeCZYE+6ULROmv7/KAUNRUbAO7gujDQfEWJ+D0NL
EA6UOri4mpOfHkDXHmYreZuqAvbKwvC/vTRFbYByFGYyKPi56l/fw+pcwE5uIi+3zcBn7gGH54Ib
B3J+Hdx6eJqktZLDCjJAu7lEIvNxB0pnZc2w/m9PcHOk8m8QMGv/W3gXkxWCWLG28bQpQAGvnaUY
0x+H4N0ouR7QaBFJ4DWhO+yaesXgo7V42kapkR5oJ7TRx+HhpcdtPRodpSyr3VXC/m4CpUW7YjbM
AY6l3HZs45yEdFqd3HULpSf/W9l6FZVs2aYdldy1PFnuU56Ougd8rt0uTTG7JCYf95uP8OFQXSt0
2hTek3emK5ue/LuufmiXAkR7uW20z9UmEvtKly+3xupDi6Rg9Anfr29i+Ye/X1kMDASgyx7Gvnl+
X16RB/Xr8gDJQAQ7igeVaOT7Daq96sHfKi45pg8D+7FuWyOMN5hnOeyv255obSmCu2E5VSMDEEb3
qfUgoe7IRGoF0V02DMPnOKB+2rVLrG5ekIaPxaiTi/o/NZuTq7W7HtT0/6Zddzyd7Ki0iHthNXtA
o0wI2WRtAxbpJeT+Wq9yxEUYDWuXVWnuX9KO9qKJz5DlGVrzsJIk0nstDVPOiMw7y0caOeUhKSU2
R4zm79C5VRt1+5JjIsFSTrtSdEt+PeTY8KWwy98ipDhervmyS5KQWZHEE7BRcx9HWGoMK80DoVQ4
PHmXLHNVOipgpKRX1gZLcnxidqfktKYHO2nXDwt3xyN3tNQ92l7IQcCOsFiV1IxxFA6yJxa5PgQ9
qEdcsGUTK4Lrrh5LOx4rotGmB9xSCrGrF6hyucoYgl6EwMPDgkINKHpX7vqq6N1vJQ0/jJv1R+mE
NhrhwGrkJ3VfkX9kYZCy9MvNe76pBjYqn11MJB/B/hCDn+5CIliGG/C+RJlyn5W9okibEiTw/ZR9
Mh3d/PHCdgLMy8V+mHsJ/+kxQcydONP4q6ueVs3lzYL9vQ6eXne7frmto1lG8o7LChGuGFF5vXFg
ilElqM/Gzv7I9JB6YuqraAvmWJLA4RbhvWAUBofd8ldZQz1ZqkhWEw8lOg3ioTSSovEAAqRm8Q8u
aDgOYwdqO6HgugFEwDWZX8Mrviroxj1/JMQZSY4qqK/HR5CprPrMhBxx0Ye8j/ZBCEvQ9o/pEow6
7fq8ObeeHZfzzUEkU9IDtNwisjM1nlqCq3b7sMCI+NAUNtaafIHX7H3CLXaBE2b3i8UhSCE29c8A
CMgEjP+3Y4qpuLdSFHO2B0OKgSjHLfZDwAYykjBc/VRxj6BGid473jIChnKv0lun088s0WSNUsXu
ZxqjAzRNaKMC4NmkkkXIHQvj5jZX83VPJ4XN/ck0Yokvg1dH18LXGQdbR+sFxm4ejcvFwn62T0rG
45Q2tSJz+ADoGlaDOKMFWkRcxWPM8jRQP9ljjtfuNJ3xZ4bHB84wvygNKqjkhe4oxc4hg5DciNua
JrLIvjR/bqyf5Zrbw4g+arle5MMWCuiqa13ejr7DKcmdJA+WrGajz0ghAtT46EjO5oLeeEhxBCI4
7Q6e/209qRKFUPfLhqleLQ4Ff0Dem5RqShjU8HMXB6buWydcWghruM4VT/sZwrW1mzuztR5nI7vz
DscAPXXZv8Flvw8ah8xdU5Z3WZVQFS+oI0AXA2k452KPdKDqLVnU7C/TsOVhOGvabstA7z/gFaaX
Yu01qF870p8IZxY7jEW5bG7sLhViNl+8mYdhaW+ZMxnQdNrBBAaynCdSmu4iYF/B7L8Jd1Mq8d36
dG41XHBGpLp14fcFsF7MFsGvXEyn3ISq+/WAaZEA1n9MAc4fhrOwmEKKmWl8958nWdHmw5CZclTI
QE5LYHDSBecfLCuy2t4eEK1wo+Iwx5ngXgaFjG293j4EKkkMx0qPQBVu+zvFsPx0gRB2EdjPk7Um
e3OMfoVrk3OmNzEV6x4C0oGWTmzbLPGSFgxQmDFksfdn6fOxX/fQyCyoIbhsFuBOsmxHG1u00Y8D
iGCpUNSSA4a/9T/frttFhXCpb6EkH/zlEWrp0PQ/hgJ9lY+EOc+v6vHnwgaENNZISq12EOpENoUa
PU8UbzPhmCpRz4A20j+rJ9dbK7zoB4ZNmUFzdtKxNUF0w4gxLtmdZXpVfHEtt1hj/Q3wSpcFDLev
/3XXGwTqQ6ilLG/d/BGEScd4lVB02IPVp6t11TmlfwAS2hWeE/1TNVIbWVKuwcjaWXtmBs5YBaKm
73FGwWENcm/5bpACI1MHL2hOyN9SnIBUqVlssE2XZwodomX8+fQo+P++GGboVOgty9vH34TlR8Wj
vSYty81LBd+FUs8tkxkLMGwUdocbVJvP0K41RZYmZoIigKMN2DFNaLU4DVl+TuhK7HP6ZtwZ7QYK
hKq81YFgOAxQS02nwi/XvYOniEZoZunvsDvHnROKivfarORTQpWdZL1HJyuvg8liaayma86EYSLf
HkYuUUqxfAnad8R89druLh1w+gqGBwbU9HFPgk+s9gcfZ5OWEH0oAOGqmKW+LqzpZXpi8okpTsrP
tm5Ynlq+hdAXYYjuFATHXFu/MI/fNK4q78BzDxkN+Vqo6xLhw0VfoInuDVNZCdO2AB00oZCdHa0a
em50fcE0itVSt8nWGhVUDcqgkUaZWZ8CsDThv8gfbDmd55rNn7tCYBrgGZC6OG/mMgQFfMUoRSdt
ajMUac0GJFj6ld1df0zQCkpYrQamBuAdScIF7kPLOW6oLVUJqxaFmaCRPHXmKkBG+puCHlcgmFiM
0J63KNRY+RuKcoNahvLqAKA6CnTXyWURcX24Z0i55/kU0x4RiIr7N1ItOiBnljw+aTaOGf8WlUPM
QcYq65vZFakR64CCUHa8RNK9GPXdp4eTrzF12Zh6gAAjpO+GQgzs2/t0hMLRuO5wbJJgYIwBcNOo
MVmkv9rFAlgqK3afbJcEmBaaTaVobgKeLvI8u+SYW81oZPrD5SIekXgp6JagLLwcOrKIkf59ozKi
h2OkQ4oAxPFTQb8cXAy/Z5Dqfy3WmriD+KiQ/r/w3w1aMbU8Ilj5aqG0B6RytPn1B3cBG/i1ZxZo
dnfURZPFfxsAukohyglDG/GbBFgC+eD55uJFolle6M4xb62NbD28X/GbXIozFLrButEx1I8HUl8k
53mfHneQZyw40AODJeuDZy+cW+hcmbKQr1LSQsEat2xCsiMxH6W4Mn33ydH/ZhYQyBTiQztHa3qA
wjSVIl+IZBvAt+KyDYBB9wsQEUZ58MbijEtCgmk3T4QEwVX+c07BrwGhYqzPb79xb3XWLvpiSyxw
J7jCHPS0+iXyOcGTCec0blCykEUOwvh0wtLZrwESk/bAxSiMjQMzZIdq2gRLP2NMGFgO2a53ehDr
MVO2rY58O0j3LHkm8dCzypEzRqTkYhp7WLp4+gbplR5DnLhpOXxpNUEAE+uFFfFtiKWDM1qBpD/6
l2vcVeNe1/px5H8oOc4ilgNQCLgaS90N+zYAZ7lmfwInVcrieeCSBXspxJvX0odyZIdJYr6nU0EM
0Wnm0Dl5lsTd6ubjRGhJ/yCvp0p5vi/aavShNM0ukWodNiUHEIE122dviDXejT6163qp3QPnmObI
oOm+bzgxvQlab7UexDkByXxldCJFFEBd90opY1+k/m4/MpAShH0Uxl2jmu4bp6fPqvha66oyuPVj
242E1UsOeI/b/CMnU46e1EZaWIToB02ue5UEIF4LYRdVI7hCa7Nw7bgG4lD7ee8KDPYiWjRh6yIF
0jIwWz7x9kgzz1Ca8BGFe1fWcaOewz+835aP1J21+HdlDVoIlOMXOYbhc1uB5ZOSnRyoe+Hw+uC2
YGa9MutYFFuE2KooF2ahFfQRaa8aECaCAfDpona2cx4FW9sLTTd10ilm4xoD0uOPfGdByr0OePFE
+ASIbohL+S1ICItm5Xd94Hawxl3QGmSBvpkJNESPRG7iQCjYve8blhbc4FlyzadVT4K6sAYq9gsO
MSpVvuwv1x6MlZrWh4iPgMp8McgbYfFUMXc0BcgNXtC94AjsaLwEzpo0abhx9u8uHa0h4Ns4DQ/u
4Z+XGDS+yr1BCT+v3nlb7Jvg3YSbkz3toEXv03QBXob0/HoVQBP1V5hHt4ppkyEQDixaSy0YEEHz
QT3zDXBooEgvn0uqzu2siMxHCBvgnFQ2sDvoa8WTpjp3ohDwO1J0t8zv9C6zHmt6XEJ6adSCsM5Q
X/FrFV5UEw1mv4sTHYvY0FEVs9iis4iDv9elpvsxOz0Kaka5F6nIxFsVQTnmFe3QFwxxxtTz+HPT
B2p9ZPSCke2WGOFy3AVDPxDPfT5lF63FWCB17+6CGZVFARdMae9sT+O4nYuW73dTblrnAIy7ncUU
vFajbR7KsF2TRsew/QXyDkH3230bkdJQIDfKdCivpDSC2z1HmnSexN4VGBe/nJp6PAcLI5H25F1Q
uim6TozSXhyT4mNLvHjQE27spuayiBsV96dN5WBs1WZyOyFToZn31oDyCwaDSKpOK3EVVtjIGYXM
P3SQHXd4TrRX5OqvYcRNREw1cwVjmxMvM9BCqdMo7WVBl5bTWrMhy5IqEzmONT2gitbXgG/ID3OM
2sWgdZ+mmBpYVHIw89FM2WLsToNK7+9XDKdqgy8BigA79cKY4+JASWYuuuLFa+2kmZKkIHzAsnij
jFZnxwFR1dYeRQ6HCebEDX8WoR8mxfLfAbMgY8DF6e2QzhdeycERvdqLMd45f434fkfLTjhm8rLf
8Lx74/JptRJZvNklnB7ImHEaF1KZDfnK/SdvIfetFGHNPjv0eQsNHCG3JHqGgiUTJcPZ+dm5ZYX6
5Q0e2psN0lsyk5L49DtAJDXuLDavjZK/OeUne7UjZi0j5z0HCxyfT2JI1O4lAdXSaGP87IcNxGfJ
MeoylplOtDiMkeuCmw3Wp+aCddd8eOeX607Bs3JPdKAcOoGKmKG/ZqI5xIorHum3V4reisQuTy3L
8UdD8KTx42m7ou5fPQhzRuQdR2AYRMYO8KNTnaHUM4ZsK6K1cG4PntempKh1v8eOPKq9Ti++Vz4e
fxG4Lr7wDkb7SUZBIAywHiTmeNgNwdWl+MFwFjL0Osf2X9+iE3M3vhT4+t38OpWabmvlsBGf6zcL
0AgV8d1j9LBI0UhnmyfumOAyZzYeM3514jlLiGxF9ltAiDQuBmQBS+efqKpZ6IpL0ujeUOoN58MH
HBl8wtFALJS++L7yLXI2OxkjoO+KQ2Ko7aYIAeXRSot9sAp4+eQlmlClabPUMBIQE7A63sV6cw40
0Hc7pCLnkUwZWGub2m71TsH1KCdaRXJ/EGHuzKKx9+XfKJ/u1ZQr8Mr+cQHWzHZK80/V1idZorK8
8uDj3o6giqbm4TizLfy0zKvqmtfaVrUFlfK2RwZeZlfzuZjzIhx7hDCLhFluMWijawc/3Cfck1cW
JwibDTyYrpLRYM8e4iB91gIIB1I3NzM2gxrtpizuxN1+wKTmbhsu7y0gWxV3MYQdJrdSa0HyoGrP
antbEYSlypcNWgp/Bv9kgz4m0FjUZScQOrXrtTZC0EaelA7B4RAzctDklQ06hsJXAaKmrOLOhQMj
lDSVWPUtQymnAve6/xqCA9VJkj+TgSZFmU3mv9ulsoexJ1KU7D+NvqhnEdXN2/SPWl0FBmYtVc4L
KU0VP5NZZNUsz4fRRUh6iJaWDTHwN54K/XIX1jMAG6pI1ZiXb8bRHHFYhn93G109WfDV86CgcK68
JuErDLPGJ/y3XxExSTmwY7fpB73oNOdIJFwMb7t3Zd8hFsUc0fgiBCDwU2rWsCUp0tP5rSAUfxic
qj8qVP/z6yzzjSBSsmn72XMDkwDSRUtHhC+PXVKKrtI8l3xC9XzbTNnlBy5l8ysrIvhXEY7k5avF
V8xKVziih0m6TT4F+BbMnRfrK4/5WsxPf56DKqU3JXE3U2ZU4Wbv9kMFLyLHSGyKqt+/PZiH4Jgy
f+Rap+e3sglRDJFBkhsgkRYr4KHUn7N2YHRzg2u2DxvHdeRX1gMRB7+D7wz+Sxzo26IEr7NXdcEB
pfDotjQDF0j6S53s/dN68idE+OjeAdjYiqE1EH+yMJeRWKjEjeKiAaDftE9Zho7u9JtiHeiIi9dZ
38vE/dIP3igKRaCd0XDWiA1dHjAKo/10g37dYdBHBc8wMsMlHMzBiYfd83Ac8mQp7bIORHNcks+R
RPF86CZizc3n5Tjl1dGeybjFGQXdTJi38CUGw/YUzyRQ8/ezMT5pL7At6r02omsG9UP4dTjkkHHQ
zsbwOXzWxPYWXSdnt1BxxY/fba0fEuvZDscldCpau7KV77wy3oSNYh9hVPw6cKsAd63f5iOAqX2j
WMbx1lc0gLhlVAJuw/R1e28f2ooKuWyXtd9qgoqVW3rAJymwvQZ1o/UzvyjYBR/kYitlI5W50s9M
TJ28ryhUh5X+Q30DeDHSAiA1U0s0rCBY/znv+JoTt+RTQpwxBCClvOT/yBLolgyI7q9lGSTdYqh2
E9oLV0KxBqVwgAP9ilrPP9D7rPdvE8jM76xZJDh8FB9zNsCL4X8DIfJmy0SEDEHN2IdpGany+hD9
uz+jOKmhYVHFO7AWuqfQ+zoqrasXtIWVy5p1MKmXZ+NsXalXcRXkjpeONMAU2/WEFr65LrATTZfk
fR49+LSyqdrH4mh6gkcI/ayzOmkargIZQ1wbTtX03wSsYZfmFgbwb2YRLHaDbKEO4G7KrfeAy7Uc
vyhnENrA+pOgibB8QVDqhYJgDreF8bIkbrl1X1Jmzoo5gBcaFJmjpx4UV9EEeQIWGP95EQI8BIjC
dAy+n13vuUg4CP9b2NBvhmcEDMHpqWIEY6OV3+Pyx5dWxH80unMTgY0FknWeybDMIvM/7n13iGG9
Gb2R8K0a9t5mqSEedagG53LQ05+A4zx7HL1jSQel/cs8OblaDtyeEuyaR814AkjEmaPAgdjB/oKp
x0ASuTuVz+i3Rd/4aIaybMWdiiwYjH2mrK6WT9KczPllyl4AKCQ+QvXQIlpfvApCUW/3EihPus66
Vo6ktWdseLILqbyNEt8vzUbfq/rb2rinN2dKerSyi+WPOwYgbgkPGb/KaTzqQrN1GQiB2EW8zgGW
vFqQK3MQF8SkABE6B80mFHdn0d61VoYardWLJvQz6X6Cof8T+Qr3PNBDIMjF8b7xJ0dSBgMHoUL8
eE1EM5yCRGTDjrNyrM2oThgIKJ1Te4CZF7sPVMBuAOOA+EFmDO0wD7YE/94xSQGP2omJBGHv6+Et
c/v5ViKcE47KXVaiI4amJUijtAH9QN00K38UF3xK+bXxbvK3ApURpEbxNGhB7fw3uYWLVdqhpUsj
jGeWkGQt9W507XwNypwnW+PrHjt7DzlqZbfmRsTaxFc3th/2QIdfy7/MF41KsySLoGrp2ZLhsLR4
woFkFXo8Ws4nEK6xqCb27Fr+ez82JSOSM79iFtNNDkcby1T6ceOxfSDQqr6tC494csgQbcCs9Ir6
mxXaidE8wT6qyCVltLo1mHm7EPC6JKCvo828Yi5ZHxJezdgeO9TAx9SJI4uRBYwLKec/YWpmxl4p
kvOLz+6RnXD0oqcSczG6CUYaxDkJfuTFW44+emU9EOfnautx/GAWFt/mSBqmvMSteerko/Ee80Ov
/hruU/JnjpJ2H4v61Q9r2Fp658iOrZs0PQMiVGsahKDZC7q34mL0DxZmYIeZGPDPE7rnyz3P51Hb
oLqG5KMToQ88sHOmGG0UGkBbFW5FmV1JJHCcr/bK9Owu7AGxt1tcUEwoN9o6uFCDe5813/iMlAvV
6HsZBi45Y1jlL1Ro7xAH+oUuSPafDAXWpc1jeslZb2ITAfCo5tO1ZSZjuqVyf9uQ7Vh8dPUarWZB
JwuBElgvUdhQOlx70MHQwYMZFI6yfD64TTkV2Ek3FU3dNOJEEaLLJ+aot3bj4XUO6Lh0vl9LiJMb
OuwBna+hgEpJDWqTshHLbtURYt3+Kmr/gWVyrvByFPuLPYPZzd12ZvRni9TNyiGUnUP1xoM2LX8c
CAryan6vUSRy6rXRNZaQA+8RNQsxebu6OMRbhxmR/Gk3HfyulY3iyUWhnr7j4rw7KdJsHwLNFkQD
yboH86sUTBumKjlqj+2/qyZ6ZKV1qdSd5CDk2JPP33tOLZ1JbTZvlRul7K9se4SK9a+R/BPGIzs8
zs3xfBEUmXSOFEW5DICMlC/1U6DT5aVRg0gQMDfUUuuJXT1QcZzgDUuEutfq/AnwDdIqPVwvOmV4
FKG/b2NG1fGIbEWmXcQvYkhI0g1rwNcbO55NT+7zDgslVqhwWr30xatIcuqFHDvvmeqt6toaed4N
OJAdzJi8XDmGv8MOuLo6dmN8f4e+a86xxcK3BZ3KTFrUup0dzedCXjMkNmf5YFCJeecwFtCZUops
K1jSMpQt+L66Kji7UvtL8883+YfWstuDVtH4gkhyNZ9O9SHx6VWJm3imA/tcw9oRMKoV1TSpi5Sr
Gsk0Yg/XVf/202FOU3r7dX2r7GJf3/Haun+157xpYlo6ROwGBcGv+HvBqlaU79O6fzkJohb9ew9F
qGxDI5a4j/slvmCXvYJy0j6uqYpjF1rJrIr7eeXQ8vTIkkavFhOc6XbE6cpgBpiebO0tFxjATepF
0hQpEnlpLqth9Sfzol7qP8d4WEYmM90/Gs43F60W6m9iq6bbzYXskgdyIKYKTsn4WwXX/ZFcxrMZ
yC/M0UKQj2tF/r8+4hjMHesB9ufrM95hsa7tgc8rcJsRwUTRhMpiArRVSplTxDv1U59rh6pgN6QJ
UivdbGa8IJSx8ZZiuQSKbqI8MdeGOY1goK3UhjcwAAV8fC0lquD/QyEFJI60E31s/i2fa+AYAxLO
o4tCcwPJyA0tpTdSVLfOoFRsHY5IB9+GrvSQIpFvh/XAnCyJ1pLz2PdzO3M9uLcFwno3POaZgdZ0
WU3Iru5cXcOFmHpR/3dZH8CMfSDG63FWVVrXSU0QLvfPhD+zECN5/hy0Pzm1YmdOuSfqZTl5r4YA
jvOiEU6PBopl6SzZD8I5CNQ2KW9cshxV2BU1CNuH4fS2Vn3fF+oANVMeoHtZGicjQO1fPvKYcHye
vLtzjA2Z+lq5beht6QQ8vzEOMXHEN8ZwNgs3hc3HjG81l4AI8txxbkCZYhiR9NFoAZVf1hL0h41o
EtBEUzakgxULdAedgn5eOeDDexPhjEnerXtnRByUQTRoDNdcM5Gxeir02Wv4bhGWpIidZ0nnkAWN
hw9QsTSnsSIrfDhNGwtUkrfKKUx72Cm+Nnn8izQ/NcS0EcoMXCtEAtn59I7LbC6+4Y5oiHfvUO6k
N4s+MhtR4gd85bfwzC9jrZbUCrmyerPlTodL4Vbny7e2mD69HdyZN6ocqyoDwIYinxHh5/Wxf+XI
82TdN/NIV8iEMqp3j1xDvAluSrXurqHnQjpbaS9pKdShP+AdQXLlzvrFRZNpE+CuO0SqS/i2nQNL
GUIA0RYadaYzMFBaAfVVC5/3rjp5d46OOc5EhXyr3+MkHirh93yD66HjC4aA1UJmf5rt+a/0XUkY
dxSQ3MzK9aBuk0JxzFmGko7ZXo/w6+qzOzhHoeeWLUv9+3+DdhRYQAIjyhHyHaQcM75mwtFs/+9T
rhyUMObBzWUcMZAAwktEWpZwc6+hrjfrgwJ31hb7vHKItPKghJKsPewIxuil/FtspH5KfebHlsId
/p3+5/Zf7QaJ/LJTmHkDz/f0IeSVls32tnYLb0oPrLVe4Mmz5fS+0amS2DhIyqVI/aiTvYtnxXi8
YydRd+48hA/0GJknkFoCekq1BriNeyOxXMNfrFMjiz95vVYrGuayRZUYq/oKB3Gex0nma+Q8f7SL
K9b16HiKEAbTYWC6axJZ8nD6ZXrANceFuDuFJ3+dCBDIFqAh7hho7VEnrS73hl0dmM8EMYJv4ogy
eIzzIftTyLkKGs3Fhd7XIRDGPe2fj5OPsYoFyDoLFb1lkFw75Dhwhro+vl0//Gwcv1BsILMgvmis
zYp1zctg/KlDGMF0WpMBMw8px7DMsB5WptZCSnex2GrX0IpyHumt6+3GgMg5RuIPYjmRNyiEXccV
LczCMWesJLcxLnDIO/v/dPXucH+RzaPzWjGFlthdsFaAKWGgUCV6bvNAima+/GjvIxs6lmG3xH5/
YclUYdDDQ3nPOdNslUbm18JruxMstLhjgxvd6SmHUVR8/9ntJSBce5+exZiB7HU1RORs8+5wpWON
TuuCBpJma6R58CytLyPhCvwQ277Xyvd/EhhC8NhNCotjejkv99BywcEtyTGquat8XkMsnnjw6QGb
DzCuq7JL3T/32DYvplc+Raw+ruc1e3jjMm0EbIXJZF3DSdm4idZDZraW3rrrxlckWFgegb4Wbxwk
Cig5jyCx7dFxKTWayZBXGCP6hb/YRICwrTG5pmsNE9cJjkLz3BmkJXXOISvB3pkeikuGQU+6fVR8
SDnCQ4Q5aoVc0MiEnTKkqAbP3oLmwKTGFstIjmbeeGV1QfEYrx9l33tdBpLIIlXmTZREoOvVa1Bc
B4OYmh/isQWibu1n3IaOVkPWZjhcPdQICGJALKlYLMbO1kPoIowITgf0zmGQltfL3rAdR+NAJSko
7pc4I1iZ1kxJbXEhhq2+EKR6VQ7LYToQgMi8ZnwZXTVhrzA4A9mkfGOLoZAq2fGca19SnCaIjIop
GlvBbScA0LfRZ8y/iX44mXepkyrAYhIbRB9EfYgnTV11RSgob5aNip2x3RLHwTGVqwHxqD79X26C
aAvZAbpLGDuAt4W4fYHUTZ4UQ5P/saNcKfL+JVTXMYGdt7mFeqI+VIcFxPYu7Ogp5AfVT3w8NTAM
k12vMFoSZSNVm19/TlXW+XHRcgCosoyCtCKsHIL0yOolEsiB/d0TYjddqNrUYlubGg0B9FlWmTGl
IyA6Vjr5lyBYTW0oRLFxNFtUqxgUEklgLrDQamY0RA6ZiOAkgTS7vPumOte4iVgUNJqX6MLgQciA
Vwjiw/h5eZUdnvmwF1AvOfHJYm5UbrMzoCyLBwbHwTJ+ExdD//BMWkfHv5FVSnCPdGpzfUYC9cyY
DW0HWxyQHofYEqPCdb4EqnX7YKVZUAkh9lQ5SZEtGE7jyG+ovAQ909DxUGkw759aXe1vPtqeIKHr
FwbFM0xos8Usvi2UAxmDznySBJlibgKkKZt60qbjcawwByMSVPYIkpd12SsSic1f/R3/gUarK4Av
9QWbd/4Wi45JCNtYMP+GALHVuafnD4ZeU9/Q6xS7aBBp9S3OUyAAfsVmEPGFDjt3+7WoB35Pg1Vf
EQUY05pB0isgM6XC1DItHwGxbsJCucZiPk92OUWzY4C6XWruWhKD3Wu3iRqHxVA7bBJ+lv6RO+IC
CdHWlkK5NK9mIPXXBjORbqM/Cd/q0+oF8qZS4tdGVoawuCrjaO/sj1wPLBOFBbZDq4Mej7Pt8gpx
Dhu6hpUHfs0DWCwK627wl9o09ziqwfGMUZSjWgTztKuCDm1bOpETm+qCXHCbKkDQrtNaMBoQHcNj
DLrVX0cSr/R+jKrBlTjRbQnnyGBm44tYbR4EszL7Yl1DDvOfxUawvhN/SEfCsTHtynJPOtVxRTdl
laaVzDGY9am3IzLQI0shMkRBP10GhRpPLDqwvBNECkcsxydQA/pA1A7+SwYsJkVDcjwwbo7PHWul
4UKE1//yFnca9Slp2Q0Id3DHqYabp18fQw/+I8hXy1CVMRiWWapWrp2cNjyS09rGvxrZFeiihVnC
0P91mOR1sHJR/tWmBatPxWiepfEgacxWfS9QoHQwSVYdCg60cJEpDPj62C4Ebb+GYSBsZlZtl30B
CllTlxwx7P2ApkfZZpJmkDInU8On57e9C0ClgobzPvZZ6H+1RFAx2qKC6nmpmONHxtfr3PFEnxKI
r9YL5an/hxlJj931FoVtXK1vEFxBGy1IKzk+n6QO0AaGcBcbc+mSZAkt/yj4Odl/pKUvgLd65hUA
sP8hktlrXGl4Xu2rxJqzhnrqXaxQScEQwb8grfgAL7uERnYrP4NbRsMpovWPfQwSKMLqJ4RO7r4S
Z8b++y2RVquDK119XJExN/qI1gBLknRdcimP8jF0+ODbeG25QmtfUkjLRcZC+iXRwyy7PSl36tyb
HTbr3mHo5YF+2TalCu4o3y8pgumj9j3xd4FMBmvqPxklz3TjEDfiOhtyBJ7tZgXv78XhSkhxH8gE
ilhW06/3CBoF1uvafNmOlz48tVrYszhOcQw/mzBj2eSbZajbBx2HwWY0cWTdr546STHuMJNFqsTU
IBiW6uPqm/5taN8URgAMy9UbBWL/AJac/Tg9K+ZfDTICy8Rgrh6U3F0ndq5iNl2Md7ChslvV7kiA
Q2+6v+H+uFprET6oR9Sy4MXrqz2SuD/vhIkguzkQJk/DQFQPF0c/y+Lqk0+oo1kH1QbZB+KffSsp
PK4aJ4e9DH0MB0OCYfolLKO0DCwk/Vkfv4C17D0tI+hbBYl/ctmq71UB6AcQjghQmUOR7fUDKap2
q+L1pFf8ppDxElaneWbLX1U26BINlHHDqd9RsdaanUthUTNqNiI2E0fkalWBo6Drm0BZ6olNQeBq
1AmcxSRjDWf1HYgX8EC0LWkdaDguH6e8NTk1p6knjl3snHiNoPE+IaO/pUUZQiFMXLvftB0AhBF4
8JRCcKY1dbq+qOLCAuIMYcSUjuVCVqZPMwZwPORKlc74TdHgTInZBsSYE16/JBaqSNMAh6gAoe31
pvcjkY2htlfbm7lU++P1Gg5aB+MTCXMnczO2KxORanOgQ7bc/T+TTOgrqtdw3EfPotaZJuDyCD6L
NCBNikFSucYC3NzxEwJHnQTr7Cz5GedF//pBVSV/FS5391XM8UR4ehE/CjH0QxrAdEn8UJJWcf7n
6Lz+dGF9hbAupH1Re8Ra7+lQQwWBEzleIyLCfJs3HF3leBuLKo/vhpYakw89jFFpdk3QGD12/gh7
xQ6e9eNB/ohqf7610QVDN8ffJmjv5IadFiyRutUclHOm9mjdN0qUl3DBEdBP1858AVtPM3u0Ey9L
ycPT657QWtjF6ixtk0kiv1YBO5CI0L2rylHvv05fTvwZPUxCslXb41MsnsO5yyn2rmNTt15FI4nI
U84gQp7e8aUTY9M4ecjST4k8PTVyYtalY0BZAlbd26sFNTjHPIzwqZ5OUQ6FlMhB640pGZ1lmIJd
DlbSu8gQPlI4HjSAZfK79+EhzoQbdnDY4vjyjLEBuqIFNDjCW7fJ+kRFv5lnn5ajahdy1xjX2XFV
L5VkW+7/2Hrh9qeiALjoveNxhTQQRpk0K4NQWIid5VS3gTghpcmmKpTtzTPMMMCcU2qXuzoGlKCk
qPjr0RW6vzqv1ANqTBZLXWV4MnlWFWbFS4KL0HIkA9wYZPsZBTVV45mPCelQ0ZmAQ+UXzi+xdbql
yogOl48/q/cA+WkkAOtdpeANG0B3Dp5/wIHxsCiBp4ybhGRuREuwAJSt4NQUWu/72ccNJDYSbt9X
zl0X/l5n74/f3DOM4Qbmix3HgLUx7sM2vnYDqufBEL5eIgLwmumoUpFMZAWVDc9VLqEMOjXdS0gE
YinzzqEIvDWnyOcjD6nP1kx8YACSRX+6oHjM9zYnzjnr58sriYU848GsuS/G7sVVqcMDEjyLy0oF
/5q+WODd2zVxOy833Mi+nKAoRxTl4TPnOTNhLX+dwaRY7M1CkmWNBGxZSW+KuUu+uvewn+e55sHc
mgKpkaJfTG3YHqgBMqsEE0jRjSq5F8J6lXCG9Nmf07VYzBATr2GRdMejg2z3WJBwKEJtAMGJ1KQ8
v41hVUbSxwjH6TUVSbC+KvdX55qoeI3nUB5chZOSJEe/c5tGwVM3I5TjrtfmeUlhLssDHyNUvCon
BdetgzicJDgYeQ7u9RTZGU7F+i96r+hu5jLybIWj/RC9rTEmylwmKSPwuhC4/5+i6Jcv1m1Xeqqo
x7+aN9qjZgx8RG7tNy+pSB+qIUcLnjs88eTJljtGYniaxFb2Ibe8AGV1S/GOVvZvYCOLtlH68sBN
1FRWHiXMDOh+rBDIRwE5/MUVqe2QMlyTx1RENZ1hRouHrEVUkl7ZgJSIKUe0xEId++qVxDntNRWJ
9DCDS9hz9Hm5gwkYB9NicRM4YQwZqqai9ekun3iAI7bFNDyxd+brycDPKx6ErPFoeKQvIDTUyBvs
i4AHxTqK4kgL1pdpZ91qNwIxxC8P7Yv38noteYFLfk9gcOPNryeuNlRpYfKw5AGf1UIi+9DE6xli
qvQaBzI60+RoPzp4PcewXQfAfCknuCP4WDWzz4tPjo6WLtEqH29FXtXagItxsbsBxgG1HBLqy3U/
R+jCqskgb3TVo0xqSnnrQQijvgtPxsyYf9AUw+XQbiVV7yGikOYIIKAWLTr6B4i8y+dYaT1nHRTw
NHIM1Prv+EmX0+btq1nok0OWQx4ocZseeDnctT1wNLnstnqpcsIfPnsP6qiaRmO3LY/ZECvZ4qLP
Ej17ea2inFXN0vUe6PL1PIxriwr2lnriufcFPUFW0O0Dl94nzWTGM8TIhhnvBjF/QCj/gxFgnwfc
702Y9R8WUFml3G7XP/dLbFFCvuw6oN+VA+uArt8ALL3ojOf3a1ksJOYYbHPclUqdduGTlR5Mm8hk
J2HzelniLvmbOC/ndWDXcqNl0e4arJ5AmByp8AG5LRn5EXyIV+vbjyYgeXVv6u6qhs2CkzpUBvst
fjBLtSF2M5KtAGLjtgS+RN+Iy09nQkE7BZoC8oZr+SMdwbcT+QOlPFP9e271lN/VBjMkLmosR78J
uEtzkHyk6AEj0DJOwmaqjCYBkn0dRpXfrZQoXvdxr1mcmwwefaw0XEixrStZrTbe2c6Tv6K33z7U
iVdO6sKPN/s3WSrlTCIyhOmICRBV7nS+ESwnY1gDPegLpg+XG9QZ8HuenHPjBkmBlkU1/YEOgI4f
CGwQXJIWVPjIqR3x6WsyCtLb3r97SEzPJtavMm9bIPl5wxueNHGCUD94yIDGtrezAdqbr5ZQZCaM
SebBuljNoHLgoEVKplN4AH3b4EFUWjbhIx4K33B0xfcSj1gkFgKESDmAsAimTnmEevLwK6NuDa5i
mZX7cvMFqePy9AL0EeSfrZQTbS6Geixdvna5g/Z4r4fajOrDpQAMDM7uBySE5OYMigrqr+uDVRwL
HE61kXtGYmo2yW5SpVPluqn8n6EmM6L9cBxc/RqSJ3vJoVf4z+/ZftG6kM/xcs6zbG+6ryrXOTDU
raePG8wxvhxEnyGRFPnuCGfNJbDqYwufUSVCChiRqrjSBwST6+Hdw9R/JZvnsypOXzqk5GCIr6XP
o9u3qUqfvUSEfRvqcg0Mj6PtnyabTfglA7ATQ4iTNbss2+pcss0TgCAuhKazbwDtgcgPGZtCJHZc
eAF9hB2BafDpCIOMre/R/jrB5w264Un8b6IZ5ZsHPs7jfWQp44fNbdOA7YJaNuPNCiQde9R4u1I4
EcRu+72Eep7xQJSo9UWTbJv70bvP7vsmsoDpH5ncKYc1529AyrYtAJS5AcFtLk30Pmptsdh8Y8Sv
nsiDRUmP9j3x1YXTdstOmrodLXw0D5f3AmPNPQ6EZScio3mGh6ooOB5Ry0BpI5U6AxPGZ2jkKrLW
QhiLyA0oCR77vj78peYNxOVDfq6RME9+Ndyoz1gbf/x6K0OPbpYrJRFalS6b1yunvAYgQ8hOnTYv
Z40LMiT/HqvfeHL7ksFkvObLrwR8JJdJwOyu0X/BvFwX0UlUASygyK+0V2jhx5QeQ5l9e/ArgXNW
aLls8F9yTFVI65tKuF8LC+bM2i81iybvXMLGhL3tVosQBzunJBnzzEZTil6xG555/3I+6CxT3SVR
aQ9ZIkKTG73hau3bjX4WA/fstotJ8Imlo410/kj4Z0d020xXtzuz9+dmI3p8sljXahqvgYASGbxj
3tVjQJLQ4pGuEEQcKNf2K9lLss0cZy2xJln03OA7Fa8TWtfpanTfMzj2toaMMYucprgT4P/PnnU4
Hb1QQniDDkYxPEZC35ojtyOh8bDmmoQkyuhdvLJ4CQvh2Q5ny0FVT98Q6nNLb1o4nGXp1KoEJmEH
EzyW49gnBfOI+FUIbX221cwCDaQAPFY67Y9xvynr0NZwWHYmQOR6pjfMQ/3dSea9w1G+oJSYvQFI
X5Pfsrh2Oyw8IZ9yhZsMFnzNcsCYaHAt0ROv4FCLnDAp39i8nJPVqEmIPIsVZyxkszxQCkR9+37g
VMKy8QHO44pw8ArKYsJNvxtlNdZdDDJ0jJa7ReIDvc2S/6fIiYLcAn5NcOmOcxewNrr3Wseovm0Q
lNE2ykJ/lAhWJDZkTxVeLR+950KtJVcGLRpT3PUNFk5dau6TSgO48sUQ0Lr5VGPZO2fhxkjBrVsz
2I6L6VcH0/V4kNeoE/YbjAdLJeT6+5uyw216QaQ6qxZ23Z3C8tFe5aru3ccWUAXFuJUluR70z3lz
l5SddgDLz1zVeP5d0LsZS1aiJ8vw+di6jR94Wi+pNEb18iBkhjieWk4l+UdwbIBeymIPxjfNjzwf
0cF6JVcogURcQyfv5x9PJq1WtA0FiOexIOIxN4fFDNXy0hjINTUNVMo6WYtIOcHW3piEc8uywdrv
vGSvpo2yv9nCPRszm0nae6sc8rxYawn2OXxGD7SYMdCn7x7Ca6RkzjPYWvNv0/N5KWxl2WYLYAex
UULsJSZ3WUVH7E860KoNeJW4ddgFKmuHlyGa9+4lBGhcYEBmN3YCb0HFQr3beornKaAg1zmZHK/f
k9vaCUYDd0xoxNkgtfeP3QwAF9wrTmuQI6B/nEa4Ax16Y+6FRM9QYEFoyHfnH4RDb6mmjy0ajZgN
+F2WetdPyrBqDWKIljskEtgJwzmp4rOkw67JRdmSsOk6eVgbN4TLjPtXBYz8ixH/4RvnTnnBJ4ND
hRGj9TAoeZufAP9wAh+P86IB54UJgz691NaAq9vJR04SClaT2V3AC6RcZkACcBkf/WS5eGY8NT12
qXeTzM27YF14/FGG//MlkWPUezStCHaHQ3EfgcQSpRL1Qeyzw4VkGwDUOujiqlCXJnQ+rydLmGlK
fVHPxe8PMiYeNMQ4PbOo9MOIRI2vGkpcw4d7SpyaUlNjhHZ0wzCzMlm45a0rcX3bG7KwZyrQEvsh
0WXrwv3aq1vicfF72K6zwBZFnkIzoAUYxugZrMaHJdhubd1Yxx0bQDrNpFmmO1EAGmYDxnBuftYW
qN2fra0EQI3b/OOn1bEy2jyWm5yzS8tN2iqUzOhd8eiw0YaOXs65artR2YCucpS716BWyf9NtfYm
RfZx4CB2fC2f9CLXax5YmR5yq4oyIunfFMTfbl24bumeGhe4NazXK62xzfS0m4yreOtfPSqIf0fT
sOvuu4681G9jsoT9GFhKVOD1d4YzEzV8cemfEZBWG5Itfx7XpZ4UoU0gheCrMwqfl567yNK+JBuD
Ld5ILse23dgK/bIhPCWMH/wVRke15ZaOTu+CvjU0Xh9hO4By8sML/vVOTxUWXYNB7id8n7OSyMVn
+B5YNkuVhgABkmLavNPRq0E59qiAsTkqOcz7S+NTTWUCAj1WP5x3Xz8eSmCSWS0fy5tvpvt+T8jh
byv9WVzkBXY3pfqYsoVgI2KaAkPn2CUwBhu1foC1hdbSMMYiu3dMHegqaZM6hAycNeh6qDvRzx0y
1BjhsRHZ//Tdn1uoj26ysE29UrW4KebYphfSK2ysXQB6d/xKpJHtW4lca3OagMx/ezN5QJZVInuz
5s7tcJIxZaOIM/v4mcadl2GbIs2k//qqjF72Xpn4IM4pfatN09QHB0CXBQaDdmeCul3wxVsFBR9S
Tnbs+7s7LW0b9oyMGW2PlNXUVSDzPBiq7gNSkvT9gOdkvoHF8a88MbM73JkheuHVmQnHHM7e+PbD
zFOdFabVrHiVXsYuM4xr0LNltL+XzWBY3foyyZBaQLLA0wUA5Lo1myF5rkbDIV2ioY7SsBvYWuAH
8MUEEmOHXbCnqDL63imRrtYB0Fsl4qXVH5Z2wmIV4j4bWP48pZL8anG1fWfXb4fHQLPIU/SmLHzs
zKP/W1T9BGdWMSlLjgeScJGkdXHMLptue92sQpZeBm8+UiZHdL+OXO8ES4Ra5C++nJsPL/kDb+hK
rUT0FD1s/5qmwZd2T+/3GmJWlGQndJtXwZ2j+00j144iP9j2n2p93wRqZqoBHnjlwRVQd++lv21X
jbEQZ8EBHQL3VtgHvHM7LDZ6VOp7q3jZgue4QmP2KX38ZEO9wzy0a8g/hb1RWK0WOpuDu4UfJ+9x
6OR5ezJgn7t1fHj1ok3IAN3yXfdcsbaZmKIbqBykQUdDXiDONfvbIMct5JkXA8wJ1ARFtm98wbpq
Nzg6wJ8Ivm6UWSxxyhCPzh4jchLW67CDKtVdKyxqS3cqBlQctqpnJTqSSlSUkwXLaFA7kFu5ArdV
7B69YIKp5UD5mFkzTz1168qFaNARh1q+JwYmHdkDz6u94y9BGdaVE6GCY1FkHwaJGqW+0Nky9eBz
sJfamiCjNkbswBYqcpe6IYwu+nWBDonUTErEr+l/zrPxd91y43ZZ+5R9Sb74DI5Hb42NDt8cIPu4
3CKedEYy1zXEn/vZisbp+qpJtQt5zgIwWiTJoGh79wsyf8hhIKA2jRQMblHpHILeibddxUyIbMrx
TQWWcpBunox7mJzU8U+W/X+36QtwodIwkQ0bQaSaapPWdRkI8RwxNEVrQmw3vf51s1nywGDxDp5S
JGI+CTxzNRe+/Yqljq9jCsgXwv2sye7N6+1CeT+rwVgopxqdwbAkaco7DaSUC4qoaK/igubeZNpX
Yqv9GYW6jyiTeLT7XMoDS+lg171L3GgoBtfaF1QAbbzXbuoF5CtLDPUT9TWCokpb2M+HQDjlwj/S
ALoHxd3fB6Pj/E1qGRhrq4BLtOvol9AYxJS1UYxoZdWZQ9p1qCAcPAD0Mbgle5gnyVZvaLF4qXLz
w0FXyLJlN5RL1vq/fYwKc3fTc36ZWrLwfIHqVfwNmHhyoZXiYoM4UP8CC42WieC571C3xHmgxedP
62Ewl13YoNZVgKl42ijboRWxqvtGbqgCZNmnboULWEnsxAaqh+Bf815oUU8mrgwGMBolns38O6PI
bHTu16VgYhpVzaOpPlhLN2EvIFRquqpLbzqmMkJWWSB1thjhM0AGyOLS7+i8yxQ7sjmMJLJMfWkr
AzEg0+zYBnKg3aCLicyJ3qh4rIIrhRWSHEKvy9fAz0xUgDPdaxtY89erL1zb1k9o7w6sN/NIGX28
9iS3B6X/WCGvS1rj1afm7+ZcXHAk8i0wyvLI2iQO0wo6blWqtcWddX6r4dK7eBDdxtufAXqNzU/w
EAWdDNhdvqqWxDCTUO7NTineFjs+t5SzoyfiXNiQhyOFgX5+XPBFInclYs71XtPwn/0059DYkLTZ
Ua0ie+nkgjRaqCYUti50gLZvdecHa93H4INeq6Kkp+09dcPP8iwalhOeiomYRGAXCvewZwzx3+WO
Hq+xlitqf64ylAU87olrKonbt/cHiuxS6I+C7MiB6rD77osroGG9KvzmqRTc/qOFJqLRMDJ/g8B/
DZcQrWeoFCWzfmX79W2+XzgHfIWVcGvkHklZihGnSpe3npxEpWseQD6U8ZGYvFro9pQTwkUEbOeY
IhdTZjiuf+qoi2t5f84jLzw60Ct0mLQHRxb+6Nya+3gj+bnr3PHiDnDXlL1LhZiU32VZ4EWuhsYz
Of9SEPWlMMeX8lYDmED7v1OP6BZ4vth+iPwqtISuk7RNjgpNO8JOfFLA7PPZ5AO5aimqiWT1c2nR
2h5A/yX5r40u0TPKsG18bgNfzDOQsFV0ZGMPs/FYJGk3PcBkiLs2SCkC/oNVtTcyhG3X7zqOfEw+
9SN9V8YRMc2DKt5pHF144KcFcRBVk2kYM3qOraX+wiqOMTSR+2YqdGi+g3qEu0/CsW4Gj1BDmimf
qXV5Hdu0V10ENrI7wKHfZ95K2J47clhi4odwv8YkQAI2IksJamONePK02iM29V0RnEMRmLbCQdx+
CjqXl1yXwyvJNn5ET8qiAoK/YmNVSwJJBnBjnDXreIqBuStej5yPv69IrcyzWsQKqb4Yp9i7HjTd
0W7NWy/La5Zw0QlFC2DV1mbyMep79nR/IEF8PI2cfnk51O21CBLs0qvAgmRzXmDKJZBxf6jYhGWb
a5QJCxjDUoBx+5kLqD35VNyIFXY0rRe3Vr5oGQBQrmDQiRv/fYpu2d0Mlp4P3LrtHGsF8oWxkugY
buK38ZBIM9e5rwIo0objuhMC73Feyry4JsP9IKW2vbw20p8stkuy0Tg+ezoxOBqR0ltHGUqZISKm
OoawiBlnNrzEXRQJubW/KsR8WOmA+Sk91hOQO5iR6dhB0NNy+FEpWySBFcKf2TCb7kk/NFhzGw3v
60t9vDxDHFwLm04nvqcNIMZ2pwj/5NotBUN+UEv9NZyidFZout86i/1ODktsq0691Cob1dLEReEg
zLLI+OOYCJIr9AZZMu3SXKK/f937t3M04tl+XKtIrjb8/NnBLWdSCwrvTFXHllbsv4QouryyCukT
iF48go18okQEjyLzyi3vHAdH0pjRf4DUYrU/regwgZyXLpU8LrTrvlyH9uX965QbFzYCBpCQSvSi
FKyC22z0Hd1IXJbkaDpSTGsoDS4iNqu75+O1MWoWpXOWxSz4XP5KCYLfGOBsoQ65w6wx/k4WMh4z
BFyANHVktXw/1MwqLexHnrfm8VJ7rXw45VHjbJoyyh7hNUBWbzquC76Q7PSYVnoHPcE6g4UsS+ci
9m/OiWsT2vCqzvW9rzdSe2yxnqm1EbVsGhuuAoB9gv1nSxYNz6DR7XeplXsEmDKmnD9W7m6l7msy
Ypl6ERHB1y4NkEybPqJnB0KWrwhGDX9aPt9uKVRiZSlOMOeWjT4E3xIJA79v9ABdurRwqtiAGYvQ
EzlWlJtXZANwgF/mU2LSd39YhuVDxZ+SkJhS0RYb9w20N4fyMkv4GbbclqqbmmB8ICsKQ9befl2t
Zjz0eZuK6YT/YRWFNUDxI3LfaiTQbem3qTCKpY1+bNikbTPjdHqAZJIZEHgyIkRe0ip5P9o+JQ6p
pa/+D4fnxvxSJW0fW+w4z3B9lpaOvxdRHWUWCcgqnhEfg7UQqmYQlBBY2wcnIhxLU4DgjVO9WMhK
Pvo+qMqWeuqtvUbzppIPdU5HvRrggYCS+7+daG626NZrRr5y8IRRF1xRbsJkk/lwENbEsaIfzoJC
c4KNsUp96BC32WO+yrS0FcWu6O49tC+5AIkY/+eJ590nMk3fGc3VLnlVAqG6Rgz0zKAUInl+aNbP
qFkeUnlF4tLHDUZrU7//baFNbou2xLecKRlB1whEYuj/1x2hmWVcGtIhiBVv6ROtJ6MUgiVGnuoR
Ww0MU/LHwAx5qrpVpzBjhk2VEscMopoK7xi6bNWK/4ID/PcyMCqjN3zK4m4aNBiNSt3at9YyyzxT
smsU6lUmi0QwwxM6w4cDFQFoHW5S7IrWHOFAEppGDn4V2Vo0fS2jS9zD0n+IOknc3gEttsz+kG9U
xAv8NgzCP4Lwnh0HdSkGqvWNC3goYSC80gEwDlk+hbq6Z/GguyQhcgxncV8xKyAEZk0LQtC7S1Xi
PlbkqKql25ILUaDJUzQM80J3QIMzjFihpa5cN9lhlVsGyCrNNGwJC/wSr7gccvpTkHpTgOdjhvn6
YKVTN6QpVJg+Eje+GXtptSW5obzGCotEZd5IdNNY3Em3es40xsOArIH6MQNUqzUwJglZF/cuEb7b
2s/InAIBesahMYCXJZP3i13qjFxmmQ8DHxT22A0BLhWizSSazGJWxtfMJBHhj0pneWKL4G2BiYZk
i/ag5ckUIEQqJqWhqukCM7OdV2twLrjc9nPHCid+utMoonfVJ2z2DdbzjWJdSlEJ0+RCOgqGQtQL
90/T0B+14gTlgaifJDaafejV+roxsbh45S81EmmYT0gPRzqi+4kAvU725DuyHHo7/RLAUPO5lja7
ubDXc+mvaoIZOqfhydQz4JR8KuzE2ca/x6byjbMYH95Qzh2FTwTJf1GXxQNdrPib6drJqGV3bHbp
UOsrCzy+rgGz2lDjQcv5eHvT6QCXjTIxjO4ILlLmoAL9m+QdjAodgqE1LeDY9cCjpYpRjLPWgnTP
kVbn6okbDM3Dsp4nxN6kzUzaK4QRvYaOQ6vx4Sg5GjR12TSgeUAyM1dBkR1IkRDX63qjWh80djgp
HSKLXaP/GJ88LL+upAOfmG0mRodxakdM2f2LfcdX662kCHh2tZQMZmOjUaR65vWxDb+lzVOmh2A3
ekTn8VKmW4KTVW2lI0Li/Dg9ohIpmesfcP7Cv0ZxB8+RDdan6zow2eOMcF61XF04LVCO3Sj2zXf8
AT1PUELcoQGOnA2qFEZ1As1X9APbY8BrC411xVI7vOrXH4l3SmgoihgyUXtofMeLjgKawwkRV1hZ
v/iBUvSkv3g86D+x76sTcyAfozwPYAiPVTfIUk2bye7vHdY8fkY67GZCyJbtIX5249jN7mhk3qo3
77TT2IBSBEFfVsQ7L8KkcegCgQXF2OO2UyDLbL2T3hJe/Jowj+y/DmZ2lhdc17mQZd3VpJnqjiyd
pmYYw+enLkuXvuPW4y5ZNBfrSgIGjrYs7ktJuUFXcmnX/dERiG1Y0OxLPiJwU/alR8J0tQukTJtR
lD7Jh+CBJu0hB+qwIKlgKizFQk+FXuKDvFJqCyX9AsWTK1lEFGp/BVUfpKbPDBgXdGlvcDNykYQm
ODyzT83dd/V9s59fixTL4HtlIwqDtzns+XK7D5MmiZnMSc7V8lk7+m7m7jkQ977ppSv8kIyumLE+
hnlWmBHQRkyPtcJwiRicPo1jLyQaRiEYU0sLVWhySzeBd/5mbC6JaJkzu5WBZ7k2p7d7mZxEstT0
KhkabaC0DputCDrMkA5zhBj/thkFUub43m/aIVK96qFOZk6wYsn6hNlfskeKcbE05zULgk35TjAj
63t5Epfk3GvCldRpvWTuBPxjzvkim+hU2M4b2T9yy44vjZF6JoXbSTBIxUoTTX6DE8AMBpjam7yS
wEfBJ71WXUpYAA2A8pi9axhJSDZLSMOuhPeerNejH9kNo64J2rCTgb1EJn7sEfAqJxg8r34SY4YS
JKNChZYCqIv/ALrmbb3qlZ38KsXXFPUUS6TzLOvKPMurSW8hUhawcD1F29hLvzca9BvcmoQIfi5b
lFNG9unNOVDCJ6wo4iQ+uJ6StvY5Ze+KcuhknXZVqJP6K+eEpZsYU/yv4Ns1cKdY5LQY4nG3uPOw
CmH0V02MxdyBlvxvnWgeYorUpERG98bG8ElqGemVIKHICCvgix3dBa5Q+Hqe2sMjkaCU8v0k1MG3
5RofxTZcvzdIDVaIhS8y9y+oM6+sfK1aSKo3jRml5ADUhwfUhG4Cr2qYcyC+ro1tvGY9coMnAGNx
nTjuxjesSxO8vDtFCNhhAtA+K1iGdZXVuZDEIQ5g1Ab48xljaEk1RST1MlsXAEgSdbZrpn01pucE
dxK3pi6DPkyfXL6f1pOATujJdNpGYjWU4ZriHtgO5jAcdqSltb4w7DP7MRagffazJADnmt5DH+Gj
aPqtNO0MUHJb7NY29d2E8exlHhxejvumgzNBkb5EwPlzmgSObrAF/b8Lr6//fc+s2NzEwUCdoS1/
zdlzL5LjhwKorr7ChflP4Jk4SOEz9JlLe9aMnpqUQO/xlxZa9UdfeBIb57D8FS2jp4GL4KptTRaa
I4y1jd+/S+8riKlXOYkWfhICkARIG5TIcTAni+fLOOMpslWojDrzcg44CIJRPQbzVYKpoGpQdF/3
Wy3RkFr16a4ypqz4rg2CqlV3CSJiEO66QcAp+I/e/dlawTK3P6eD0RWjkvv8tWtaZeezvmHJH2P8
9iQCZZOEYF47jld8Qp9NFMXXMvDd8wnp2WEWrBH6xajD1/Y0UmpmnZ6cRh/6sdM7bkUjQs1xfFZg
dq9x17DTztz3eXg9quFLW2Lqn4RnvnRLS2QHGzSEXG04ozBeZiEUYCUmcLdkz31KPW4On8Sv0Tcv
GFw0XigVfaKjiYHN0x/wTMWxDkgIRjBmAPR6lfkFEqOfCADoFK3RffUX0Fp2UZkiWLXHfNOY5ufk
kHHh0CCZBH7enr/y2Z9TuYGbcoWVRBGqvGZLqvwF3U46vqW21lvUBTBVDSbM5sm+5PEAswqa9CYN
JoShTSz8aJgmIgEktZPfHMC5VVa8eKTj4lfBDjLclfwg28X3ZNVY+NbxrvQMIpDHlvpn0i06rNMn
0+HgbaHs1AEawVCWzNSwFkTDtZj4STwbI5Rjs47zAKjOmK+isvh91goCJNzZWf0skbGSNepeq3jI
U0cbwkcI5ArdJg6jGPgKEnsmPbH6o7bxUaQh7/v1gA+qAgz/Z7Pt6fvqMIQ4EhHH1Q2boTIC04Zd
WYmqr3D+XbtjpAkaWl1sskkTFp7XliaBNBrpxBIe+MgiCJljlOldnyNo9hBM2HZQc9O8y1LnVz6m
NH1+c4Spk1ATZe5CpdWyP43HnN5ewT/lfOJ5Fe4doUgQ9y1LxK/Frpwx1EQC8bmU9IrnWFNFANa/
Glt7/C2eN3rBlw8GYzN8VM1eyBQhcv+22MjaA2LrNfd6X/RNShIzV4gf3E1p5RsSHYwX/Zz9en05
iJYzSMFanNpprVRMc+Zp2cyWVf2YyIKJbIvjDN2/qeSiKQtbu/+hHenFMqpA0vDC+25XbQCqqfGA
46l9tBNb5IAviy/3hYf3PnyP6phjbDOUbFCweCAUnctL9/KTjXtwpXw+5gIQFIKLYapFz3riYGaW
s52rm7Q0nOoTROt4IePeJOwOzMVyn4dKSnGnrR2tPmnniO/aAAdy9I8RjRQut1l4pbEqO6rCQQDH
l0eEoNslmo3gLWZfe2kUNhhkVk13loa1Q3aR5Jq/RXy2GBZ4mnZqAjOBc4qeXS4IFBOLibNgWfzq
DwG3Bdfm+IJPrlefC3UVRI9wfmXLpRb34SOBKFGjpo/eiOwLpamb65nlq8vnqVRVPrNuol9E8LrF
ICQBDHxtpACaUY53xkLAG3YGOK6s2zygn+wqxzT1Hmk1N8dpsjoLSt1RnPdp9SSfo+f3akpXpflg
IV6r/T+JeKPfuMGyu5xd61M0+ti3tqnWbGGPxWGx7WCKHAReeRs3HTiSjRepURK/ND8uQ16zvT+F
XrYdy7uGL4ptXNy7wn8Wns9z9CEMt39VkD9xXkvKN4svW0LhNQ82A9ahhiTd/jgDsdAnJTsIprSU
83Axy2Mh/CjTgceQp27NDn1q3833oxED1Loa2p45kUUYgWQtYMWl/RpcZcTxq2KQISAz/PXf/En8
ThheCGfwqIka7x9HZQQlNudjRUH6r73AHWOhgVe8werThaGVNCgOX33d/2Bd5c3zXIWTg4FOdAvv
qzNmQwtMSeD63upbWTEig3mC5TsUQFRV905Bqchmu8KgQ6it2ULdUy8W1+UlWjyeJqwa6CRfzAhK
yLiJWFt8m/bckQiro4umvixNZzrim1zyleinXxuXY/2qHNITHiYK/YaP/k8hKqdvsvpfU3OsLyxm
SGwuX97UiijsSs7IGwxiKxOz5VGt1AmvrQXVKd1fTou7C08gFAFJNLNT3hYu2ysEhRklLTWAKuoE
YNVX69XBoKKa1CGtIzI/3w3ha4F8X/ljo75d2c0DxtJTYTGB0/DybfimMJv4pxK2NmM/0dxxFRZv
O0MLP/svf/tWkeOYJ1xaVaNulAyXlT/u5ee0rEOFsGGKNmtsms7NM7WrwMmZiW6gWLvxfP5pK3+U
pAL45+SKORNpnE78rfw3eyM+W7zi2g2GvNYRrwvK7vQXXFqi65m7mKRVazXk1Uf7SyJbjlY1VnNU
BbI0tvFm8PCjTNrl5uXTZq19g3G6cW1bX3eXhclWgSsA926oBppUdb8Yp1Fh3/tXrzJReKaoohBj
i/AmvPHAVSuC/z3gaNs4VG1N7KEKQuGWtaGYlgXqv7p7T4SeWC2Mk2npGrIjPhjagWPpqP2LIWtE
rVL/9YPJn969ej/D14VmWxwPcnY0XKkoNbc9idNsOiVf5l1I7OSwlYj4eR/utYRXlJVXpDNaH/Ci
D4abvzYojslTHcfMrSZcmWCR3Wxzn9y/vT5VLYa1uUPKXXeEbzM/eKiIjvBGTVdqcdoHErRc5oVP
CFtQI2z0mO4xmatqK03xICLxrDsA0HZIetFXvZoigte7g4u1KqR9JQAdxTXFUyJ5xCrnS55WIv9j
5M8hp5wLXU/BqxukMnxGqQolo3VsKFhi48vx/oxdYN02sMJDs/dpSbCs8aGj8oGsCbSQz1a/P1tM
7XVnX7774IW9gxV5J/d+wirwbjS2Pb0Blaj8BW8pbu86rLqRZ61T3BOPH2AlwHl4hF3Pb0tzuy93
OoRsYmyBIDM1C1gI+hZ895oaPBaqcGtQ6+r8ZnXt9C6Fq5UFep9/c96GASmY9TefRECiJVsVIgPV
9Sk8gxMpvVn8QQGBvIp1cKri5x1PlhkKtO8tnTUCLY6P0Ps4NE5e5RoDbu334Yp5gXKH0iREinYa
XwXR7gtV+O2ehH8EeQG31TnCCvabc90pIbX5IHzjGaxxOr6g8EyciWMp5yvrA8Z+vB198OK93VWT
wnSXrQf5Q/72PmVZJfzqg1fpzosf8q2rAo+dwzHPPRKcpG7i++tMb0MOZKJbAPMrJ53kkAOjRLIm
S9qxeZtbBC3tPe38CZ+PhNelQgfIiM07yrXxFcnd7OtgfDavcEpzBszkAzI0FioKaVXgr+0uulP3
6Xvmr3BKEEQQOkZPrJJNtnL1y2Lp8zh+Sx1irxXIRLmu0jQQOSW0SOCYt0ZQzfkaUkTLJneKDlMq
zv5Skjvdc03MapscR/1uvE8nrO659P0TZwI3Q4ckt1keUWgtMo3yF2V56xAS6gWLwVlQccpNJ+6P
VJfZBOR7oUQ8QNbDRlb8XvTtjAfUHZpAq6DPNYNaBwFpqnFmZBVZ7VJe8zYyilynSlzmtedt0bKs
vVYJlYnl79DLLAk4LdzjcaqV8Mz2H3iajM4xvP6cu8++Rve3yfBMejBs7Z/bDsRUsAtbyXAAxJY9
3xdZvc3x89mxetMjhCh1zUyNM31jMJCc/Ltj+folS0n1Qdu+LMtBJb8/WtQFnNb7Jt5VM66hBZG7
ptn5ABduTm3z1xORGXpLRUGG7Z8EPzllYgkVJFwmQIhtTURnIqe/grtI9dMDedEhrANGDMHHaKPK
LAI/1FI5civOiH+DmLXqcsTJ5k332D+zLrmOzQyY37+wA7ygLHIA1p6cJ8uf9gfkD1BBQuEcwiu1
JVmFC19KvN66pgZCkCx1yvPgfnBWvxlrs2LLdoAoKyHCMwvTlA6WjBzQedGsQVW4ba198FFSyZjw
3mBaCdM2FlPZ7iocSsAgHtGHGLRc9JlriKCFqP/CWAj6IGjo/syZrUYE8jnGoSms+vrCVnr0FFFR
DKgxAD9SOyy0Eg85zexCKfuoNtAhK+jwkLbpXTUvA54PT9AA3/Hm4Pw6rFRulajWkFCCGwFYbtgy
hV5xiJ6DMBt28j/nf8b34/tbHbSpQFj4bcNLAWate0kLVDA5L20e1KRtRBqG0PHkpF9h4+My73us
htvPAgbTbP1F2Oi5x8f2e1JJx3XVdQ5Rma1oIKLXCvJaa0yivOLDqtEzqETJQopY7ZjholyFLqGz
C0oR2BUK7CM+t8UF2IHqzaQukAYXpa4Fn3ZS3ztILDK9ivCQBTl6icbct0l6Xlg7Co3WorXp3OKW
KjS6FNcU7ooI8XQV/Ky+Qkue9j5PepdCISrjQZAWtefzapfZpDpO/suqym1QBJBqBXuhRzy2dc+Z
WNfg5GO+cKyp+Y5nc7V/fL6mu1YMREJ5OVapodQTNG1VX1N1kt4W7CICa4PPb/K7Bs9pVU5gP9gD
0A1t08UzdZS7gj0KE4ENhvWymSlbyURkPIdSh/Ggo6voiyooejim5TpNGTKH3ByKOF44N5WI7DxK
B2jUjshZcZzStmqapmZ7M4FEaMJKKGtHhQILAlkcPM6xg3qRn/NMnBLp/EebqVLm3V09Y41GCMLr
/hDb3AZWr5SbojaOLRfteldbWYkeAV2tjNi0dJxjhJyA43y5Q8ojHM/3kI5DtGIgkTksvFXcbyu5
UHpJNERSeIq8EBmjAB0YyUyAv8RK/6GOsVT0h4HclleOXoVizGCX/39k0rJBp4qWKB4uVPiKBx/g
nZWTiFQQeV2hjAuYjAODdCZ5DGc5TGGFX9uf21fdvbzEHKwvm5y+hopvrl1P8BsjwFjFxeQ37Apg
bizbnr9e58rf21HiK1YlJwI2cWGlVLeCoRzUvxELUgemRIWJjv0yrZQaSI3i+4ixTCUW7QvahE41
/Fdt2jROXh7qja+MFGUwzSyv9WKh9CqBzBREP1z3yBBQWTQ+yrFvQ5XBgTztTu9j0eOLkDvYLTaW
kBvj7FDA1Hu794h3R81D9VCfB8OD+ZUydW+cLH+x7HizslSQm+jhR0g4tDp869bCQyHINyBnzFSV
Xy7fEx0GgrxMbBkf7/TtiT4nJdJPkGiykMrVkOhSqJF4dIhphPyGt9FAA856z0Oq2+ufDW/5d2HU
WAC13mkvt/+80xpW7OvJnNoy4PzgwdyHhmOcpifo3cl4Pt2BN45VSFD63IWKz/sj0/l7hwi4A4+t
yePU8jTSS5bALJt56GzCyP5y+vUAxyGZTn7hzVDf/DvjjgWwvTpl4YdpnU8HADlDGmE8kPeYv0uV
DVUrjqYYhwZJxKVmoPLOo/elJLB9jJCJY3QEx98t+/Z6U3adwEubqyUFhnGti5drgSMXOzRf00jT
7C2U4bPtJoNapBIuqac6AKXWSZdHpcz5+ckwyecxjo94ioxkk25u41UCBsYD9r0A0StbhfHnD/pi
N0BvIHwZrAvTkuzpjrFZ7zSzY0ArVIhimFbBB0PWLgoHqL+yMbVa99VjFQ0jVWUsnc+efo2h0SbB
rlxYnYAkkDltGhH96r0/NlDScpp7plYLmh1TPI984R3TJfI0yxRtv0oF59wt+cCArmc4EGosUMQ4
2tPJGtEFECOtMU6XZBKo4VOGvy4DTm2jikknUz4L/WPyfd/ixa3thdw7YevugolnhsuE1Ym62ZRy
qjpn4JK2WMiwDMh2+T8qScwJXQny0MApJ4P2a2NIuJO5dUpLFjwkuhd5fBnbHPbJedIQ61NaWtEe
oitPM1vxglmXz9FDtVtwZs6gEu6WzuFor8Y5NoiR/SyBJO0kFnj42Equ0Is8wjewG/lIK/hCrQ9R
60Tp4pXXf0GFzDU3DcorTEzRQfMYPCKM6n554FzjMdHdUBmfzQsUG8MFfHayWbq1HsvwtmDzkiuw
I8hhMWUscgmfdL5BDk9zx3BNzv8rzZb3raZdejVaIW6o4GaeP/coxOkdfmHL+DP3vZ5S1vSBb4hl
ECjEMVZfEE8Mk3xS941xXuhm0BYa7uHtZb7yLrW2sHIBrv4/3OxlCvS0qdrHFJTKvjZPy6HX4FhD
YTuZx+VKSABlp3sM/85GdpqeizT3YIBeCTZz14NhIqWvbepM4aluGqv+bwj07guXw3fcSib9T/Uu
GpxapbDZ7RoSzMncsB7Bc/BcLEaY4xBXf4whRonOUFUxaI3860KPdwFtZ4f/FGLrTsLbY2uRfdtT
yOM5j28XS6myU+LiyobZtIuyKG4C8RuhxyUKQiWlf/Kr6oAmprS5H8fUMATtEdRr6J+6wYwmrtaF
2lKsdbvpJjaKcBpKc7d6ffZpllDUnfJkIWczBODxoAZlTXQ+6q2yoOlWfh3DrUt5xDeINIK6QeOK
J4ysKyKpxbKckcIr4uLdVAnglKhFVf8Po7A8VaNvE95w0ns8KmDzrn8J78UPdZOZhc7FA4lKazVi
ubEl1QBaaXJC1QydvvC4YRs2zbq3QH7BQaOVke96iw3/F8w/L58M5auRys9lAgdovKlaZWPaKr2B
HA1vfWU2cOZtlZ+qNXBi3ptruMwmRyxpu+dkB1rNfLonakT0WzAyUqvwFL20qmZj6azEavxw42MV
fwIV5BO494zywiSNzj/qLTsFeZWD5YGDrVKIn/m1wwyAwbw4YEkdnIW1r9tybx7pT/UfUSbNfvWj
lzWCXcT7RIzAWG5axtADfTIjto7t75yxkKOU+leax8bvw/ads0QV5i3Ty5iRb2skXYLy6mVS/e43
erDHY+ssIqiWEu7XNYTFuKbOoWNUQGjgjjscS3R6MTnZbWte+t56jZEjd23NBZpxm/58iNDHThsh
Yj+DMq5oA3JZ/jIyOiTbZs/xbhusLhPqTYlWQ82aBD7pVoES8e+edHeFgcf0dRVbfdzga4rhjbnS
JQtLSN67sY4lGP/r/wX2ZmTdYIQtHngEd+xahPPt9vEhV0xgkBuJNvpCQ3drHckq4Zvj/mDaQo7n
yfvUaYG82uAmXuW+2JhmTruG+cEsW1Q6CrzXVj0VSwBF6KrFn1Gc/iOQ4zoyZ0wbs4+fNy3UgTMD
MyEqv8qHW8XX9eIlWW9ZufCJ0qUQ/IImSwd3Omf3bukEsLJXthu+ePmw9WHhhat1Tx2hmuCgtpkb
wtL5tYJQPnL/mhKWGpEPeODAVfqLcTuqKgFt6T/2/lTU7Nv1SJrGbLN1XSIE8+YONkL1YJbSuDXh
ChOUU8eKy63ics26BqbT664ozk44bDyP60YKU72HEoOa6/zNmx0aKnttqUT1iozni8gOsM07EYex
nXEaQMCS1TPtC5T+emeYDN8IZCTZdz9/Izv4jrwCKqysAx3B08JrR2Iav1ReaB40zQllgIf775Sx
ArjdzaQv1DbpWBa7AC4YNajhWbY99qPyVYkbWYn5Tbey+5dq4DoX7BmKvTiecck3oAU4ET/pHtV1
Zou4UXDwXZ+a8X3ZlfN/vlwdXy6K1ZEv58sGZT9FW02e5DWyl7ByATpywp3s2ODtXe7HgzN+pzyq
eUhUbB0DBRMy1Ed2RX0fxkcd0JXiS2ckz7Z3Vma4ZK81arkVs3bChRiNFDqI442fNfp1l5ocP6Zf
T6Rj6y0K6LRVe/Ao5IftkfQ3wYIg0LVNpYyBfb8hhEijm+nxojuTmZihqMj3jwQlNUZc6OZ2+qRp
gY2U6eZk2lTrCW7/2R0d1wOucH0sMcq/3v2qeYTlKtJhPeKYmPzMVAGMj5EYLkDIaei9NrH/Zmqt
YquG6PJLyHnO1n4dSjC4a9xDte5yYn7gESyKk49Z0VwvmNw4Jpy6ivBweLNVHENM0yHgnbYVP/IZ
0HDADR+6c/j3M9E8ojiumqiPt+45RghhFBr2jTRVt3AH4Rz8AMmj8rT+WEENhj5qHrj8hhhAmwXa
TNR0DgxBqlFOPPs70H923DzNwZHgHDjJxbS4Y6Egq41P02RsdxJhWKL5U/fowwMLR8cpWeIw+cmU
S3FCx5KPuoSO4eS8W1HarZaOOPOy0qIjuF7H3qL54etXtBIg0FuO+ZzNpv05IFRX8v3jkhW1S9LM
bPV+UbJMz4KkoQBqkLFEwgBQOlC0SyAMaYQbcfRdr68A3pMlU9WA64LcF9ldNgzkj6dvxK7aUc2k
VZ1ruRZoKYv/94dPvAZ4Uwan3IsEQcvM7sWh8RLUzx/63NWez0LikciaRxpo5cBUVPWqHa0d4ljH
/POYT45MzxH82YTpvCWZqFozhMeViIz8oPlFlOQSFZxr1HDQaOq5u2PAc4phXFNDIxw+GMObE/OS
uDEfSjweaXBqEgWYA2qmlBIFJPf/df8yOV9RZJ/b7BW/m89unECm4bLQ//1BksqcWtP5PoA3TgJH
3mONYEkEegW/HRia0MM5DAoiKuQLaBFpAnDX3+ThAzNWeEu/LcfURfY/45iE4GPszkwCT/qCIxX0
4Z0oagiGN0Qe1QljEGBu6x8UluT6yF+fRmEcTm/Idj6cbdday723SlOQacneN2qx9hg5XtEaqJd0
K9nFC4Z7rN6roZVYW38k00VWay1+NjwFjCYzGODCnRwCWWNlNvY9Ljd+gRRAxohnQW7UtujxDu69
I/1o66JJxT5Za2Cokw/ITcQxrNaNBsaUAPIAC09RffXn1PO9QsZiCfbak8wELzAvUkn24pL5ktPW
8NvsgNBiX4pkBTRs+7ZW4QJlTzcYZ77WfEecuCVCz8nPe2IzxVO40tSAsQcJ5/CIjaaStO2w87Zh
og9pSQOVYExLj4yK3XBT18S+/vhD2TEHguKN4Y4IzrbPLeWYO9MPCUjUjI2ddh/f0DOsEiT5PRis
NjPrdrkVBT6dj7/hLBxlVGkmNZ5j6Z1dhmKX1s7fsaqyPTGeoFpvnNQA77HUO1wTYx99kC2ZlVEF
m1ORiDu5loAXlez4nBL7W4zYx3DcWmWnesvrvJLgYq3zmcNTvIAQMzl3yHy8nFn7wyhO29rr3r6x
j4LpnvNKw5SO8rKzGarlqBbUig20wZjOPNl0Z6g2THV3m3TuYxGD0oXfZReAg9E6z8JmbTptS427
GbpG60sd5FqTEvjVrPkDFf+8ja+RCDrT4SAX/7smtKK3FD1D34V1MnND6zN5U6vU/+IcClNCXYQR
a5LAGTnV0py8DF7shm9bRKbX8WAzKo2P/FKNqRG0gz04F0j8NfPHsjmwcPUHltd+VbyFOyVVN+ix
4GgB44/v9HdhNP0TxNY17trlDYfLGxXay4ZfIyvYxNR0femclZZScJYxN+GLXQ9QP3I/RnxHSYo5
UgBrkYSZSAUivUQELk1nZ+wX32VqBh91nMNzKZS4pr3KQUFpgOz4IYOu8XeVobcKhO71dgbTx6SJ
Dxkfd8oS+8lANCnerCv4tkvmRY8Rmr8SYv0+sCQwZLJVrHsxZ85vs1ed3yq8Ho0cSb8hXIlJfTMw
gA4Rcly9yc2VJseN5mkTlsTYVeJYvgXNRvTz1NnlbUE8X5B3kAMFaUIa5F/7zGNePQM/Omg9O4Rd
FFmM9I5nKNdbzkmDBgCnzWG4KBzpPS4DHn9o7jkMsnyJmTNlygJ6rzRS3v9LMep2kNUWYQCxdExd
CBNuLWDBImpWJ887BdwLyoTWK140nqr7MBPY7zsjzzlyyZ2jZclNbBDH8aBtN+6qGvsk29SrYm98
cdsTEIzFVeVBj4tzEORRGWYfpg93g4UaXxImH5lFdN95IuMEXZg/kXguYW2D0OMCIAgeXwa+BYsG
kGwFWzGA5L7jgYx5Lnp7gGpS3IHREutGy6RpsyaT+Tt6pj8jG0vEz/T5sPoAH1gE1rvIU+oNPhGW
jnhPFud+P3NwZiQTv1naeFkER5nQnFQQ1uFsCTlkqGpimwr+Zc7ci2+8SA5YI0Cm9UYh4ipMvFCA
ZggKqrobqS/NTg7JUM5u5vtonoJPR7+hOAPNSwZB2nzC5yo/Jd9VuYfVCfBhcGmjxMVSYHqtSUUv
O/WvQEK7H6cMHlSPhmLgQ+paYc4L8BpiWbFKtbLExSlQD2Tamk/axmrj6vbzHwhUvqTsRY50gZi5
p7nM/PTrrebz57N4HRrSRgr2s6dA/R3rG7RCRKFUrY8CCfPvA3pKDCpYW82+OjSmIOCm9nv2nfn2
ZX277smhL3BFP3qM/7DXB1ETzTA50MoIcvF4F5cpBKkaiXvVOtHxB0gRU5zxCCjSg/lxzZwDSiWD
yla8hlvmh+NuOKgkPHxfBri2eBSjGSBy6pZcbx2JPQX38XhnNQjRSjT/rZcIh20y2MTMFk64oDcI
693FkEaW9mVY2NmnqPFfRGjFwnEYPAxmSllbQxhCrSEt0v4bKLJA1UvFqTjC4VUbQtqL8VEg8+Vv
8WxsVmyd3BqS13Pr7IvtNpjdEddE+CeaK27pwSjc+bubl8UxxIE6PoMjcVfU1BOmTyhUsRIQX4b8
uGZBQj/r2BEtwOEFK8VOWXK6AP3NrikVbYYBHZtyK6uSxNJNYl31VCyCSuWuqPAyBk+1PgPhiyVq
vr8v42P1UvU5fzuSiq4F9JVDKSTqRNnAp2Hcqu6K+xRcn4FtKBVUNYHXs9jjDEjnoce1dJ8ll/rm
A9VMSEU9H/ib8WNXUaAmpaBU6zy3Dx2jp9z8dhi8FzhcLgnQvnnOjQb/271RL7BUAmeeVfkO3lyV
3rvQs5AbarCR6GryeTUqvgRv11STWOPPhTyLrpPG8Dpj/4QgWfCrAH1SYs3tZViC7PgJaYsmuZWx
dVCJHKQ7jFkm+EL0bU4Irh1iBtU05EYF1nZQbuy2bKpD+3Cit8eCkcgNCNOWlGCwGoIURZq3XE4S
irgjW0CoqzR/jlNNVmc17e1steGo5BXWc1yG9os91bS+mUKB6FPWm5ZJGJFmR7n+3y1iPQwglpMI
aV5PqcvUARvkGtGisAddKF6QI9ktxQZcHC4U6mqIzXLDDzCZIBXINr8T4adkVRbfatJw6JxuWmKq
pSxaiTapChvnnAJhyimR80qncIatByLqUsS4SumVrbKsbGY3uMMgiTiXmVp5FAO6OA4TC39g9iqL
RzKS3nbinGLnCFCNFCYpOCVP6FrtjnamSMlJZO8t5A02BdK6C/wQA/6TAkPHzq68EWaTIcIeOoXJ
ij6KfixIUtswyVSassY3qQQUhkmEvBsWuXK8hK4B0LCXo93CgOH+yWVBkwd22XRNUrqM3wA1PDi1
2ckvftVVSOTfdYnTOMb55/Y/ka2mxn0NwlqYg6OiKswWH/PBxrCl1HsazPciVtrXSaMyIn9g1aKK
07iHhrJon39D4K/2Rp3k0tUEVZKxUzPadV3tSl2AVofLQZugAGnp8ZMARgnRs9DpSKNw/dhFLOWB
2ZVv2MSKrJwHB1YEvy+nCNN7ehxdCTSwsdSMDjWw6ozuneOIOAetvfk2IQY9jUAquQkmexo9IdJT
QsL5E9n8HSWwjNojAuo/fdIz0ZHBBsjGLv1a6dngF4fSx0Dye0LRvK377MUfKs1iIU/DYgLYdcIX
BLvKCpPY9McxXj92cNFgIfha1NNeUYK6XVNz4RWi0wUd1TCXjsDY2oIsPHGOFlfUsYAlDpHHOvhd
2EVjT453A24bGl7uHT4UT5CgYrQxltSAC94WTpOWyPJsg4Yzr/bVZVEFBJqVYjxmX2KjET2gWGKC
Je0+s2ZzJUqwK1LCBsXRIf3Wl1yNhjcM/uvfLi6TqKlgqOTkF2+oNJe/6JXj24CrZwnrF72b8MNL
BSW3BuyQxEbD8NW7s4Fcr8iur3dle43ZSMfY/b5Yvlx2mtYGyUqZzFcsIQtAXCILpMtJte2ctw4n
y9+hsWUdZhaSqHnwYNPs0tjar9lwcC/iI2aAknCe1Jw3fuQsboNRLrIwseTSK+gmcEnlb6a0bSFL
+a7FbtghXLoPJ4EIbd+sRkfuNVUkZJ0UwaOFDzTQcj2EyNxXUZaEIgcRG6cJMhY9iMzpsVcgG7oJ
NVQ46dawVZ+JR5QSDjM+VYI4tiWoN6RKrVALgJndVs134sZOYPoYlDcGVYqHwcPijF0hyBCEHaDY
41sIgKglfYyh8p2t8WOhqt7J+dfPVFTQMHL6y/2Cs5ShsAfXh3AisIyv2kf1hWsrlvLAjAzOGuuG
qRe+8nDFn+VALK9MxLd6G1CQ4yEQZ2tm0e+IE6ebmZdWN3yIIQYRXwnVpiy22DSox/F+w96URC56
k19E69F6lJ6kqqBREvu39zuX2x6PQMl4Vb9w3k8u1XUQyKCzh6/BjGcIFvnGcUi8zyCz9wNXJlAP
qHjF7qUDyntrbgjEjuU0lfvaCo+zLZsRcC/8DQwEfpVgpM2gsGO6PcgQr8EIXPT+ciAOhMtFIPpP
a9bL075kp1kVv7GAAo7rM3EbgR+pWuwOfwmYZGkLsN/T0vYeYZyHLYkYMto2hZBMh4upa1TGdH8I
6v6/FaMk6j3zIt+0HladB/+g611OKcSsBNDLGTIQsTT/HnrDevZOxd87K32IodkRb7nVcjnJcpAL
O+fItGgsH7WN3CUyMZ2qzCUtSHlIqAaU6+H5Kp6DRngQLS0V0n1ZPezddla9bK6msbUpegiwD7NX
ve5lQajvmyomCFQSbU0mVKp3OoVd/Vvb+DiRoVRnFlao2tE9WvriLsCGUCQ2zpllp8E9yuO5m9jL
cQ3XuFsO572qhq8p+iVlLXCZ68kANxA5wkNuG8JHHh6r0gifZSpZ57V+wAGV4xHJh1/TO739idFr
xP+SiyVVPv9oDOV31TqsDVYzQiNpHCGikwKCv/y90wQdHLbREyNz4NITyOKYuDj6bQG+359z2GGn
uZmXtdSqc258Ds4Tiw4fn/cDtNygtMMrcxg/8noL/EoLoYnw2bcbP8ZG72oksZgCGXc8EsJTOqlo
19FWygTITwgsE63G0kbPrFQ4BdJjQrRJRr+wy9uBBOr6xXopW2aOv0MvyTjmf1+MSFQ6REpJC3h/
j53VIDdebttN1vsHWpnDY+QIERU15FxJfVtS+0tQMjsdonQjeQJcbP516ZMgnpD3mTGCkEqKWB26
/NwyadLxAt/nhg52YDbKEZCT3TwpDqTCSe01yAG9HGGKcJAkbc5o0HoKY5ROToqQunM3Ev/gKeXf
g8zFQF+AYvcMiF/cnXcxnDzIPp3+7hJvp4O7/VB3LM+UbOQCuVhhMBM8SRYV6sw0vxEW/9EL6cm7
peUj5LK3vadaVStG1mdQp506Csan7CyXrfb91kY2gviVj4NNLe3aa7t+b6HaTP0+MhMSw8iL37D6
Fu6K+NFREGtlrY9wQjtvLO44eFUAV+skVGFP0snWj65Ne//B+567Oe2JW/GaYN8hrl7GZBGdhhhp
9NoBP4Z0Gp/IOJ1weNcZmh9uzypHIeTSRdKJ4bkn5IAvXmh4JCHsZcijsKgTx9Q6sjooBND1ZIYB
BM2qzHxfJZEmzHrKHik0PwPoxTGbL/rda0e6n7PPIWovXGaL38pPbfJ+nbwyfhrr+CRmgoTeSm1M
2r55FKfFcddghvXbZB8l2RNNlnCZ5Q1Ue/FQoegkSSBj6sTbC+g0qa5Py29w4DD71DkavGVooLxo
FlAiw7X19teczdn2t5z+PYUT7/z0n7p0+GIiodfmqVrFar2aHX61tUG6yfV/NHrKTThWhviso2eF
Tt6gK+w5EDx1m056NJKr2G+QsOEVN5eV+fQKpNfCi5Da96GGDq6eCtadaG+INv7mdJCCT7E4irBV
OI1eTBQxNJ+Fwd+QxWldD/cZILUXDI1juxZHhcn3h9WwWC5IuGirfUghZ1K6aGy0i9tALeZ8XE5x
VmqyjZVgZmtBTIsWOxYGJay6p6VAi2SfvD4mRnpruKsDiaGlxuLvgY8MMeD3Nha9+hdqBg33a9fG
wTomOQZg9oaxWaOE8QiXinUulXOAd3BkgS+km9OLC6TFF8/oRYMARebFpdxGbfCQGtCrh6iqeCW+
plqdrGd2uIa6gdp7OU9IZB8gz0p6BWueWEcrTLFHtdG+IZDvGAY3uB8sZ2ZiZqU3n9HNDKOvaYdS
LkB+TBlqoqKEA5N98A105nAQ+hEAJLEE5kUMUlbJSm0dem5Zi52E/ZP6eMz1ew86BLWsXbHZ5tr2
Rep5Fb74medasjWJ7/WM68gUrWLmOP4M1o6t5WdA0nnx8LQGUNMdwWHpt731u6uuhtIUhUAEUSDg
GnEn8THeqqYTbcV3v6RegXaWhdn9jll3Rc+xlRngj+VonOkKRCppm/+n2aK/uB0DHI3YtuqwsmYL
Dx4ZzCcDdfAxGmrqGURcKnmUDe4IrZ3emcKLWJwzleTSKJpNnc61ZjXeDM1e+w2Y5+tVqjqVy1fY
TKHKTWjXULFZvpudlbkZNri76ersxQ08x0FKHrZA8XQBOyrtIhY9tnQ8XolwzTGtXSZ/a8cS6wMU
+9sfXaksndBAp8ZbT1oH6SqBbiXtZaNmyPgQP1WkrdlnJdkauCql4NefwAE5V/SuOXqLxvhlqDyy
N/basiIhLk7T+4GmPvPjwlGU4dvpI7yIEi4XaQkkFO6ldgVUMc8FH/n7l3WmRXq/LfZIQPUUhScQ
31RgKNRhuXm35u25C+kinJrtt08OZCjBe8UlO+/9cOg4gTTKx1SmpAyEMjT8Lqv+9taoCy33YeIF
IXjwHErXgE31YNIOy4dXvx4RqwsS0w0Rt1+S7MfG0yVLvflTbdNEXY7ZMLuaeR9qYUNJJKCHZ31G
En1WwZPa0Z8nj/WvoFXzQYdWSJ52Jc7MFbjpZHswOMguX9EH3VxjnFc60omJDCk1gWQl/m9gGJrq
nAWTwgfQyCb9Ga1f87KLEICUB9PVyQPniRaykWSck/gbqdbJzUUH7rWQTspPqhjco4N3SMB7RAFq
aZMt2IQcSZFZJ3KmyzQpTBJ0GJzXAGI/SBbnh2C3nLfL5t29yJwIndbIv6HQpFL8koQA7e/ZyW1q
XCMarTvz4JISzxcxFHxp0GRZ4LPH/ymEmIwvKa5d47CxkYGX4pPeyb9JM7scc591N0FGKHLFmUtW
ml2bxysyA6bR+F7LGMseOi8lWMuwH8yqflBI8N4y7KdRPy1/YewZFHDwEShSmWNuNFD4cF+k7XVF
XCQ/oD9J+FFgsrSjWJTN0czA3knhBNwfyNRpuMfiDH6ZaXwv86yG+62YTtqJdZRr4143CQWI7fAx
cQTPw91S2K5BxnmFHaN9J78sh6eVOGgk0xLP7KTjPDsyuSMvXzBOa8SY6aa3pbnvPHpkHqm84qgc
/eMrwEzNxlqjNZYdirdJVC3iScsjngSbT+6uIMDBsqv99mwd8P1LQRfF5iWM3LAFBueMdzEgZkeJ
sNAfAuxgh/iz/LUGfaZ4t0CdE1WtNMRQ/9CLN2J4s43Uied4BczE6V+eTOrEdaRsRi98IReJ/stg
tpiqdF3ITSIT1Rv8SVi1fXKS6P2Q2Flo4z5XGAyx0W2oD5SSMwAlSdP7Efcema0mcbW0jV8xOQwC
HR4Iv+KzGg4fJrFD0LgS80B3yBdiOiBmKVD97qPKKO4Tdl1HPaPac3moq/LhEzs9nj/GoXxqIWxu
q/E7TnJAVSDbblEo+bKJbPn0owbURQoj/6wI7drzKeFneKcbY8xYu4xHe7qqhxA41cPHDTcmgwlM
gn9UxhewllLrhDIq0OffCbuiPsMAIbjeSLjfXVuJRXBmROTz/fuqzjefRNIz4tIRL9aLI0qKlwjc
cH031U8PfS2bFfvth3DF9SGvaHcW0Vn6Ql8MBco4xIyh7OhMqCfhG1YA0IGvWydu3bhmJ+7EA9nn
Bo0Kc8QeAYuYv9noRaYJH8mKpFQAYKdn7tpLOd0puIdxz4vGlRYwcCk6kN7132/MeU8e9ozZCReW
39UsPtOaVu+78syKHRy2R1uHLK5hRj3dPFL5pFNkMKFmytyYGVMO92I0+E0X2FhbVdRQo/NKYGB6
mwGdZZo2/Xth6kYoqG7VQFvCYaHDfmFMkS2xyn8QqvPHicULeWua4awqwQAax3h89xGHKgen8YoU
3qwf9IiPHxo1I1J+spMZCxtQIctk0QogCYiBEFgkG3PAPbjoykzmjUcCLvFtpcNYeC63hr+h7Q2e
uOXXOw85VMczBmub5uud/qTuk6/b4uGBV656bs7gGHDnaPZibLRdU4aIJsJB57fOtFmDc0H7pCoH
ZXvAvrCG/5mOMHNxYiKHDAAUV/mlgfUg0KpV56bZBvzARFA7tUaUGMQHlNEvn4OGZbWHNCbTEZEz
vZtu2imvWqM4KXlHs96YZL3g05A4/AXjJQTwMpRSjF6l1aCXF/NSGKxm/nC8s8jMLhKmUYjVCng1
tH3BIpgQ6y0A9A2j76OPzvwrZhcxDxj9a7acTHKCg1mO1RUZMHoJ/kNgeCeHJ/EZ3/gGLUCH2onE
5J5CyOlL2lciBNHMjWRHu2DOHnFwiiye6reZKpQFDSONxcFT1JwsE/L/Nc8Rs8mbA5kENFn858mY
+ZsEEKg7XuV7YALfF6aYgXJmQqt2EmnNLSZVkmHwq/Rvo/6UasQYmKGF+ajaKI9Gxm8gnl4YT4EP
Y+j44XxY5wd59rhagNW1F7zSM1t0UDJhTG/xxi53bUaQQi4msRQFZvbNQOUEg2T0wXgfUwwqfiM4
yQa9oc5oTJNE+44GnPxE9/iY2KmrDXHVbWx3t60dBr3RQadUPLrwnZeya7H6CPN0eT1CZPQUsfZc
gKJATFHyhxP/hBMvTdJ9CCnOON2StIwK7mW5mscbxbwPC9nypwRjFOCcmK6L5P9sRxOnVkJVUkDH
gSzbxNRNgh2Go/e5Yj/6g1B6T+4tE4Zr77D6/nzxaZSjHGfpJe7OuuYrnzFvrosFX2Ne2JrN0btv
G/Ame8CtH3TkTkGv3Nmx++RES/cSi1Puzt0jhCGWvvVdh/BToAjq64eobasmpfrOQcMg6qe0Joc0
pqiZRDypOA6Hy2vMZb8cBEMhct93KJvw5coxIgqzca2K05GQ4vrabG9IUhluBF+wiVEyruF8NPjc
ivjKzAGO54aD+2SHbbf0yQx6PngcdQv8+B5JSkatTPZFE2g2TKjSka5MGW7eC6kjmwA+TM3ru8DY
Q1pRct8S0cmGofaK6ZookdM29G9OX5nTHAHRrah0TO7m0DeLd6xeutYyVKVEfcFzPjWs2row2QYk
jW6XxiiLp/HSx6I2OpfNPPTqwX/ehwmv81Vqqu9klAnj3GjpDhg4q+O/C7rw1qh9r7dg8+VwLKU0
bSdGv7gy8IU2HCmnTitWS4CJru9RdwcchOSB3dKb10wEBt7SneWNhfQymyCfV17Lrs0/Vtk1k6w2
WRuYpxKuwWsJbzqTq02ouu7FMojR9yPkCGhkIUf4779Vz/bAqmQo6HdRXawytk8z/rOtU5DrgOD+
LdPtHSqQl6AIRW0A4jTv10g9u9mN72Tjd9E+Tzc/n8uxnLNuDnJhXfLqiPd8MIPXHyNJXF4P8bvc
8qFaESRt0gL8MNDObxSExWXk+JWurhrFXu9yTCNSBNpo0qS7o1d9c1ppz9CSUgU/+VuZaGoqIi7a
jADl9hCZ3SVvPmD5I8EZBBddLrEYtCvHGFJAeTThLJNZ+SOuhAWLiBruEapoclE100L069D0kllN
mJZ7czdyKveCz8J7aQJiNcYqmu5KGYFbuZhkFaqXu8nOyzKg2rAIl7Ct2ctnu+GP1z84Ax95GCPE
+Y6cpQlRo7y8u79HByZfYtC578RUMq/S/cj15CXJrDeir+Ho1/M/khVVlk0Bw6nKViLqfBi8waXf
J1R8qBUxKOdjYyu7Nndg8BGCX0fmBZN0pvkwp1H4HGMdES+X+Yt1GaIGtQDKbguVEhcKH8bW0xBK
2T0uAOh2zJSZvazBQPlXlpzOJw5c2zR2UQejboM6NipjA9/Wa7R81dbKB+apKm4p4NxxFNiLDCBZ
iiMghLQBcs4dblykf3Ss8u2X6g9QqhVEigSW9Jy7w+fd2xU1rbFt0gtF5v+gYpORo5CUj7XDta/w
5r51UHTbd+MyYf8U3wNUmg2HLB/rdlLORrurRCh7rpB+PWrSW5PMZFSH3CZCBqp0/mbDt3c6kaEK
APOXy9cIQj8RHd2Mhg7Ph1RmPlRG89kZ9meHFTKWtG0a1vCky8p+m/mAdFCYOnfWGTYeRfkQ5vEE
Ox14sEVOzRiLuN5PJPUmIjgV7THwDLtKmirUfGr/iLnJ+SpTDpTFNaO6SMmtasDZH72LjTKe6mku
lW4xjcR8K3RrXS7xm4gNx/ILkV0y93w9I96ezGoLPEi6AWrfX5x2nf4rKZ2oKadAsB1gRH03Jyo5
MQpdIS0wge4S1MlihH3htczzX5G1X4TwiOvvLPK7cl3rms6RCZmIba4zWHBd9zmQEirVVLhyViTy
tfJ3QoiDBPz1drRlSPd8taLVj+sUMq1AcpzgJI5TfzZTSEifx4Hms34RxDG1Mz5j1UFmaenfkN95
dygfzpttR5e6NxuBs+nVMwUANnAM8S8uDMZco/T/XBsmZfoJDlxWPwwDHZN/ehAs1Gv2ZFWKgUpC
l93W2qXWH77TnGUJh/ykfeJqUWsJfppGPWN1gzmsgQEuspSS74fckddTgN34fOohiFA3kt3YGkEW
T4bbAVlR5on7BNXcHhXsSh9M3VA7F2S/dvuUosKbkNIAJKcvktWYUaiG02+cMvDAAOjhObtJqyYj
uT9x7l//JZmXkm69aINGD9jifYnagzR65vGUMSLRAEdBMAKQkzg78a/fe2fJaBsap5WxGgbCFl/a
HGHZdVjsgfHUptgwVmL/W1kVP0URrJmSb+ZFS8dJfPfmm6qLwr1P3lnv/SDgZhYxxg/Ljf55wzbf
lT7buQqe4Y4CQ71myUGQlFd4cAfkz24joUQDG6e65GGDOs85LdpzhM36MUQ4G4thd5Tq75oXJCt/
cLP1UhItZeTgbIY25Lb6wWWPKknDK1Gq5PC1cTgGKe2yX6FQFS34Vgc3vZQX1pyu/Zi4kHSPsOxb
eoUjoROqoKU+yMIVZPhuGXugb8SS9/AO/HBV57HvBd6R+VlZKtAuCg/yxrdMddQLDC013GPa5IQG
l0DBtPtCqfk9wKq95M7HHhCBR8VHPVGClMEtVTpmIdN/Icg0G+YfWfo4L8wOskV3ZhoWBzVcXS/w
XPU4RmS9svROKd+JZ3yNOdN3GWe1TcLDA57e3dj+Q7E4OPk//4cTOWQb3Lm4bzIipOBNz/spU7Lj
JMDB6X3SFYZFKaaOzMm7XL3IFVfZ+/gvx7KkpXloYGMn1bNGPVHhyQ24iId9sQZrtNDjpMnL3Fmk
p13lblFYDVHyuid/3lZuQBcWfDlj7QcT1BXWpkpyTEFDVreI2gQOWE3Aao9irs2z8O6z2kXu2vfe
vOqDM13k3TktDgE1wXmngdfW7/iYYoSRBoUbNKI1ZH+6YYGhZwRZu8XKYq3WUP2u2IUZKJOgrC4G
nHJISpibqr+xF/nIdtoyrs1iYagHmIv+aDQLw6jinQDrvZEwH1yGQat3fJLIIdsfKnsivUY7mK9k
MPYbl6l60dpx3z8JA6Yfr4On8KhHYvkWt2ITIBYiQ/KJiwGcZW1CMdMwgHXi4115zhF/Lvgv4yNr
kNai9wT+FTDXxrm5aJW13AxrXskGYL6xrjKP1cBk7h0ObC5t/liUsMuKxFPANrfrwJ/jDydXmQ3C
MUyZNucIuQvJf272PF3yJ2M3JfAkoyl86DrO6guwHEuJTZcyl0ZCsDKnBNKRvYrnHlIn8h24B4xl
d/EtjIjEKTfo14lFJCLCXKomg/Zvixw+62fQUuz6OtZBpzF9eW7TOL7WhGOyZPEU/GMQ04F0ce2d
+RZs6hUaBosHtmbDnu5RBrREHeeVUskqqpWS0Afxdp3Do+J+tMdZizkPzPw/5jR9KKCp0aANJcVr
mnCQNjJ4NAntSUsE4eUR5Hq6Uu8A4vw1QTKjnl+sPMD9Rmla+NTFVYCgrch++r//Z+KqG/RMDAWE
bEJyQx6fca6El53QKxU4+ZQBjoCX2sOBgElN4U2yXCKqsSsHSWpRIbNDmXFjKACWPNcecz7hiGj/
Rw1M6fckN840wCXj46e1PV1NXwU/3wdUJ12IHnIRf4ZXZpJvcEhQTC00nl9sqMbRLAqqRLCd0Xpc
m7+cWEDB/CouDRhbkX4Cw2Gzi5YKQ16KENfGVnQZUBreyBQl1u9XNN/fI7B4nFJYp6NjV0TAECaR
Gg0pUcrecYpwzDSQtu6lbtF3+Ig/0jtUHiLrUMd8PqJu1vPkCqg1s2xDvRI6G6HYLqHFH3yWsH8J
0AFMArOiQ4sdL3VMMKkwWkERjTtGOQXOIf1TVehcvfLVhXl5AQeHwEWDSuyF0SK+R0+VCTvrQ9s/
fTjtq6AzTx8O7xyWvtHgmFze+3cUAXeR1LZpXLjpYE1F3BpKvmR9o6OiMXwp2gNpLSIOU7jQ52Zb
QbF8DEt/GakjzhaWceZ6KPYGJCfOkD3/3Kdrk7BZ2gvLTAIsvRdj0qrrDbxOi1OGeBGmjk1n++8y
9sYqCRTajJcHSHqpXfjToBuEC1FmpwR9SD3NjsXIGHceVdFA7VOVMAgFw+OkGqq0fM1wlGItY8Lp
fU99kvpINB678fssGi5kqydkEPRxI7jpEJHB/koqn46sXMiYR+GDfzm0hBq6Noqo4/Zs100J3gpt
cciPwBHQ8MzhF+W/0qu54a1hhJGU3vfHrjuA75M3h7bxZIenYwmP8j1UyrwlMhcKODO2kCcJMKHp
2W9urp2KO+LJmO9GpHcNuRUqK3ZJCOHAkka8vsiJlPmnOGYV4YAHhEDmB8KUzoE7YAEzLj1RN1rf
sVhDbJgmIo1ZQiG1Lk52d02am0d+r6XsOBrhav18rrh+iI/gLufepF5MovaEparj7mzqNDnfONu+
hErWt3YbypMeOa3l5/zeIqzCKGdPlfwUxlltI+uZ/sQzrVLy0WpLTL1kqXFk26z7QDW5h0kl5bV5
0iuFvazd0wmAXW0qPp1j4VkTp0XKPAQBpViYFk3ABFWK2T05rlAFK0hi+vTgzMzO2SDJGy7mC3A9
lwKzWJFEzv9fzRtGIQxaG02RNVfyCWB96/1ZUqPX+gw2k93zdcml/JVglIwpnIwuXPNkPc1UPMy3
hAyi3EUGAqohStMK9Bh33dcFG1nmaRLKXLzA0j9VIoQgx5hWOl54Mt1MePnIWaLAEsWwSq1a7pAv
nMtfCAFTLA0sCSiH3/Yb5PGLOBChH5sLbjCAiPsK7bKTQTcBuOySqXNMTNnSrN4AZrJCyKoDX/0f
xd7JgqmUo97sDc/GiLP23GYh06zkS3CFYIFSp1+KuUz0c7c4/1EhAVnj5YfKmT1O5ibIvGZx28vX
kypRT9uB1iGvmcW1A1bfgrEJo9o1KWdIzBDX7Lc/WIwneznk4j7nTsXUL9LKCfjeOHlAvP+AgUbC
4n1pQ+G/VOM1d4WbE9q94B1P/qw+wQBW5DFK2NyOu+syDYTHHUts2AaQcYEHjdvuXFPUOdK9RkQO
uJWOf0f6MbmAbrkpBVWR7UwkSpbh1wP4GVFWAP1cehPeXzCPpOE9MsqTzacXCU+FhJ1a+XNiWoVB
BDuvE8XSA6SgN2yQycOuqlLaBTIzffLsVmlHHeDinoAx/jfpsUKFFxYge8DwS+LOF3JK4EKrJEb8
KWxu7JjjdE1JjMtU9j8s0idUIJxvAkIBKFkBZn/t7CA93+zbuOebNM3RjuYNpGJ9g1DjevslSmgD
CIr8lMNbmGV4mSnWCb9sMRjO+N5IFWetn0ahVFQZPLqdeC9oH00dwuqBKZFnT8GDsCzMp3PVdUGH
JowKOGDYi2XlPI5P2MuSumi/6O0vWC2v/yD6h6/B6xqS3wowuQroRZSANCRm6ABQDGdlr/ofztxe
bZyHyuOYApPosDDDQ5074ZbreG1sPjJgI7l4FW7EihxGzlCKWlEsAxRTyhkSeElqbHDm0JsyQmkE
cOQlMwn2UqnlWsXK9JoNPQy9M4LYdyGa8JaB8j81XcD9UNAwjh8N8AnKM3+PNCyHLgEy9HxnqNrC
mkYJOrUPquekGEjWGVv0kVd8Ab7/EcPEV2nRfJ2O4XtEfZE2wE39gIkCIHo2AIdBr3/mJrHsIvgK
8ZwVnRIWaPSUgQnZuTgfkJ4PybcSGNJObPpi1X2ox74ptM15gDVuMcNdw6xSjkjav/p0xxArHp7R
fIh2/CY2QP0Pqu9XsUkQN1tXnggXG5k7xmygUQoQl2VtAegifRMo7KJu09ukdSVyP7ThuR/Go/nj
ekJpZD62KY3he+JzukA6KliUDHvaEjF9YkAtVRwi23ZzMGpzszq/Hm4u9zi4EPFRX7Qwg5m7ArCX
eViOIs6ALKLNSssYof1H1TWNBhQQOse42aF2xrkcjNVidQLcWP0T2TvH16bG8NslAc1oPmN1L/k+
EHMHNWqn8t5mliymX5zX0w8Qlws9VSIBjLGNIr6L0LvyvlBRXx8JPB8Jn7GJ8IcH3iz/76BUXlrj
H14syv6etPc9o07Bpl28fQGRf8MgntioJxtOVx7bCoQ1FOni+TXvSG4ygjHHwNEzuKiGrl+AWh8C
XH4cLwz9iMGBKSPHfbGNn2KvBaBPkdgtresKHfFuFnI0YbgEA1WRg+4Ub03ZvT1/oKJKmlV+HyPp
YWxQSdXDWqgnslsGpg3Lc/GpH7AS3RIeQMQLWR05+OlmHYdkqgYLzwuWZUGtBMq2L6U/vqaqw2yy
RNezduroywPyIxBD6/hjDX7K8BZ3lpNFl4uzTcyEp9tV5SyQXiVOUD0b+gwYOnQVCBrPAMG5qm0O
EVSvXv8UrooElatAyskl5jzv6KAnhmo/UPfgcrSd99B//2JZQnqiIlygu/zbHiD9JmVe10d4NLMn
qPSNB2IsR2ii64Q+6d+XJlbkA78fXJQwB38gD3PmHytvRo8f9kdjCLYMRmy4O//hUDr+8xH0H2W1
6FYF4Ap1vZO/bGGoszITREDxETvLNSOtTd62+1NPpRQ/SnZztb2xs96sZ3dMAS3vEUoi+86ecXXt
7D7mN+xQPbH0UCaAK05CJhsOfGc/026+PVqRzb+nbLnAdyJAhE/jhKAXxP+niRkoOkL3ddu9oxGs
GvCUzNz2CFKSJaKSMnav4AeULQ8WyNIftvax0n8NicGokVfYURrZ0wrSOuIu8DnWyrdcAPicex9l
QL5nAqOSm4wwIV9GSA1/JwNuUnPeszylbWNKPhWWiR5v6vDw+SaHnoVawi4dC3yKmWoRCV7ZRZhe
moHQTJtNN2PHZJ+V/eEy4H56UdWX+Ew+03IJ6Mo2eNpYl+1ftF6Uwc01EjB3JHdV8rG08J8zcl1h
Kf4jQ3e59fuk2Mh8bLG2IY8ohH3eTlWjtettlTiCzbEkwu1xG2bnqZgSomjyimVW9OdIriDBw/ry
NyVcFcD99BD+dH7CDKZ5r6XF6IOlhilP73vhiyuhU+ZUeEMgImecfzDv7cLY6MjEmxE3IPrRL6yA
eOmoK1Iu6TGhGDDPeQbdOiZmPClz2O3JJEWmIOXzf+stsZ25n4CCPr/ZFtmptJfp9v33aL0oiXXg
COn4+0U3oLp4qNltSoDSw417/rwukD+vA4cgYbcGOBJEwoPvTo70aC5ymcaYL6awnRuwh44nUeqi
a8a1F+FEatjI6MGoEEjW7lPIZ3Npsomx/ZWeqXdCIznk/LWj9kcDJl1QzqEqPvNWupRonc2q7Dhd
3pAwhMTbA37OE8LwV+zoJ8CLosdJiaG089pjC3cRs5SaViZ8Suirlr+Gq+IUoXwl1ZejtFtJMsjs
CEID9V1HNJHXadZTgPrCjlmo/1mtDrbdqVDB+i6ZV/sOsw3crQO1mFOsHYlnNWuzvOtHCO0kMtDN
FcR7luGLZhcDWpJCBCRB7kwuyEPwv9VP7n74ya5i+j5cKG1aE9Sz8gJ+habqGDjDMgbKJRk1TASY
4sFx7OnivBHIfvFbp5m454Ckpbdw2CVHoUwQ9a5vpkFsHtcP8GJJ38jwRIEORP8bKyvG7GQhlX40
guIC5qOLIUzgv4tC5UcesO8jAMo37Z5vW+BB+bqWB8jgy6I1gNBue/bwfpHb65N9nXT7YCGdLKX7
TZColWV8dxBaWRTT+sEn5+GYbNuO6KncA3Ivcmt/PyPozAl4q5N2/yA0HJ+AXhmV9k0WBnSuxAUI
APAV4W3oEEM56xaFsj23Ug7R7Ap2n7NW+/1YLnB82yVqCTc0PmyNPMd/uef4kAZjHcxONTaJP+d6
BTWgqf6GtCGXTlIQir5IbqAuDuQNl91AK7UXAUL5aAzkGyiczPApeJjKLj+EQiBsfqP5X9VwiqUg
peOWdlKRHNWnSS/Z/aVgee5xmo9Pwp8zEjWCoEr/OoTthNQFphR7va3rzKva5AFhfcd7ue1GK5d0
5fy+S/KKQMflpcQEpDpX4MhfPYkXFWxO+xRGV6QgVbBkd1HLlmxSDq5H/TL7UPA0twOSvK5e3p9W
HiSxPN60QVeoDd2ewNMWpMTldZEeu98mLMepkaSLQn1gcECnJE9uHP7x/04JCuIYXN0BT44F0Gyy
bd6BmqHbY7YbOH1MmbRQQZAaThbTeLcX5S5Ks+C1Gsa68tkdzXCBsVIlf+DzbjMtiHS72mZLSSM6
3sE6cksC5k8pRz+8bROc/w3scYArPyxY6bCwcEoq/DPu+qV1iHLRQx2zW6sWib6JhKwbXRbrhL/D
7vMu/PM+FImnE237NuN1V8cFIej5rmaTHly9l0qYmTO8pP2k0UmIGIvHe+tK7+aYJZLbTm3CO6Ek
oX9t1Y3Y1hMhn7qI6lK/5kK2kW2VqXtmd8BBU7iS5BnzE7jyPeTcyx4B0fhXBGVTlUpwWTP34XWb
ZTFiRmCKonfhvl3PaBaG9IL7eZiu5g7yXKWSGjoW/3kKuanuhL4M4DgwdTvB7o5A/eY9Om5trEHh
xyco2SElSLaew/sk0ha47PEvtyzPN/yZzKAHQOwu+iLVu4OnwYNogi3lhyROsetLObGFkfcwTBSj
LD8uOqktl6TRLqu1t+6PEnv3oblbHqf28t4dRzgs436HDntbN6HqEe/MNI1jDgOAXl58mU2Tg7Y/
ZkJd6q8a6dNitdG83swtXNkmm2oYqjiFUjWw8dKhSlKBzZFiJiIK1DC2i0PCfuVft/YJqN3oynW1
cyw+AxXo9jOgOnJLLV7AgjjH+p0n5w2Uwd9YJJv4XyZ6wSmEpFw7qGi1rVkOn7D3/x+C49990FKi
HL+qmc8UXUWeNySGZVD8Q5rsXXbUL8iwCPTbD2qQpxn1WkeNH7yDVwxfH5tJDIJLIk0d/RTefDN/
2KuqV9oXIi7VgniWZ5BalLV8j+qqe8s3IynL7CnBLribdH8zMRmvf2g38/sMHt9vXq7kB37YyyUX
pxy2lzFm8MmUqjqUFynCLT6sTBJrwjdsUi2AP3JkIOoKkPZ9fMIDuFRQ6anuCmKDSA163puz2vwb
waAx/Ql7S3zwMJ1ZCpewbNhBXGmZByInn7u4R4pRjukSh7D2E3ruAFp4et2wL5OMpvb+2RYB6FZL
HKsaJW+wawz/vhFoFH8RZ4NfzWXAl321Fli4SydvMG38nPtd0Ink+04b5RosoQG8HnhGQDXzYwfT
K2pjTLqNsCjz4SChcySSa/NqnnblPPELgLhCd442VF1vN2kGKVuSO1iREbjdcnz5MQBhDDH4MVOb
lvsnisCQNbuaTWFz38IRSmrnhtQ9JywmDVVTuTJRtDurUYN9VGXD8ot4LLN7q9BGRNd4YpeOEv5j
EkeQ+UQWcHDGx0oYaUyOInxIqrBUXzJm28CZxCWVvr9OJgrIG/+A4BJpiMIHxsFKblBB9GqVqmnJ
6QVojU/7jJnNLtWoH/rQFDplGuSgIgy5koog47wf8WEbi8cfQUVJYlYeeL5vtW3D9Bes7Ake8c4l
XrU3dp9y3ufn7NJC//tMXFYt+3jZnGDlcYF87a0IFKsKe8LT8reynQUI8YGWYZR8BHThSo0LgVB0
/os2qGTy0eTOqCWgoMhaOayiyjeRONdELDgb12W+NF78ShLOyNBVUFy42+LTfVnG3vnl4oPU5Fbu
9we1nl7zuYXhNRGqWKC3X528HW25OMK3nt7yjmIN91Br4PXGVKqQeNf+PS/Z2C+1FMe1eOBvNTzo
vzgwlo5192qhpeJ6NDNkycRrTF8/9bvUKYEwDOKXOxNtnUZY143IGVONVM8kpghxaVBTPzxFoViT
XZLQREjTysTeFRdAEnQDY0NYYS1JviSn4TvI2LoZ9Kdu8fzoMJs6m2ub4iLj4ptYqXoNUA33lPdn
bAONTJLk+n0USsaTDskefE/wEL4oJt2xBI0MoMvYuYBAlooHTwBhcOZ0tL4K9GY4kgTMCPpb0Oru
t7zPl+vERcouzVGdFgHRzp+jsDtWXnrdtvWuZl3X+uKGsBr2Oij6zgXxAvecsHNPyLgtTlFZusxp
TqZ86G3VbP+oyh0xnXTVQif8N1MtOOHtjINjURg1vKCWUR0ht9y8DDQvGmGw7Td3VC30jfjrTL+Q
Uw78/Vp6xnKO7yNCtJ7E00cQ2RLJ6ObHn57V5e5s8ApTufJhgMXOnE0++mTbGUAlJx4zo4idp1nA
oeKV/6ThYM2+WbgyQ7HHeygpWRvYYHy2ylsDR9XvPmI0S7JaqMl9lTJrU0EXNo18jFBO9Xv7Rzrw
ZK0gtsk03omvPptrlOOAjjlvIJ57x1cC6d6w1kYIwhOYO4/c3wsejNBWKAtgkmXwjXzI8d98fG/V
VzTaG4rgApfvSS3dvB4aXHR29GMNjjtxe8QBC5TyBB9xDxPnl1nqILzcYGKHrKmS6bFPCSeTUALX
rnUgTZU4V7xUOQwgr4ceEGMaWe80odZEErGTBPYSM3t1h33PAa6RxFVAIwFgsScvF3V2YIsVsDz2
51Or+ms2UkzObzG20r3+4zDa0WF3G+hRMPnABGj3kD6LQmrDjG1q4v6Z/pZLyrTfgrDguhqSG2r2
u9ayQ4kyruJjaaDllsBlh696Hoq10SN1AqeGLParDmo0p7Nuk6Tvap6zEjZErc/L2T7rNJX0uTbc
NNiX6A9TpMkR73gm/18bsvR3FC+7BqSL/nXiQxKy82dazFxlLmYognxaV+C36kqRnBmMg3oE7rOZ
R2Rzu7Y22Xe3LHtY0+C35rXMXJmTnWdybOQgKHUqgHhazZDWxDIkkN52kYquYbbd39PIorTMcP77
rUTFV8cINIOmT6F7lgsZWxZ7sjUxqpDQdIyI0RBOnoX2ErP7jaZ5zsqjO/1gykNx68eVh9X+5CRH
xNzdLHE3KVhESa20+oA5J9H+TDubgTNiitIM8QeMh5Pm/jxDTP0m3h6ezFwz+fnGe3+5ligVxQwf
Vvm10KFCvOrS+01DL7qBRdKTXxceYE3LGkr3z7b1eN8yW+g24Hlss8zTe1Bi+5Krw14jWLkhVfzX
Q7XPPNfqqRMpNZ5PnoP3PDhQ96q4OA1rLsvhfRdCME7fYZQ1iT4UHFcuJfMIOQYz56E6FHKcg15l
Gja1Xhc/BW0P+7bG+CqSbhCoPyVVS+s/foI4j01/cfUwk3yc3LTtWPcW+E/yWVZ3USiiEBqj+EJr
ey2+nZmYT9Tywww5D5c4qefcdidFJYHi+xkxFDwVKVczX8dUqtnLiA/quOl3HN9GUlYVag0PdzvY
yTM2A0q7Pru0RZ5//myYpFTsTw0LpAzO6gW4whfq2tALWtAZewTch8uoqgll0W0gkvUga6itpBjf
Ej4afc6oGz3Q4G/hQ1sRHuniHiLwtvkjy3p0M/DtiwT4cWUn86i5iTe8U0FgqazXdzwqz3fDPfFp
uj/EMNGODYZA7sesluZS9ykyJ08M1TzytZ1aB0FuheU2kJOKiWTn5eWj99orfbfifj/58NcQfNs0
PWlOS70CxQAhfW4nGqh/BTg/Meb7O7j1sFmTpMHs2oNndLYFvFfywHs8FbWUbwZ3lGlep6kyBVtb
DOyRv3+y6xEeJ29fiCB1RplMccg2yPZm69OUTXXbpLvOUo5CsGNxUP6DOQvG1rqBN4+H6uqpeS34
TNgR+b+qp4gT6CgdmNMSERuZIT5RAzVSaXV499PZqhLAk3EAg2JuZJs85LTpydLns6iCUUUgm96g
ZkIGVIPclvZ3du6oui6d78/hB8mmlRRMbHq79x7QYCB2M2a5M0Naptm2fw7t7rFUl+ficooNFe7o
Bl1MEBw6D+sqR/I710UFH5l5jUVI0LUiL/QdDiEg9l3eW9s8vdaxAr8xJ2WbumpDbrk9574LVljr
AIZViImrmmjPWL2NVw2oFKC3GgGNrwNI7Q+ZrRVco2kvcxW3PBSKTlDpPNJKoFwe9J05xRv8JNfM
e8wf8elOe7vV2ZUOJGeHy6sPUo2PHLR0bZ8rEjSAXxmpODDm8KoIlks0+FFZQ33uutq/E4LLcisN
FXa18NWF9c5m+/b2a6MSIVVFOH/Wr02N11dWpll6koMvuK1sAZiA3RYY8qPNQU33JETsyYcILlsb
PJtyCQn6rhEtwuJZiGfc4kQ+Uc0Q3Ynycs3uOsqSYkIpxfvLQV1hh/u7T3QDDJPl0yZuCZm4cH+P
eclWc9/QV+WlFlXgjRJRM6ubfj2eYtAMPgGulPLLcIb/JEdGdgu2+672coxhITCUnF4sPXfZZbF8
wnDVs5MXDENuUw6yqQqeYuByS7Xbh+5ePe//S6JYCYoCtARGffOsyQ8/ChyRJqXj4G0jynvMAMd5
I1hgPboOqdunMx5OmuWWSnoFmdaO+ffusvAKoRbZZFoMZG5nvO0H8a0xsFzD6L7QD2xDcikIz187
vgmZRuME51CVisHivU/Fkip52lwDybzXkHIK5snaGZAHtZBI7vJAf64mwYeipdx37mr3BIp9coMA
9W7jKyw9bpzyX+RcH0onls0fK42TeouQusV9Ysq8iaXQt3xUZtFyIT2BODMAPOj9g8tRsxBuBnA0
YEHvNJRmLoMESwRiXO0KnagGpalngx0NhCoWnsIHc8p7fUNN6eIfrsEGA4wy9z/YtPVD9rCnHTk2
/QlKoF5+S7zn1BuwxLXAFinGlwv/vRMNmntQd7Uwnep5V/en/ulAKWD5gJWynEFIjFsOUxaoPbN3
3RLvYPRa2ORmzKZgpMgiF3A1mKD7xc7WVtQ9mDP07I5OGtfgezDgZDFltTuJuePsWFDCLB7Ftnk0
KRxR220EQ37Kuvpf0cFLrS33HZxnxmOD+ufaVsQWZNh0XP6LYWS92YORFpALfJ5Mv4aSNZLmvY6T
WsZSWG9u63Hr3dOCMcVc/3PtaWTxkJR9WqoCBpa3AuwcEODXTebl83UdVQ21W8BuoY1ZlggipTI/
nSdXBHxslTYXn+LVdQpqDyWTS0QCNFJhL1AEBe0aAU6WwLFNul9rRYmcQCQJTkIgEN0cLGc2S7M6
RkCuRfzHfOD1VuakiW1VuKqCQ3/nmQGVpPJ8J+D+Xj3e33qCJGHNG+m9vJV6BItDKkCeuOdZnz1N
UHuPZZoLVoWLvyw6rwshDWCIlFnmqY4IL+7vmtR74cvo3wWXt/YFYYCeR2/O+2Ij4OqyIAVQN7M7
8NJ7TdAD4QGutWE2WvhBKe9pt5wrQ/Y1B7x8ii1QwBr866N11jKnDHVvfV9prPXVqQQHYw0Q0ER+
eW/hZhZbS1e5kYJPss+8tA/Pvc1CenbfyJNXHjfslraqgfOedJUkNkb92urZOVBzIFWd4T49ALHw
+0Hq6TSfFRDQxHODZz6oiyfv0gPYzb3TFP1PUKFprJ8DtOMpNZuwcyP8nJnLksOwtWPVwddoZPM4
JP+O2BQPcOccrcgnecw7ZQ1JbN0uqROZ3K2MX69DkjNHJk1+QemF4VzCebLyGEZ9CvGepAvrfdKf
miYXcSkkb9VV8BhHi+Hg4DKRHkkLhiL1NrnNVMcb+6Kb6WvOZzek5mNfumG/Z6mU6TnBGixoV4CL
8lmUFlRkUYvlluuxm4tBDf0Ec6CS9tLcHncCeHwNiSTtprxx8Qgz8l8RB75qkMN2nzlfTLP4Y635
j0vQ26rzgjKc2yvgStqyDjqydn4L8zgBSk3VRcbtDytcFEe9khMs3BbfEty6uXpll9sZC8EXwLkq
YADIKgvRXEy2zqb6EizDQobB86k+1Vz254dGhGoncvIzXNY9jt8Rhb4TUgQVTjstxXGpb1L0LP/b
/2B1w1/3IkG1dpWZmPro7+GbV5VgaIUYVhp02CcVAoI4SWa9Sneg/Fh/uZIwUuzZzTawn0hzhMg1
z62ixCNsm8f/zC+d71l/Ld6zkjXNqP0NKDlFSyyRqCD+1274Laz4gMcPPLFri32+tA3Fg7XTjxAH
x442Y8zqsDI+oWOcoTRybCQp+EOi64nG17+wC1Gc3jJ0QLMihDGmHjET8v6IyjocxbmGpaQ/Lfym
pCqKAOmpbqgQXx+6Hlyx2RBwkHM601KYoOCadF/LJ4r0Kz2wQuLqcpF9QEa/p7lRaUKANveVXR5d
OCjAayUFWd6kl9BhX20f0DNqTA3HStRwYTxcnM0ZuwsKKfog5YE5v6xTFDp9eRSX93BjUuVF6AAy
NI+4E1OYzIamKkdRyCYQ2ar9h+GoBjhpOGzUqL6S7pVIEds+EAjUPwdM5xkbNM+s0Ma7pWDj/abq
sIgVQW58UPTwY2kdPi1QZ9m8A8UCPeWc9o7vslhoWTCcHebNPLKMrNdlNJt6GZ7r3nCFzEkX+Oqe
OWr8m//0bWHPxCnMTUYl4jU/Ai2S8UJy3YQ4XzVWr+w6Bkr90Yew3IFRSrgqCwvjVY3svRF64e8A
3htDEIWgzfEjpgNzwCL/jCQSveI4v6PhF4s18aJL7fmFk5+FulLI21e2eI3AuG/Y/0k5XHA6zrwE
Fxkp7gXhQyrskEFMu9mMSxsmqWn9f5a6hks80FlfyYIfucPZlCT/AozvljoCBT+OlfWe7cWe8n9T
a4NsWyEEd3ZJKIkCG0/NTmvNVW3a4EQ6cef0cP4lyhbtCo0B5d7+jEuC+3eSSzvvQEb+UNULsMWS
4F0mvUdZ1Kr5r3IGIN09MxC9himv5Y5xdBUBG4iNibHeibL4QBFKiM10BcJWJzP6QuyEpb/6cSeg
JR9vL5+ZPTskrSA7FaH7a/ofzivM86cM3jLUr+KsYcKKu+zXBXggf+HVEpNfBkE951udnC8fdVNt
ihY2YXSn3sE0W//AEDaPqoxlzt5N0pw0DPqVvx8ujMgqaaJrVN/NnrqwHAmrNpX1uw30v/9THvCd
OOvl/XKe4NHdEQgC5l+x8v1OE7F1TlvAOeegBIRwn2zyh4vj5U1OqaJB2Hcb5PFzfDLyKC858Wq8
Ya/YmvwWoH7uain8cK6mrMGFmDePRmVhyPA8vL2q4vdNvbyCbCMf7bEh4IWPpK2bOakNovcuIKEI
KnFZvcGiK0ULFT5uzjtJgs30uhw7O7GhZ9RFHa3usBAKCP6N/GMAqciwc1sAWmR9OWrLYupWbuGE
0BP5OYO8S7S0PiSPabIqTpQabEWJ8w4z9oXuE240SP+XmtZVlH4yVHYWta4XKvrqR0cOEC2yaUqF
93MfgwQqMVXyw8s9iV2+gR289yqmAgz+KQDX9ibiMVqdVSBvLf2M6HAkaYpsnQW4Zi9sIUR6872K
Rppb2joy/Wrqiwnk+c1GIO6sT1gItI4WIitRG9UQDAA/dG4V/UsB4R17H/DzVPjLUqNksT0XDKG4
GTglEXVlb39BLdMOwvWMbaVkdtRWmUn73tBwwgmcoBqRKbtzdIEcelNf+fRrFvhUT8bUmXy3et9a
tTRLIqEbi8VkFAjwcJEd6r1XTDCjtksUx7X2ZAcXOfkwo/K+jG8N5OlLUi5yCl9Y92mnAyPgcYq/
NKqljugeE2LT4l/1XQhIXd8k3yO2FvIRYtjK5arqdyjYLC/WC+2aPV7w4bzkBLZgCdxkWMSbEPcd
I7d9n4mSeWF0EUd5vHdU9hwxzvE2IjUru4XiWedJgUBFWXhu91eLMNG2hpz7gYda9ce7wlfvrjWH
3NTIDIkJ1lJOwt/mGQki7YY0T4TI4SCS0Ep37e038VKX1QdUW5pNu/Nu5hXx51SmGHKT8nCzd5qT
2DPau3JMn3haMrAqszlxih9K73fylo03Gsh5RdXo4zyqhGANwy6rUKQiGTq3CTYsaK8qr+R9qyvQ
HIjM8w0Y1n1yAqNnvj0TrgC4ZUqnr2+Jhz5g/zNJMutbAXQnDItXn8yH7BiV/u6E734g4Jw9e6SS
LyKzn0nON94Fsj8GcFzk6juDw73f1D/Ib44zt4R/YeH3gY8r/j2f8GvwNsDQXTS8VhaocpBngpgn
H98GH9w+FKWrwZmmlUlIP1LK06b1+yBCdwFUKWsnk/P141vDnf3XVU3zRMXFLeEQoPN0irMK/kqq
Q//JZ1GSGuLr7Ei+Hd5AbhxNqPKkKzGqLFkxl/F09I3J5DSgImY0RPNK8VPBjP4GRoVyqD8kaB8Q
bgBPQwspafcfrIAaH+xuFjo++7nfIZVktj9R25OaSG2Gzh2p+kkCZt1z/cNpK02KTr13kDiQaVEm
c4rzz18iBYIE0L+Cx4UeQI0SSaWAhKrQqv3QoWbb4HY3wiWiDAGMk0CLZ6opm9bk/GAV3o6DOyV7
WUEJog2zhG6IGV2oW4ivOiqypkrPZtmSND2HoJHcvPz8U2M1gtYWlkfdDKJHm+dpXa9r4cL+IUt/
rnUJaeo/haEcV19tZWBWazatCrjM7LAXisF8bDcTuUQExolPEk4E8EuNDNCvcxYocT0HmtCxhqPg
GlOkxH1JgxXiQ7k2xqa0DiNE9+BZxVgNQiiIB9ZTvm6iTtMvltpFk/vEzLAvYYFfMBUoI1ALaufy
uN1bCWxHwzVSRADwX1dybvWHsfO+hsXM8SJzdI5ogWyiPu4kwlWaXswTTbiEjNwX9z6zmUhar4wt
dp4Ak22DKhC8gUchSV/x/wQQU05N1ZLnBdUvvQPLKSrxKf1P+ueMnAT1K6ajW/nz8TIVzHhNfvvg
qBEOmuWritO79u3cn3DhgiZhECFbxGLRrqAOuXeQbmjvqOh88DTWLqbvvumeKYkj1m8sQHHyUjBV
gY2nsgscvydjFhCNHMXu0mXLlPkBp2/qtGkkb0wFboZq3hI+tTR/0NC3dHqBMEhEgaSvruRmAC37
HO0TJ6ZXe3vlY5YrX/HjwI6B1MeCNIyyD+I7JIH/F+iyGsx4K02Q55QVcgN125bYHLsFnmtrKsIN
8INqDGZJ7aeXsRL4TtT7PaAsYpGwCrjJ4utpa434+8rDF2z7cfcgtKT+v3mLVc1p3x3SCqn81l2c
DrjbNE1ar3AgdRxitixUwd8RdlSwfSXi4ycArQY6UdiMq1BBW0grg3h5RzcZL6yaCdvbP88iOuQV
5BNBe6EsK9m0Dzu4fYtv0M24cnSJ6KHcCkQW6DYgHxg3lidYQzAi5Tk1wZ6tfsJZogKs4w2xXBZE
KJwYnZPzf2KMpiLdAKt0PyJ5uFAgjwi62MdTwIkIAGvLcpk30rpLuRVj5n/k66f7ulyf66jE2MjR
1Vl1LshrxWm2/Sjg9/6PdALox80O/19Mx5uHd2yjx8H4I09X3XqewoxRXU12YOelY2NQ3Y2Ovop/
vewoQTkRi4L1GAngJS7ndhcJx6ATXp3nf5gE2R6G+9WAl+WH3rKKRIs3zBMwvyOp4EMesSlaQW6A
Xh47Pya8Y1c/MDXHaIsuKNqJ1c8GYnxYGPC1PycH2p0TIXc8TfflD4GtZmdOaMPzx+dgbaV4CzsW
SnFysTDJ9GIy4uTwYG7gdAHscDLzsSklS3BSbL/8iZuzqXPy6S1/BUuCja72afRaMjoY/pcEvtRT
X3s+IddqeqlCMBwjDV8mXG8tyQ3LCTHY3K38tXDfhfg4/cwoOY0RHf7IAmq61ROKZ85mv4QwrRuN
OwhQS1dLEnPeG/NmZY4tX2NDvi+lPw+rKcnWRQ9CfyRb3GyyaY86WqIrtD7ohQp1Gr+zOhr+SBlj
4lpNnaNj10AhlcXc8KyJycDeXdqMtr1CJjQTac/qrtlIqI4KFEAhEz4CG8p2MmI2uEMF0JWV1suk
orgBjriaaoAXvgOYynKEq5QTmYHdNPydNlreXqsPZ+LrM01CxPYh9Bntl7KtYZQNTe0Ee+3XwlEb
qMpTSDaQGK9eaq+hJCm36PB3hqAA5q987AEyTylpEv+C5pMLSvPyNwlCB1uN5haB8WRAOexd9uRf
rTOiJYz1J3UchdirVdDxLgI451UP4I932ctbHA8xVDuqSLC7EyjVTQ8D/v39nrokNVdaFPFjizHI
FNbKUXi8jnPZf4gg2qyZO2VZCFvMHyUFjei9jxZr0x/nqsJTOieVAkaNjtBZAZlAI6KH+gUebmiS
dG3B/u4IH9PLeTWTOXrVOqZ13CtY8vUHhPZTpQdj2Dq1JerJ1lfNgrecW44Dv/AZsY/fNxHhtUHb
cEqt3PaQ40qdpsZ47cKvQMcIFysf2CXteON3KKaP1Z9Bv+H9NAeD11Q4sS4XFEIRGaHJ7F7rKaDF
hXevx3TkRmT/bQLb9tfxOMladTLFMNb20DWxSDZ0Nz/f2LBIT6H2L0UZEIA1XGQnK0mAGUPM0fE4
pSSuVwVSUEA9ogMM1WNfpnp7AG//eWWe1aW5kgKZRyKRNL48Sf+btP+Jb7MGi+s6xCr4rVwNveZm
S7NJ74DYG3LdOH+ihMBT0Btrgk95+7FuhhSDV7C4cNBpFlco9yIcdv4i4oHSX2K2A0o5EA2LWuq+
io8t0RWeU2S7StTpi3OV8lLL7XxEgIqeyWZSt5vJoLahexltIajARXFVf+YcVm2W4gHXTYBwjcp9
1ND+vvu/DVjszbwPMhTYSNce+eKuPi2rpOv8xmWgSzLRFG+1fC0ygccBuHsLPkOSiZzVZY+GkCyY
YVdFq2w/CSkQ6HcJ6m7kwlJHfgoUdqQaEljioaZ9OI0MQ2rz/YwWEjvQaHi79veJ5fKOMGaZebrp
AXac1g1qs4N2j8egh0G7QeAdg2dJmu9YG3wRxbxAiJN85VdElZZbZd8rEROc0GEeTDsgy5ejTiKy
IVJCIoGE/I4od4LGd9gF6juMBhPliyJ2Zo8ieGZWBbCHU2T+s3nGEky1zVm8ZABypOM2av+qL4dv
24TLAHRuaFf4uULcS69rOxZBPyIEPo1l9ufthk3fzovgwQOQY134pEAUmcvG6FHHRsxtNkVErJ2m
7t2751ZT+Odf/rG/GnB0Mg4VS8YGXulUtBEzwZEe/IZ5ucEDrjD4PDdy1guDRcSQ9NAV8o5JHOvi
NrGyqTxMYBNKh7+HpYKyeqeX7dEv1P0NiO5R8AYD69V+/FgoJ31FkuYOs0wN9D0/jgoUzNBw7UGA
9e1jpBVEglOVTEvSGZVto6Mdey/oRu+LKim7AZdFYCJSFel+Vou5sF4vU1KdiDU2bI0eelwvXSWK
sN95KBW5afAJ9YS/mx6SYMJNLStoGq6iAb+04+Jf/A+VqdvmK1jr0jwBZpCmc+p4h3EGKR9J6bY9
pq5mIxp3ZxLAtJfVq6uOUPrWO26XV7OUIlQ4lvYtaJT3Kc1sWOCxzhtDDs99HUm0Qym5U2JS+EZp
I3gEBPKElAaHlSVJSZbsNxk8ejX5U8lfEPpTfQVxtKwbBgMiwnn2bwzFzNXgiiLPxDRHHh3zEZA8
e5X0xJjMYaMMI9kwN1FoFyO3LKO/DaO5j+32DrWswsTKrJTncN3eGS8pMDYfSCQBOXfNPxLBFob9
HOgQobR9sqxlrj/W/Z4uQFSmpkVqLoVNYWlYPjst58UxEsyl7S7eGQcHLEw/2us/Q59PtRsCTq45
p13wDVVHKULgXPvbSfKFzLssCAG69LHTfNS31NTTBP0oSOMOw9yhEzGRD5a+ZqGJvGDkOS+1zvs7
xnka8gJ8HHkurBy1G+92iWHEPJ1zj6Awq/8bWxGNj9hlIUYwji7yR2jSZa27fBRL7dRIoi8kglwK
LRd8vBJXruHLMBs6WNfeZ+N/6xi11WMeVSBmlePaNf47j+xrK8Ummif7n1HmMLlmC5xgJvDIJp9/
5J+CgTD6ZtEKKPG8WICvKOExn7ouQoa+6/UejNK0K4dZcYVoODbjhymu62pnaOulVGiw/bsbE94j
yarIDmuALdGjqMp0TBLfVKESjPAWIcK6sXb5s3ZAysZTXD8qTyXffuOR7K5VKq03coiKNLUX7uL7
RP4BcKMqmCrGnx0mBIP8xC5EYK4155wP0hZSs618qhosIn4+5d/VzShrpYURPh2u7ixCH2FqLodE
ci484NCFOPqzqcrY1hufaCdiRGz+Ei+JTbtcTYyRZR1IrP+499KoVAWURcDaAKohEJ5zdD0LGCy7
gEuf0uIvyXwNVHFSlRbQAkVnV/ELD/xDnxBF0s1FQbUnqTYfL4lD0MJGBWm9aE+8lSlMSahb0QbG
e17n1vSTV9yaIHNczfIX+TGyWC1LBENzOq+nP4Q40ZI5ajcM3moLr9OLhDAzuidUH4LUAxhRsTTn
5odRi1ZifZPoRgjqTRATgSYQgp/z0HgInZFwfK6joNNvgeC8Op2o01EuPDqBV4Nr4pSX+nExeTrm
SQDXHoQUC5/BACCXGmq/FH/JXaCMbejY8IWJTXrxpoz0lRa0KB4PX6sY2lVyCiAIy3hhWBQUIlFz
+HRXiHU796KQQZOyNmB/R4MoSJsqWwJG/ZwzcMTFNw9QtkGWU2MicZYkJP6FySA54guPmZjjKz2S
6VefrcabF7knfVASKHo9cVIGz8R2OuAf8xGeqon35X/YT+BG68FH7MWgxEu4W1uVUC67VNItorRS
RXOwFh7irhPfkXVUkOhmz6RK9da7FD1/kb827j6/t6XPChbPNLHKrPeRd3zR9d90kkyasJJwpdbj
Y8x7I0atekHKHap/Qhwfxu9+USOXsz4t8ptzotTnwBxYTk3+umgsAvzobtLIhdHcmpZLtYg+4ljU
q4OdETOHM7AxEvcDRn1WA6W4gCU13nquOO/eBNrxb5UaamwZrCEh+vBwl5wy8R1owSNcMJf6oTSa
jSD5tRdFzDUcKFvAt+dog0vX4pitLN6LTMUcRpf/8jY+pwRY3w00hqKhe77vwjbGzn7n/lgPMqpj
2p6J0DQeFI3UurF27Wfv5oI1OqDT+CXsmD7SG3oq2p72ESnixtnyQPCKK6n5oc3uL596/e+Yy48E
XiihwS/mtgy253JbUKSwkWr/92WU1gDO9/9DYY7tePRPzZRVe6P1T7g4Kd9xStaU2QvVDf/RYI0Z
uI466o3gSRekDg79d2jU+pmmZyQk4rBy+Z0YeV6VcSZC8Z00yLkpXuSb76Spk+4RmNwqzNx/Zjwf
UBaRBquVwK5CgPL8+K1PNdoo/yhT33k0JeZrF2NdCOllM69dCJLhrFUvH9Cz9OYA+Fvq2VtvsRjh
aktbeVt4BDRFYfZuYpoAVQcxzE1InbgT9UmGzeXjMREEk/TU8EJPAKVyi0U5KjYM5CxpI2mkjQXZ
qL2cfB5xIA0RZLHjYEfoQrq+I7X5zE+JD8UzPsxwRVGQkTUrtkmZ+DDkqqEBvSahnRjMEGA1wCSj
KBFFoZHO97Z2CAWFr7kk04ZT5s6LjDxB1tSkAe3BVEbOk3WsHnArfeAY4l+nq5mWoNdT7Idz3WR2
EmRjnrvmcIHnhttH2odLPJVoh0hfHXBDdsZyL1sYQDF1T+V9LvQ/DdJdDQqISTMJ2Vppf0/CYb4z
ElccdrNvFzhK0khTEEOGTljPP07P9RfsX7fMioUHcxBheMn1ipe/uP7RWq+HlDKmFCY2mZO+CfiL
ja3nEKrnWpqCxO0EpyPFbHWDyr/Xbqp6gI4QodWKwyk42aXuUDV1NqRKdck92sdEBNTG4aJphBIt
5t8N8MizJvWAHAsUOBI9N5AzUpEONp7RtOsS/brwVKosH/SNV80bimrN+DB98ftZxdCS/RvAsf5P
2dGuWOPOfh5xDiKSUw7CMyXQCrYRHqBf6q9AyoAGKWC9aeHsjbqmP74mHymxGiGee9dBvM1am7ok
+78B5T9vPRButYtJ3XBakUVFqvR+uawIueRJzDTeWUat61G9VGEzuZeU1A957qv/kRRcthHOv3rJ
n9nH9j9A0Qolfa7gNwi1Tm5gu7foZgcNB9rEaeSd8TCNYGu4BxAPSgyhKWSZQJm4KW9uD8PldRjv
FgHhLL3wjOHf2vDW4evCidV0DwK4MZk5kWZuYt1PTzNqRhjQfYbFu5z6wjmuQE6C7AzGw+2K8mzV
N3NCj2PpFgQX9ucqU0n7gQ3tEN0ylP71m9UaSTwNr8wmXVjB68mh1WKPaLBPBOObZZcsiwtmGwfv
UCh6ub/vU3PLbJxHwdxf+6DMPn2nxmPWZmhYP757Ppa9UyXL6I/rLqv0oGdWxs1OIC9j9fPq0ynK
LDCWxofB3Z87hcwfkNgySoRHk3vIncGRZUQHlOZ1cAj+e+628cmj7lTlv1CAJWIhZAv34fjJ7XoC
unazZGBecea0m84er4S+VJh2ZTcLHWeFjyTyclA8euFBuAUaXtsSvvcnVGKvMaGIJEv2m6tXc6IO
B2ld03sFgLd5an9LuqBVYt+OPTyDpjccGmbe4cttdQwcvxjLO/qbHKFy2UbpsVgAIb86BZhMGei7
J3AKXgN8RcfFJqOHPepR5rek1SdCt/kV92TSs/Tvdi+PhpyjyAuCQiCQ4Fzlzqhwi0gm6NzHfNmt
cvcrvY8ff6c2wjtGxE4PFHQrGTJ/buJC61biWBCkPXSKFKl6EGXHcaQ5A248A91XkUMwx6syJu0A
6l6fvJmZz8wAL8mzn/HBgcHXgo0W6d2rLUkYapgQf2Kfvz+7011CeOHFnMHBF6qhRbzGUuI7PSTr
TzIJrfYpJo+2k0OxxrQm2XYK2aUKNWEya6XRsI2Ss51U2LPHlTver2xin+FwILkfGRUYRtsHmODG
4ZMCPi8UIweE8R0wzEe9xcZYvs2BsiIclODrypYKthWwuaHfCo+vxeoBrPhFFKbD1uNL46bU38nz
HLguRE25TK6wF/EEYvFksE7McbQzSyFp5+ovsegGBhYehcrhFb/osAt/prpJpv5SDZfAtHt6YH15
uLLE9ZEwXhYMvRkOHAEgP8wHZhg60po2bW5yccUt986EkXrqcxyi3RWCnkK2LFPvWcNgDhd1AWse
R6DkW1vEYiyccVS/1T5JBNi7fmkxyNne4nYLDk5oSRh3hDUmihoBYGn+MrGjuLlONm/nNdV92W5O
M0fNBaDaNH2/wk2trTFg7uMaLrKthQR8AWWARgyVrV8xci+6VKWI5qoKgj8D7ewcVnF2M2mW+Cx8
5hki8N/FH1uURhjqugHGiJOzl264wmoLAR6ZXl6ShzxpAf8zL7EoynjSNC/Ndi9RbbFVZsVKRMdA
xDS2KBMkEllLxp8gP+Bs9SwunYYMpgPOIMiCAQ/hEDTFD8pvG3h3YLpQLMQVdYxG6fCcN61MHrNk
6jMMVr5VIWySWiTnq9M+rR5yzqp+h/6KIVXa5+VwbIiuRxR1m2qVJB5dyXQu7mZeIYS5RRu5Lwdl
wyuY+mhc87CrlbPO5Ob9MiwVKCUQdIiAh8/vzudKN5R4yjMnZYmdTl/tTvm2jONty/xqdfeK2dUk
RZ5XVoXFIxXsYv33x2Ll2DRkUguoyyuuvDjxwxDCQYRCtdLc5V/0D1JNH7L4OPyfpNP5nZ4UZoB3
k9bMigf8agPBu6JV9tVQSS7unfu/Vfj2L1bFWNAOpoZ61HRAn0XnSPFtEL+nbeNHNT/H4MAndykw
FJAS7w0NY/ilzafl4Sbu/FtfhnMzS4GOerf7QyQ5CaaFIlVprv46PmUf3ohb0HmyzVDbCTvg79ov
nKquzjS9FJqCfRhIQdoY8MPjkLaz9XcUbzR40nu2myAjZ4ZTQsDbCQQJ4uFW86dILzInKxsB79pt
k3I0ABedo9WGrLgFJwqGLQ03EARwm9R54tG28XjuZBOVN5GRdsxX/HDzwWYbeKt3I6kUIhAee0fP
wV3EtGtaHddNRd1rTvETngSINkeeWQKPbOeS0VsNlfKdS14PeFu+reXhD0EXqpV7gvla2pxtJG0p
udLKJ5v2IkcYu2u12IWsDDeZwS64kWuitPO6tUfzn9v4eW+dWejx1kYz7h7T7olItUjUVUu6pNKq
LkstJfS57l6kNuvM6/h3s3cmpQFeStzPwCHYXnihJw2no13LZihbXHDb+5hDWVyMrsQFztZM95+t
3AGNFCyFGLlspOczkB+GeSxKX+0lwVMouVWoNYW5twOgOKB2YeYEeKaKuL5tQ5bKkxdA13esFTm/
uhHyiTmAsp1yXWOYNkn1hDTCKb5aam0kj9YPBl/ulKGsBsL++3oJiDvP5pjfik5qdwd9ckcq+M1J
oD66KaRPLKRU5sebLaFbb2KhdvYiXiqIxbgWiXOQ9cbl4LrO4X7+0QVsNSLAqtFfvKuJffGenKqK
LQyeGopVOwQVXUp6dO0HMBzz11QvA2w0m6NzpyiCC6bHEdI3NkIJQnEDGI0EK0GfebNlhhI97Z9a
n1FSeaPPaPWHsUP74QmqUAg9nILtzjPnrL3goTSwEOvAAbO7FtwSa2pJrtx2Y2Hlx/sL5v/a/o3l
qP80cXXrJ0j2WY3RQgNza2O8dhEY6ThCtPzALS8YoGZZiy4dDa34IJPOQYRYpnUA1/6vCMG12Mqo
xKetW4/EkhVQ5LVAXT2fNs5PVvk6Pd3vdUo2tSmRgla7RroaLNoMT1+zfUw/XkiIBs+QmHgBy6xG
fTl0Z4u03okG2aEMKQF7vwim+Bin8bAmskYN3LvTE44lAYzpqx7C1Eb++EXNw+xwFtZhgJz47M8Y
fI3G6ec40DQa9VHz1qgBqqiQGaj3JtwLBmdn6WWYVYl1yvjjRiJj43DYUYo5aB+P0Qt3WWW7TEZK
zGzU8OlKL9rv9yNPbBYKASZjekZu7w3qC3Mk3gR2mBTcIoukYrbejzG+29+YSRzPfDtExsFCdqko
RhcYw0ELWAloZAhJHTD6tpE0nSynhMnjdZ301GLwveJoeYrGQ1PBLp81wq24Mw4p16V93wynAous
HmEnVLEPqHaTacW1C9HWfO69hxV34HTYgb9ZqN6Kt3Hpg2JCKuEJ1ZB//3oV7m4eONigKbp+47Vj
c/a6yLunGGh4M46qYOYlJj1F/IoREK7Q9juuimPYNZnTpCLrgFqwd9cuhdUd0lxhvsYPXR3dwOlW
YoTaJ3jgxADxuhjjtf7rHQtbpgfTUniq2FoKpuu9acmCQfYO8HquPI9rzkDg/m9DTIU0YBhhaUGu
o7xHQjdlLy3arxAzhfLxeCoGqDJAm9ptJG5RuAQqCF6gXh53BtdscU39/4SzdWiAGPu4tkFGJAqC
6R/bY2wEv9oehUNMRU2tOkR/+ggcgkTV4PJndMjn4PV3soL+S0AI7vkgBVUyiDrGDUnRSPLitVqW
+o7Ec64KQhh9e6dIhTbdU4HZ6JqPB5DCC8y/vVF00zmJzChJ2rIwxQP9RVazgIrYABV9U94vgqeZ
ZlF5ixkVOjVGqXN8bB9g2Dp987xDRYBNoIx+sKAatcqf3PLkbUv32evU3ssyKAZNanmqR5WcWyf4
9Y9m2DYtRtlLctbNjqWFKmv2bdE/Wg2Mw8U79ZR6lQZlISDajfOjPjSgAxs/KFdO6c+QyPetaVg7
Kz9qcYQsZoAkeMx/YNscYhHFi5NvfXSpiEWvYU2QEIcC8Mo/BI51iOVkSApWpH9f+bBuLuOKCD2X
w4O4GzQ0FjALnLpaUP/PXNpFO0SnOjojVfWwvP17tJ/BaL6uTYOW3/WuFfaT/rBaKo1qYAV5MlqC
0bdOKTLkPTvxdw3HdXZ4p6T+IakUXtW8xOsedQxCo2yV1syaUIKohI5Osqkqpjg//f8xwDcnKA8B
+8jcz1owc9112jOprMvL+4HfiuP2B2UiMu5ZVUGGvAss3m3T3VhTEF1UA2c8pZZJ0e3FwHpGhNUH
xtUU6k2Tml9ynR260zEPwr+Djf3hgWkLCBAS/68SR6rkPtjTbMGUGYNMlitgJ4xDbXg0IWZ0kHNt
8QtRHXHHpNk3IDX585XkljIY/KyCScuEZVJo0bs2EvmtqDc/miuaG2NznSLksNRvG26/aZAnxnc9
u07ikxU6q0JzItaxIcVnZHJFCY7SE3dqSVN0naHjbpNRHjG4Wph56Y2VXxPuJE8CG98LmKE1ww0H
Dw6kM6ypiGIkdg12/EGx1q9ty5o2UMZKyDCt3Qgu1m9btPkb2s+UMVEZerJw1LZoy06h6wVJWvpD
+SbFxk1fgQG6JNvpEsMCs6q+LKqzJckwQJgwKPTEQkl0t4KJ2uw+PA2QmrnAL9L9bvC52No0TY4v
2gSKf+VuJ/Ft5xHFVOBi5TU/c5rnwkcaZ5SpaS91yDIa5bzBgCUVR/qZPYq0yL4U6X5xYUIYtqSh
22L5rgLdC3EHoqphUO78XS3cYUsO4oCYb4gd6lwshpVccEh3awU4sCQ6gFlrefKsLi/wg/5fZrER
smySktGq03XXzSyK4c2Q0rtf6+OH7UQvkMU4s9300gLfHGKvNaEZnT51Ml8tfCuPGX/VzgWfVoHR
s7cXIpwblHPdUO9lGh/6Lzbqw9jo23T21JPHu63sqe+z2B2EnYw8VgVnUyXsCr+lBCpHXW6KcHc4
59zdb8GHxUKTx3cxONybuCu7oLfeghT7iKqynqalkYl5nNBByBo4ZuYIwJf+FQB7iKa3tNZvgMNK
w9Q/NKZQ6Omk2qSm4TZffWU6/8mrENmKfAPBpOXTBDyJ82WqzG4HbzCm6It4eTQBbS0wk1+EFJC3
0v5u3zvjKpVD9YFq1ShguXwBaiYQUMJWbLFv7B9ibc+i0mKXIAhsbxar9iqqYTguiAkBG/7vhhnV
dax4UcPCV1/B7soGHHxnWgV0jHXO0J318TtsQHaOxq/Qjf8hlGnN1rs93X49NR580hF3RteTuMEn
VAZ3Io9HHVlzmEgdJiylCftcZteA6cg1OxViHeKKTDtmolWDj60xt2x0JtUJbiKV/wVt8Jba22Nh
T9voOJ2S5asgC4mt+d6Qyipbl0DDvYG47dFMmlpaj1MZaVIn1oeQM20ut4MlhERpnlMYfrXfz3lD
uRuMalC2y5z866aClfvzheYpD9gX8V8xGOVlNNcvPyp96Z8DO0OVbUac0OgTSdd/7YodvBl1Uq+Z
n73okudpOr41htcKfUDkEYlGyKY1Tgzycht9m3WANFnMwP8+PCZuIDg7rZGfN06am2SDdAWBcyN/
Y4ASuSsdKhInyvmIeqdHUTPf7BXHsLd9flFGHgcZzF1Tm4rYXv1o7gJbbKnpwFeAO85iPuY4947f
NIvLfMeQPEl+EQo977a2DrYOT4BKJ7AnXEVmWATYm228pAL9vgeuF23wFXhdJmbUFNfe7bpftR7Q
YhbM+ht8PxWCCebrTUyW/h8EH6ib4+L/VuxLzLITskgFmSc3TRmRwHShC2dBKeMS4365CZshGF/9
/BG0qcYLC/W7K9O6bISvz/ruVdQgGXrF3pnhTzvv3aPidySLD9SZCnsW2z6eoz8qBxT9x5hextLv
F1O3iVGTwsVZvN7tXlL8FjyVex+aNGUiFqhApeNBkWy8VVXAFERCGEHb3P17kV/gWQYMuw7QeQeE
yA6xrsxnpaF7/8CKRBTVfkpkbPRUmF8E1uzDJyQWoqFBsFfZWr4icVCRAnp2nAgVJ7vbKVo3wRWN
YMdyYW/ZZya1rTewpUf2iqMO/JrEUjuugE19Pw9LU1Jc+ZMfdc6DEGAuUqwAbIHlbNDXdGse0V3I
RnOdwoNtYH7rtBSJhQixD+6jTzGsdMBUKZ/T9wt69go2JglluQAE2pnC4rGQGsE8fnhBCC2n4wj7
VNnYzmExOW8ken7yb52879SBjBIBpcUG6cOhdh76k2nhd5fEjupzgxdQsdu0FPQMLqs5cdi3+ss3
p1ksrWDb9hJHomxJOKzDfmjkKxG5cqG2i/oOyi9rW6HKPVYqFvtMkQapWQWAe90RuCPqRmplc0GN
o9Q5JZmPsTLlvidKONKGruqXu22k/IkATFnwZ6nNV+pUJAUShruAJ/ufdHJt23wdf1gB2fE2wfiu
PI49taS2GiSN6PtRKqVM60KT06UZNp95i08pwHG1HDVCJFsLUSCi/4iQM1RZkcHuG1j3EfLeyLsc
Og9FaFXDcQglW7PaO5cirtGv4Fex4QB7P4xDIuQcVaGO8TCOXnw82BdsXIgQIVBp2l3ucW58olx4
tyjbDZxuwOm6CVLr5pWxZ/U4NQ+WF2N3zvUIiDn58+3NwHPHVaxFNdYZxvJTQUjkh0T2Pjw/ezhq
KNWuuG9pIPCoehfR3p9r7JxMu8sh+wTCI7WqOzEC0tN098jPRd5xqK//XxOt+gFEZv6r8fjvJ7pk
/Ikvrw7q95Gh+66NPiD43gObDnjvJbCs3nJH6BGSAjdUfD19uD97NrbOU29Tbvx9WB5O4m5brRvh
nLKKLZX59HMHMjDXjhjdrZRiiqMq+Z9+/xym73scFAROpxkRGEssZZJrEjkJsvvFDLbBGweGHbGF
3Xf65PdBDPhP/WGu+gKLixy/v2iBqL7RnJRdFhyuq11QfsoPUvj1fwyWmHQbwXFPKhZmogLC36lq
G5+hMYfj0U7aqfezJpBb5CyV3FDGVnrDmmj99XvmFh9TajC269EJfbs/JoOsF3N3o7btJ+wifoFB
YH3oyz7tW0COc5UEw/VnLN27urVzLpBv+kvZ43p5+J0d2Aq1l9EQo4mCzcSV49ZHwVVvWB68eK6c
3NhcdCegIWvfNW8Y6ZFNDdYENtzIRezY6+F2JV1/x8BfMST9OzOiTflpk6/Qs1gfrFvpzU6PORK1
HjeqqME17mABI0CbN7AAcJ+AOGUpl7W2KRAM+j/dX0Ifue7YzK20doI/zq+PA+7WkfiASiLsC9ic
lZROX5JghsEm7djZvZ7zs3oyLyY28K7Gh+gibKOiGgzAxb0uEggWXuajL3e5t2O6qwCK7gZgNLFO
QkH9DpIleWgDmudomwA5/lqP2z5jNegIaOs2wa6XNdnvzw05G90mZNgVL38IdUn+4jqru/gt+Ob4
cSbC9333egiVrl7f0hYEHlMTOO9LIDxT99WHxT7/bdQu7r+PzEUN2yTpNNiFqlHD4udcXJrugsdl
NMdpLoOYAO4EFvFAt6LhSASSnbNP0URhCsQiY/aGv9O7oXcXNmjyze3yGMTVelHmaG/S2U6Ud41w
7lTQZMjcE7jdXBfZPk1e2nXQOQ2mE9ymO2WEpJoROZfZSirjWJTQIeJ/TbUo8Fw2fkEgC8uYJMSX
uMYrf4T0UMOxUsI6FAK+BMEuck/Qy8XvPlejQU0uou/9iC7lTsDfdbtj/uFh0JLRWrdWG0moyZru
iBBLW/HUFTYGdGdl/YfbhZLinStaKr06lrrH4qeBi3nOhfbFKS+OLYks4quNiv0lrMhadj5DrOvB
54U0lYyegB2FHYLWiyqEPOMyGAHmbxiiNwybEqBux00eFxxHwFwZfi3s1Cmh6LmLY8lF8og+pIEK
XUxyxZF9Y56PuSRfTsVuYBhIPdix/0glUHemZ6Y+zliPRcvJfTYjDtlkJL3vlW2YaVuUsaz7kyp6
mgQECvZ+CeQDY4uOUzGw/GHBjxkDHFoBCniN4mWDa8rG4h22ajkT6Skn23ucaQplbsuQ1nzQkNtO
OGoaeo/qzPJ8F7h32BlCi7R0t71Th3dJGtHgjjCDX+btspCNhaVdciQ1XccRKg9U8YLPlgcCcp8C
tTGQtjwEcq6i+r90cTGUvCe4OXBEIFq27sLQYAQfpY0Glm21nDRMbkhhCCaJwDtEa9OLTk/yLtwP
9ieK7b7VrgegZ+hXMGGGdvWkXvSiEYLAL4mM8JyBA7IjjEEU4bL5Qy7bViIG5aMtyjgrHwFEaZX/
3vw5uwqyVdZfHtcuveAN7CAIiplsjhF2vymKkC0ip+aGc/X1ynHceQ0+h2aFZgiCIIZmJ8V04p0h
VURhPKvpPYN9mT3rGBRa5sg4a7y0CLoS+RWyIv0i2Z51buZ05Eh99b7356tq6K8S8BwVrCmbQfEi
MFnE61jOkZdwa8gWH9Gkivgftsr32+ID1uIiNWzO8eORHErpBw2FoFznc2jzAz+8BsMDwscLhwWM
InXU4cOUdueoTI3bA41u0UBqh8e41a8lrNpH4PYgrVGGIU1fwp9ssueeSXyXZ9Bw6llmSlnu4Wyd
vL/p1atw9r+NqOUMCj51UOBtQWy7ByszFVkjM4OztkX1t0rciDm8NZeSdCUuVIq5Z3I3WxlGpuJu
zsxLDJ76uq5quuryqr+EhnBqNo4BewFj0Tg48P2ITUVGzwifmZQIWf/MOXvsXZP1GX3mxBmUB9tC
kivigwQW2z5zKJ01EYtUipWWRdWxoacDdjrzy4BaFjHk5X8MZhRhmly/obDEeAEp0XSlEfR/sh7A
YOxOG3MFQI2HaLDLGpyDh2AE3n0jWn/wkCVjaMARlkn7SxnAoYODQvX4VNvqvVeradaaN1LsBkTh
Ssm2wz+XB/wArIbskTPRbBOIaht4vhxcGPzgIR/HajqZGMx0DG9OSx24etCPMQrAgQC/Qd3MkAPd
as5a8MGn/VS1/vO/jV3u30yiUsMTvegztkRBy8pPbyMbJvgmMyTtNEnqUfwkFUpYhbZlXjOtJxxk
0SIejIdASmOlflrSfVh7KPJrPCJvg+bnQ7QHmZG+9lb0pWMdvOE7zavHmmA1eJ8E2wqLlnVKCju4
NnG7IH+fvjAOMmEO60FFu7VzJYIM5EO+mf4Vv2Ufls/2Py+eZ322rsifYFERCwLGAV4hQq6M+2rz
9sseeB7KwCHsqNc0E+D3wnLA4HPc8XNM5k5BMpjf9KKQ+aWRmRWgi0PpanXfDFdo8e/+vbwzwgAN
KnqE4dRW8rf/mc4W7xjIQjGrFh21IlRW91MWNoUac0xgwz8c18KOTLZK0JO0tgl0BlNsoXtfZtfF
uTRmrtTITTIX1vNooInInJF4UN///gV5nxB5/3mUXchSZAqwbkwBShpw2RS6ZdoTF8JpKz9d4q9H
2CoAm1O+k797BI2/KWfRMvmTGerCe36YOtvR8hA8ztYy+UfGJQZzAtQkmELhIyWZDAXKN7QX3Wzx
7uDu5mwm8Fk3zacotrNI1f7ZSN1ab7C+sIJZj2TJkToCQP4fJVoasuPptRLCXaSjSKXxO7regWcB
BMbdJQ4Pd9M5z4s1g89gPEocJDK2A21c4ivVeUVTbUxfrTltnINSKi1ljrUor1VnJmtstPM3GJNR
jEnPne1K2latc4M+lmPZSmrgfnq3hEzaZI3IKgbfHDQQJp2LZ1vRJlHN3NmXBs//h3cAXOQOgZA9
c2hvhXpzBbqTj7JY11aBAcVP7T9VZyCWR4/ymzm4YMxq10pGea6Et5MDGXcuHmILP9XMQ5oP9apj
5b1I8rRGOusuCzL5Ii/zVB3Uo4NqVU5CXkKY4V/2Mly1pSwY7B/7/rwEoT29DH7iJ1eStSK0//ba
ACEsWsntleJzzvz6/IhdoxX2ARBqQAcFprxWs/BPnND8oJhjXC8aou75rh8J7eLRyTQu4FwE2+Mt
Rbu9H5x9ZtPNmZJxxXp6biHM5hNJhkKSkBcPHTSrNpcMahPE7KAmaW0H8EhOPh6LPXJ3mGZwcfGf
WJ3onmqlR5NH0PmGaw3RLPwF/AD0iYArCTd94W+ciQ1mzX9ZCFq7skKKz7N0SX5C5FxuX3iDArLC
vOltrhXBAgn0DJq3asz1ZsFrRBDh6fX6oZSSwTFft0QX334mcIafnWMH0ItQuz9/jD8SxIKoiYwk
ZdeE4MObVq/PDHM/G7EQihw+oUwr4fwg+gKCTHRnsnHAmhTNeokld1iupHx3o9smwn29gx3ItHTf
0L1LQ4LzldA3sTCmpHFV0BjjWRuc6kNbczrsINwn9ndxnKB8NEbN8QFly9qUAIemgzwodQxeVFr6
C7vT8Pa77xY+HMMj8eyou0heXPV/MLhF5XqcAHl8KHrSsD0RecTz7NGoj+aK2371oAlsY7tI12Vl
4I+V//pMzcsZapgc70ybGCmzCFuBqCYuXMCC1Ng9NEKsBBYfdrFhxSdVhhhQyjWVdQpYrmXo9QFH
ExCuAjMcBEf59eNw3zmEo0nDDKcBlD7cckPl9jrH4rtBvtLHzYhhsfeSU6QFflWMwvpoGt4wxOxp
qC0kDYRWD3PZCZsYC/2sqMSBSebe9Lkp2hjdlyWOkhB69IrgmkGGM4vlu8RC/32OjJf9MqoEeJsw
9Ofh5F/DRCVzaEF3GSqUgoSVZRmvQz1a2ONMlbquczbIbN6VbfNqXZ3F5AjFssHrueIifZKg9dgf
VAfoqOCSvXVfNEADNhgO2odOyKTn5HOwx6cicMLrNF4XQtX0UQjZifyA8UBi5nzHxLYhBKLgLaVY
Oo6OMUqqmVitz/wsttlX3//+IPzvSNBiIep0On8/t9O4xtSgKwhJKyw5OHHtrRVqimVdlUQclbvs
jKQqfV9nj7B/GjS9L2CCb4eAjA5+AhZM9HrpxPY3uGYQOtu8Mt9AzuxJeIZ+Jz6lqnnRUW9iGSOY
/PwBMNKR6IwhOgaypTDka+CDN/i8m4wxaL8Ul4wZcs90Y3o2r6sZbd3+BPEAjhXLaDlB5dzHNsqb
ST4bsLyuOAoaRpkMIXJwQLIsPPbmc3777YTVpqB71/hKbbLM6lB0RxK74mxOXG8Ylt6ZThPvITuL
TI0j6xTa2qLQSf+9phh+ZxN+WJPk2TK9y3IUCkTurkaCL9S2mK5eLQVAwn0t4fjWp9vIn03H1Wpy
yRiSjNAQTrdOXcE1MxQEyZWRfBkD3A4HyONfl5F8pjIRPRzUdEoK4zKimEjrZ3to9ds/J3UlY64A
0wJzAjWzR/ykqN/QlSg5nBl5bNhbxXaZ/0WmzbamzwxcYdy+SD6alXKLZUWx2zHirM2qYxG2PUQA
9vrOeh4I7h6tUnPS/SdyWW+tQiVXeg23ZmX4DPjldwpdN85gocEIljOvfS+ey9xw45jHa/fMF7sl
MFIg1azLIHW3H8P193GyvnYdggTzUIUor2EXZIDpIyNndqDK3TkqZHkN5aKRKmVQfdFXGexNjL++
6yK1i+SJecj7Y/5TD3WQQ74zUXD6snGVTXrIiJYnkEXc+G3a8NdqW5gJ/kroAVBit6ocIsegtb9O
xOD6IKEt9ql7hL1iaDjD6FLpLskOnrM8XCfcC9y5IsC1c46+UXwm8pcQc1YTtRM6jPHnVYJ4epSO
xYfISUc6+mZPmQMEaWlPWvGINQUhnYrGOWCsanPmQRjJw0HbsAAcC8xPLjnhHVU4q1juE7ppQM94
mXvkREYTz82hBnC4JsBsrhuJ2XQpGzLK0dO/mtN9tN9gyEhyXc8oC267NKMG34gqrqk9B17uyIuU
YjRIotZYGj1ctkwrdwmZBxf7ltz/RUl2R9XjpbWOAWTg4F0BqyQ8InPN6JjwM6y8WbYWrA13QnF3
YxlYZn7r4BA+iiG9t4cFQJHOKa5EsBYqs/cKHj3OyrkTEqi2Amazb5HTtB7LPIWuNe3ZigH2ZUxg
VXPF4TXFCgTxMpw9S7AR7duacBTxSD4XbNz02+HoIYo2CWlJCYaDWK8u7BAz6tjzfsVMFEIJYadH
NudWXt8v1XP5QXyj5GF2Y7RmJ8go8W93cbK4fyXsoMzy/vC4nWuXaj4Kti8crawXFlPcUA6GBQxK
IJXeG2TqZsVKJMCi8JHGkgU9q0b3hCZcQlQdovxI4tDGeSj3dmSXyf02pJwu9/o70lgvurn5FqGa
WF1C3uNw37nqcg8iPi5kLwG1zfSMe0UHlfzeNiiJPT4GQFIEgco2ut4DU8hevjrBYKXQDfUHpsgu
2LHdFRtZJwHWZ4+N+lJVkeBYrowdcwQryU4blvZhqCd+uhWnP3G2ijDowFFHPKGCymM5cnZ9yTfu
bjCMMnC5BtrOZXtBk6VA1vCSOfLSX+GSm1c38vhNurHAK56ePlAhQHCs4Vt6+CrqW7OGFBsFrnj9
Orv/2llHNultwyF8UCffcDurDRdcpu7J4JnErMBEyw/L9GeNjDzryFBA6kOWlfERJGOIH/H4iwVd
fFxewbgXxT7LxOaw5kBFU3kp1DwVDVeA6gR4EvFXgXvrbfczM+HLqvLh4Yahl3OZrqISTSe809lY
c8Uaw2aFMu//upsDrX0v3P+rR0IZVwxoT+ZbOD0I+mSMr258v+/FQpeGbHOOiMTaXIuxd6OAzGYF
i4zycCCwVIu6Dv0vk6isQDvsylNLi64On4ya06ssnUJdt1j1EPEyzRYKj6kNitLZH+zrf68JLySJ
x0BSV7uxcof2eGje/3gW+Ad6ttjT8j1BT81p1EbwSUrRwube+0DS22ln+izd4uQuPIV/SyKvf4eA
jINA0qKLiptvx/EIbcO34vi6qbhG1+BHqvV0VwLW79+SmjLD21BbLuB32G79a0T9cImg8k58fFHF
iqCokOEQHSmrmQ54gV7qdftL3GQHneoTQXpAcGIuUDPihJ8iJiIFtWywkaUMhgd7JBIAusdoaHNE
jZa2DJORZELL//8AoAF5971H/9Hmn8Ix7VnLpzci3MehTPaCN1bke+HME2WCZm7KpCR+LgGNhcB3
Gg5vTko4y8SA8U33KVBekrmlOJIorJ94qfO/FlKzAZ4fCF1Uz/fx+8sedps+7tEybf/mhDltJ3FX
uHZWpA0MBf45j7CZ3V9tQ6U2XNUpFXm76UqfE6pySQYU0stvgnKMjNunSrLmQqr1a+dmxyysPCUM
aCNtfS7ta1TEqWrcTS0IfjWWxQHIEeVhQqlwg834yX/oackeawhgqVqgNHtT9tpt3SjG7wrd8wU4
xyauTl1W1gN2uWuOPkeGX7fLtUbdqhADs/0mGWjJUpkFrMVO3x4d8Tv5a52vXWBtbbrOQFuj/dbJ
cVhyZCAAKN9SFTRQtvJorvEetiu+ucAUf3iTNkPUB77VGlyHoL5oc3rnNQ7oviSKRTu9l/hYiY5j
LL6oLm2XLO4OE9UTw7WIRCIRm/6fS8Mn+iu0ldhtUqX2X2P8JxB4NkBAn/QMCkXRpdMixjjTOA1o
hPJdNd8tJpzhKdKTmYKhInx/5IRgA1g9Daq2pVfqj0lX+XOD2khrpyFGg8p13oiIUpSimQsmvddm
ZScjFf5lEwKGq06O/stC6Zxi8gwzkmLubLLDawYPfFeMKIUkOj/43RfaZ7TDDBLGJwGDa5b7Ej8L
lAM7PB1qwp7M1mja5utUxF0uMlLJgnM+cYzB2WPSB0IRDYsy/T59OuQ+/EiXVDIh7FSf1y+moNXP
5EKYQvVSP1eZDc85Wt7L3FwIBN5AGomvv214Ejm5IDCQtkvPkLaruCKyeiU3WGu0twQIEwabqm1I
ZJ+y2AfB7UlIVww7TrxKCaJoYp2MwqLzU+McwQh453FbVxj3v6bPkEYwkr2vjoXY8z3IOPVJlRG0
wA+LNTO28pu7lcm7Ml06+l9Qb1nIKudVr+7tjoCFi2M/s4HBhJ+r6kHCpvpToWd/k1GWfC8R/qnu
iSAf86FSrYXvC8WOESKSqhqRqsjZg1jXRlFM5FMc1i1DV7YOecKr5J/RIBm20mv9nITsCOtsVB1v
IOFdxgnDgAAfFNJKrsc8E391rPF6fvgcBAaOLM0EhZO2ww8sA7hVZl0K0jK+vohOcPz9aiCy3wdR
xX4I46kxQil6ogARtNZkGt+5bqJZD502BmIAK5g9AdhKJacn1xniaE8CRA/E3NkaEqkyUlr+pvdC
PF4LHHvjoqm0uemXP1k1wa4iq5p3TCfT8wPugHBJffKJuv6MO7DawbsGzXoAXqfkSStTFm4CYExK
H/wa9h3R8B5OofKReEBwuIbdNUqnnjznlhelLJCHq/pFkaTNWNuQoy+UPz0aghJHDguLCT6h15bq
CmSFLUQqj/Jaq60GMoyCjxOGBaarpctS4ayD41EWWNCO8/K1nso3sagMw29yfUyevWv4/hSMetRd
Y3lEoUKoj6LAt4GnJzAXW6Sm+jcBRLndXdADjivN8VL0Uly2Tmu2Er7IgG+GHQyHsKDKON/4QgT3
ver0tv2MYUjzfSHQuvyLF/SleXHHutZdg7oU5xaK0BtO+i+EymtVFW359rblZd/gAijf6bIDioI/
TAq+hxIPuCkuQVHECVyBJKMP6mm37XCkou/rM44TiVxkL8Q+6sok4rIE+VejbeEg1Yt7CE1IRp/2
vDoKex3fiVw+6bAQMKfnpLD8SAdcqZUWH6p045J7VssK/8mao95N8XBV9dx5B57Ka1+5nbKpEcMY
ySmVFv2CQ9sPXQsiHR/FiKxhcSfScXcZToF2VqRLb4CtdYZmqt/wPSiFo8W86qQUJ4EockXqKK1o
ojVxrlQVpPljpqSmxsstxBzsPWF75eYZiVDS6sm9R/JHw5GtFXvPMRxmAyWXKfpHuW+tujGfYoIl
L61TuI+FI866NoVu1lV07j50TzEpbamnb9D64upGwRgesNVdIidWB1DJ0MCb3bEyqQ82lYxQbk7K
ekoiBh6hJFCTT8o3mQKpTUPn8Le4aiaqpUyu/ews6lKQffg+DOKCJrXEUKrjG6J0JoeRa99HZV/9
EMokOnUhWS3j1lbhMY9cTQDkSngUwg+jiz3qli7PRfNjW28Tc5Kv4n6GIdrvNsTPveW++J7cLeh8
sVrZ0kjTMdF1Wh2FDft6P38/2KYVohAnSZLq0IOR7/8qMMJ1hPAvvBbJ00exFf3Xq+Bm/iHFptfy
n0sT61Y8nWteygEF4XqjG41ifX0zY2gzddedqEzCW2oOZNN4LeCGTeHs1kK0Jg4u+KAcavWCHQ1O
yrgWGFcEx30othL9MSO2E42ruFoN/RgZvJlDegdEXcpQ/isQ2s2OP2pbhtc9vvTXkaGQjHwhQlRT
ShyKMXkhjvYfXTxjQvmESD9OeLrL+r8R3E6qtYfYhHtvjdTxZaes/DSyD9TKdzYuDr1UCBoBBkIF
zN4IjTxo4nin2JSoWiSlBf8KZrNUmpzSt6n2+vR5msiK0lCOcvM8cKzZOuRBaRSJaBasP+HvEdcw
pG9iPqHKkBG9nRm8EgJIrdDarYx7izQHvx+BXK1Dqo5MEZDroyfar34pjsXilOHi3yQ9kW6y3gjx
fop9cZE6zAMiZW+QtIJBPw564CrXsr59pJoD7bJriAa0KibDxmGbxNefqOIvtmFjRWmRRJQsDdA6
TyFqoW0BpW/3EJwJCAhfvuQ9Lia0g9Rf/ywZepOOmF/2l9oXsvyOvDiVm3UlwhpnaL9bxHu3R4jy
OLewOd9NtNHOyhGO83XfR0EAEXaIHH7s7UCniRHIbdPZNyNnbNGrFsBM3J2C+bSdtXm4Z+PJ6/TT
lws1YQztlMFr4FrQG+CnelIuz82bcNunu/XIt3AU9y/OpP5OxB5BE8bJAxtu2RvE6hoepbyGvLop
3HgLSneqnAKc99prGmm8W2WRtY5iDzbAVj/KrhiPTw2Euf3qvH0Pm89RnxAuY4kBVir7F0g5r49Z
pSttrrnMZacB5Hx+3aTeOxBETiEGE5poQfYpb9a8026K/1Jg4gPhFSK4jlz9bT66cO0cYTdro2xI
T3Qc2+9svV7j/1nIKXFGhouzob6djGyO0VVmvq1IogXnEDXqBP7fDNayIY9+XoI3lOcwhj+u3pSI
Ekqvfpvx+poqWrgVvj/Mhrx56vxglMf+us9bPBtui8J1YoGESdfeT8QgDLy4varcF+kT/Ukb/2lY
mrhuJ1zps+gDp9lfBeHDKP0sAu5apBx/tapdM9Q6dEv+7HO3qrbjAeSJxUujaQ7qFfL4z38dHcVM
K/IccdZQbdFZ5NpLWipMk8APHZODIzbD9F7kONvL5yWVJNSvc0p34sK43r1yjF4ZSd211ouP5Ah4
PbHk+cXD71WpoPstQZsEHsYG2zs6F197pHpQHwTikJgcjjEPQxrMSY7/tnkkgRzGQKLLLde149hJ
/sBHYkq7ytbrXQLz3M5CQKtMHju+RRTdBFSmjZ5U85E0TJZ7996XJwr1X5y9y7OfXe6efANT8gtq
ixkUSoexhGyUAxtvIDWDXZ7gq7tEUDY0oeh9KiHrwNDuGJkpxvqs6qi4mqVN9i8DcNFpjhrfv1na
I9p71q/BnSmSmRqNDrXphip9EXLUpePW+k68A7Y9UwO6PexQVmam3d4bHxjUuxQuvqqHqi5jmMve
5mhv2hMWhK7CKL2rApEyl+B4LNwS/CK9pdBVEGYAwXR0E7uxTH7J6DV8jSuntaOlZKfO72Rikv59
3xmNRQUYCiHFel2nDrJtsvJglFhuiu4T04NlWkHm59aKbJuv/ozhKXqcTDY3kGgpQWk1tRBEXuiI
TiHBuBIQoXZbQQjapZ64d+5+y7bIXuD9m9i1e0zTSvmSsKNU0WRWbdNwnscLYDgsSaUUGV0LlGIl
fNKl3aQM35VEcB8sJ4ono95rimwcNTys1WuW/NYTpGwcwtQ50pb+myYVzfCkPya5QYQL3/CH8j/B
bUdxzR7cRmlY/zybY1UrfEB241q5tWnbajTHfK/Z+nGrtvQZA9V01b5AyvIXVYRkgusDIh3bpCru
NaejIQYfM4xfRNa/jhcwwYHGwW99y0hXRhPf0VH9KZeBHS96QqWX6FgQW25vO+03CD5Ab1Sgckrx
H6dvN1jVeWR/OIrK2K6joQAXgHT6aV3zUgy8/GhioI7WO6WSceJHupMz2Uyiuu8DGA7+rt9JLmmE
YNv+LbQxocp1994AbRqtTIxJyjLSqU3F7nlhpJCOE2eJRlJxX2dhY8uf/2DpxZPcG3sziKu/AzqQ
Fi4B0vEU0vDncJtvMc5potUxO0OHW7UTu7VyDxf97IULqtkpXIHwRvbGRq4T1R27RAo32OL24CbU
CmUh41myrXnLL+bsnJ40NYswG2ssDTcV9TtZQQIoHyWEv1SPWs+JuOnNt47k8yjJOo71pGFkqkE6
aFlvJSZoKyr4QCKbkZAbslm06m2nb5e/uXHPJ+lzYG8Xsr/zxdL9gOr1NgVc2rHUv1NEuqbUjpWr
jwAIJnagnCEW2rgXYSGX8Z9wpHNVdCf99Id8FSN0VJi9JGAod6SS244zaAPz62mS9fGop+m9m135
hwpz9tk9CxXJn6Yh+OkUuU25jlbVZSHNkHKTru96BJQha0YmdaTv6P2utiHFo457y4y+7ccIt7fD
kQyqn3qYG9Xeydju11T6wouuSbFi4r4F4iaD8Jx/t33YxZbQMeLx4xBAe6F9baQ0Lim1a/wdrrZO
qbFbRuzMQEAt7Rs0BwA3iUTU6msievMIYsPHAcXQzH6L4vJ2WF8l28tvYLcIOCb31p/sPpmN2efn
FeRb6U+ipbxvOjzNaFpgjRPPzQgJsqW2x09uKdOmdxu8wkw6L3J3uJd96Af6CSzkxPq8KEwz/xYF
9PMiueNrnvipyyuvdTzLj6ZON1ZqrdChvQ8SNVsXZw/RWarK4e8q0mTRA0EqlaLIijryUpBgblyD
Riw68sKi1rCpst7qOmxVsLEFUWAR4mxVFkANRaY0ieRJXJd8dHb+7OcjoAhrXsgozaswqvhM9e3p
NjJwcpgUCv6ce5aFoNlSnVuUqNjEHWJcSIy6A0Fbx1Ctd7eAV/wxaEJw7dmA1bjxBe7kCF1UCA1W
qvm+Ek2Ho7P2Ro2Q7NkcBSPkz6VuzgPQlQAq2q5i+DKd91PGLaHSaa2LdISkpplC+rZP3LPpWAvM
0r4PtrXt1IRlC1fYI8wKaZVoAmEyONIUP/L2/udAaRVyDHG1BhS3AlJ3mik6lneG06UsV9/0XEek
tkbHJBJ/Q/aiasPLhLDHJiFhBQSK3Kqm5Pe14Z7hg2qRa6+zvT72HWuZYwPTNvE+P5Gd5iwAwWOh
g9IaBZtzxiLVYDFrWGdFdVEcAXemkHfXpZhFg1nMssgf4WbN38E8XumV07my9IqPv5EWTYACmmve
Mh3qLYIFt0pDWGDmu/n4LFbM3LM9JLgAvItlN3ryUaR7pbpY6Zie1UKEhibwHhZI/M6OMs0XFFAp
XO11QMVxSmv1nhUUJ+g8viNXFf2/tvfY2OCiw568rhpTEiWEckCdxS8jc1tF1BnZwJdSXQ8mTtxl
5/pNUtNqr1PiEvj/vKlsf7rmLvtMDpjnvUxlyfAemoCZaVMnTLEoOPU+xPZdXpOZfbwV7kTWTzsI
zebuICxO9Q2lbCg2Zg4GKLfAKZWIsA4fbAusaAuW75bTzCMzHBlH4zuSSTc2StxDVSl7K++Z1XNY
N/LBoIr798aMsn6qnCBk2N8yo4lfGYxB1F8RwM8DPQqloIgUvG1bSXR06+dEVl7Vp0XIn2XQ7A3V
d51sdkeyIzzQHMIaMakRKfNy52nFIe+ju5xOrLwkrNsomQ8SUaUFAjoNMWuj+MxtbENF9lgNfx6F
o4EUptuqPhc49W0IRXsJ2wJ2FcBjxeoGtqLzGjYss4DbVMV69ruM5cbVyvGhgCel4cVvSX0z/QKP
d9EVIjxue4aDns/AOtJCb6+Cn45LGvlcbgiwIpjhY0hIZZU7i588NDcF4JDu2cCD4fsotfu2Co3w
xEES2NKQGfpegH/jL/yo+cLOLsoM4E5nLA+8voJqbxlJ1XoIxBJUTilXs/zJN8D/3K53FKT1XwNj
o9p39fRcdRa0GEj5se+oj7onFyAcy01esCg0j7GAEfEagOhSeUl++fFmOuWQWYGRkrB8mCcl5qm0
axo3CCwep82YAtldk+at4gyFRs3+uf9DGQXnDTyHUYDJjE6qMZ+Z2+yMEaqpD24/lG+S2WxYc/BM
ooCiFJLEFGNYhj9Ubm0SzNLh4yWVL1YTw6AvZQfk1HP+Xd2kq6TmYpmG3h43Z9xO4po8AAfV9wzT
GqNLOS4SA5aY8iUMadNY2m4y5WF9G3a8PscLc/6LyT75+uk6pBfPk91r82NRLEAoHP8gX2jROiDS
G6F8+ZH/12AGUWHav5WW2aeEHqFoJkQP81xpHxyMEuFPdSLqQ8qgw45EhHiHNcm/cijaPlm0/H3C
Se+6nfwOJ0DCdaKygJ7X6BDWUQtPr68SJf8hWjdugay8kReP9NM5+B3hBGibEZSKcHhuMcVLohVR
Dj/0vjQnlSAZbKAIr9LIVYZ6Ci6vW3ORDfSNR7bCeIMvaiDDlecqWpBovDpSqR3GSWODQMTxhD+p
6iiYTDQ0Y1KRGXDeaWBpJZ2viTLk3DKtcrFb2JQ79UHRSVu8f32tdvkuRq5zsZuemvGoWzUDPfnu
QgqCZw1sAwoUCVJ7NSufGV3AZtUZHL/07Pe1csjxouJDtgUmlcLOT+VQFB4zYyRmzSzIKJZcTDGb
jPtLQNkXVEKVsBkyas8/vMFQlVVER+QZonoAy957HG93Xkt82DFdQChReeiD2Kl8bXUvpPgVB73e
ysG+BWmjXFqcicMfpg+BAqHbr90YzzhfgZEqMPqJamE6rShJQTJCGnPHiXjC+ADHGWS9z5mhPa3q
r08JHp+jW5yWmY+AilhagRns1CfgvnyeLjEMIkH5qw8OWQVm0VpAMCRatHL5DeaTACqp87bRiXwT
tbqc3AG/2ahsyI1D+IudkFP3x6osmc/eN81IK4Efe1XipBTeyQ6oya5idKBGIN7N284t5PSvbKUz
CtMiGvyLP8pSm7Mrb1apJ6ehv0Pz118671gSTccLz1fTIVd+SvIad5bx1C3S/lOiKxQ1EGoz199Z
IKknUTeYu+YVZiN0xSXr+qzodLXo9KMeG96t7180rjsDPHX5c8Fe+viLFjhD1ySr3KtJfch+Q48x
9GPI0C+JOcPQVV+yTU6G995F0a3eqPbgf7zEIIpHgdL+znPG1z0Ufn9uFjuuehBwV+NPfE55O7az
V2BSkZ+VIIILzWjPy5ink1Li4VVKeKa1T5yZSSw9eiK8J/yBXjxOp2MjiHRJd1qDranuI7S68ywY
ABvhGtZMI6voO+chw82d5VW8Wn1bc6qc+yGRFirKNi8XWZy+mJYI7Ix0aDyZw7aQf3auGRPXNMoA
5Q/EZtbNB1y3s4gzGFzQdhn+vIxfMs68sIrmTicI9rOxP7pCRonziw68wDg+HoJ+odW/wDbgPrAl
xmmt1lcQFMlE5sI0gBrKDoecpGidxO+NtVND6tGCCna6VwI5N8Nl6A6KvY6M751+6qFuEkz9n4Zp
lI2ooZaKRJ3p/e0IxdtiyK1nKGgTggN0CYFbm4OpmUAOlznfdBrr8d0ggleoJLKaiEUNONrXe+cq
3Q8rtphJKACn53zO9tsJZ57873hKVUVLHxH3K09gMpOrIr6QuAK2zWRpD2KBnOQyic3xAUb4Mf3Z
CeOogfy/7LBX2YlzGNuxPYkTgW5sGTY1nKLlNLBkZ+FJOQmQZ+egvME9ZKLCiZNup6bYjdHgi5sW
j2X5NSvo8Q0tAPFcsx+8Do0VKFR0R20u0imz2uP773YEf4AYgcCyzCrybU15IwiZ67Pe3aTaudDo
5ALdvzJAczwUjndNPyhCtca3JqD6rVnKEVFNsZx1pEJDI2CI5vx0/l94jrF1fXiSLyiVtd1cqLpg
Z5JpwxCZKr60nNST8ak1mBIM23H4UaePi7idaiF8ChQMzMkUITDgU7p3w43lmbr0XJ7M4UTjSFyF
O+ItZuyKj7PDz6/GoSnYF1+oBI/Zfhwinuo8jmuBSvLXpMNZXAMVTywgiVbx9QfOR/NSZJ6OOsh9
FGt0dfK+s4rZXtjHi22k+GPtDubz923qbfuZYPKMLusY26akALC2KIB6tfd21LZj8lQjckIyd85V
QpQX+nrba2m3RAnOGWPvvb/gM5Gic9Lv4CqUtelRwZEs8RnBzlgYzdJVeLiJMcT9jfeI0X9fV6Qq
dIrtYYNxV80b1pE1lFkLhTkEJWOPd5sSUj6FCn30PNLKN5zKCmosV5Dw3O/AazD1GEjVHK0hziZ/
KKdz48HnehUaLgMciMwZNTmrsGIfHJGRPibFwK3jKT6xkHmDrAHf5kFZyVBHxzM9K0pyHF7xco0k
zgAv6ehNh2sfL35Yo9KAeOD/F75Im+oDqcRaSmwa473UgSCgAIGmagUs4eaQ/J308mm5RQ6B3uOR
SugEOfjGHfbgprmp/iVj5x0BgAUQ+EIBQjlcJBZUDGa/rbaOu50doBIyU+g1wAmN0ElbwL2SRpS0
S6whBdI9m3Zjjwso3dD3OhT4xqlO/LhkqXz4g75FJHZC6TOImgMC/sZ5byUfKE9+wV4q3ACU6sIP
hSccGPCVXTr8pMIYZ05SvyQpc0M6Tui7u1DCvK8I3M0kehkrWVde77QPEG4tiARi51VRF/xFnMun
DSMOEk2rYGFp9IkirVoKtNnuAIbtoa8/HNcK2lG5WAurJGzxmxu1+PZ6pe+x+i0gtl+p1FZwuM2o
i+3bJCBZTkhAWHbKNaiOF1rqSITH7hCfki7N2CLmpngsMbvL+qwhGQ3HtoQbrxm714moKDo0IlyZ
0F5oa0X81aWjisW+RVY1qPkwF9EtqF4YH17qxjT6bIx5F6yznAijtpLP9jBEgt6eAQ1BVQBZ2Q+y
ACJbrWqR/righjugvtGDj10v1ZLiDF4/hIa6+6ycF7T9X5Q7PLPE2VKZWu8L4UTn0e9mbm45jtAU
sSAhAJOpMnIICSxl+NVj84PcG3StU6EwbEo/4BGEtLSEIR6r4RipfadghIFwn6JevDFEB5XF0aVP
j8kB1Se0mR9tHjvQZETPvFV6s1JbT5QhFFT2Uqgf6aabsZ2kOWUY9WXdS/4Gcu+alAFL91RH2M7q
DxiPn3N7cyGy/yFdhakXV05E6c9sGj8flYKVElMoGOiMfOvmdPxl1Z132waErg3JSbfQMU5pjU5V
J3TgZmDs2qM7heNK3v1q/9kokVOlIc7qj/snPATwCKhiKG+ZjCYi9n7gyxn+XrS4/YRzTTAv5DWf
oddXCqzOtXXduVqWmbzWNedgyy5wFBMqdfvW6sSgp0mjWkOnA1QZja7Xyad1YOiTKOvJW8Iv/iEb
Toad5YXpPtFqYQc/zVYjBif0yxOtOFaOn0GeGsdzkgqVhf0VfQf0+NqAkAqrsvzqDptCgNipFR9w
9jWqpzjysapyKSnWZtnOg2M9dZVn50j0CMd86xl/4uzWpYEzWcqlm0IwqCJWBn5Xhtd+3i1v6xsc
NBVYMkpFnF5DO65fHojmQ+knQ6ARhJ6+qdKMGltPKP5COmIgOY66FKCJr658PhXuJto+ZDy+2GGH
N/27A259Ihi7qnkxTAvjP4G0PXJmrHEtplJj34Y6/fqyKSnScAhBXsje2MBDgbSopaVhalHFF5lE
HOqvTz6BLyBtGiuDGcE96Z2crg64IxYb+nuYiCLnQBNEAZJKAEGu1lilMQqId/3z0y2Lvo3FmSYX
vMwGspgmbD6wYfICe5hNcdg02BTefRdgdf+TiDBnmJyJw+jX0f+hGPc1FryJoeshFsrTueQGr2PT
DUzatn6Jg6/oWBHGJ8jg+jDXfx2ku+IsR5CLjCQkFBJ48UtnpWvXwWKQB75uXOcczP8CdHJvJMEi
ToTKW/aXuxQmQ62B8YCxiuYF2Jd4EfnFWmgsJvBgwET7bogztVZr3GLQXGpy8oFlRa/Fe2W5r/jQ
2KEXygPI02dYNBRN2vjdFXsewHDvq0AiGTMXUsTrarls/JIb842+KzIa/a5M66V43PvY/V4Qa23O
FjgpmXEOLnkRln91rxXVk8e6xyLUTbikTdLIkYTHAI2HkBrfNbverJujX+aTMNNGEE+v5SJEd+G5
/bX1WJJZi40i7odRGZcW10RYAXv4RrjPN3DhsnWxtEPxJsKtxo+hP6ZN0W4fcDwfu4/91n8puRwo
HMjcXmJD+0MP61I2YN051j4RRrCdE/n7NHoA8QrzzFoSd4KOw+WLKsWWct+blDa8DBENoFZXSGGK
BtxMlFXn6NdKPK3/OmbPNegSVdRPk5n6txbrjlutRhgkVwB564ACNBTtMyFvJ/4m68+0XtMG6gm2
5BAXplBJr5HzaOmh8CxSjdfb1tkGmDWSIENhtZ+1chrta4szQj2VMopqWwp7+tQMlQluNn/Twc6+
6rQOKZF1h++KqtKGtkbei4/hS8GGAH3Ik/a84mugPTaSH9IqDrEvSAgk9gktBvME9CyCC5AgmOVz
elZcHdNZgs5WeXHJNATLInEfCri4T6+QqP098IlyZqxBK0/EaIntvcBbTNlnKj8buGrokZoZ3lSW
qvRRUlxiaI0V6RtjqxP9m3GJdFLK7GFYhj8sOu3FfUYvgpcOn8SolP4hbg/a/yEA/fy0IA1T7SsX
LEffLnBvQLDIQe5Cpbn72AWoJUce8Wh1+ZOM3XB44iVIJkKzn3Xpk9SdMDaGjh85eTay13gn4feC
4LWku+srrFaXYzUwnrIIN9k7Ek6+u4eysEyg6HB5v7psqLPqGrWVUN/wG4CZQ/CNKcvNB/zuGtcH
RCvDUQA3IMtglUjhbLwvHhBpKgAAplboIOf/S+2yZ5J+LSL1+QOEe3QIbPkEBVUPYc19u9k1SgFf
dVPuk92nYiBH1oXWKLdIS8nSDnnBN7JSzj1uBekyJKYgSnYHiySJMDms1H58eMb7tF0PFOG6I4vt
iIrkdREreft25tUFTAEo7H7FpvvUnfHBX5P4c4fFFCwV5/pbb2QHg0+rbbSTpLwFCPfUZwIgiOAz
pG6eTPmivnrGoJWbuV9pQdtLoIChETrlihw80oDl8zG2bM5NFcbtavSeA/S3M8HtJ2kYykSF+tq9
MxUsoF8BEyjUgCpx8cytNSWxyuovGj1UEXBzVHzmsWSg5gXIxmwQWuzDIPlVKh9oRQz+L6t3iYxF
bBLN0dG+OF6tlF5GlOc4AXx7FDCHpFCk4FGztqJWmMQMjWHVMksItw/K5Hr9Qy9MCHwE4THOWt4B
e2Fkcoz9crK0CN8JnwL+HnahRObJOGb2tl75SQ+sIn6HiusVUI1+I5XhQTGyC4ImuMzrIF5qj0pH
BQK1glmYOgM5GO7RmqXZjA+d4JkZGRTYnDZ+VIyxyjMoxID1JSxgLJV3D/NRwviIUu3W+1+UC/JP
dRcz+vGR/06KMmPVU6/M7B2S7SW4OHcBlxBsS3Z13p5hWmgA4rEDdQj/MFYls+lTKVTVe3LB3ioX
66CDG52d2Y8h08TB+3HucyFBZmv70XMvdAE/7G9PA1oakTQlXaHae4YDTarL+01R9okprKbKtxkY
uVLU3D7xjGPU3vqP9wNIbIVtMWFqHi84do4x7p7iMmn9eKXTv7blW7d/IJhX8vJAg1TggN83ZGAZ
qoOEY4GnTi2QEliKKfJNe5yn4M/xNttDTJne9Dxv1ggXjQ9c3bUlvJEuG9Kg97tUnfNIYR0ILpH3
NRMUx6vfx0nyURILF5WFSmVlpkhve9etoCLed+JFaoY0xXprI3eF/Ggbavu4DJGmLGNjSTPdKb/y
WGeoAZVa+3Tj0ejVtjX+D0tJoV8sOADuDTPth0qIxQsXGO4PzE7m48m+b7l6AZTdzUIPcqubF2Dk
jP1btlhNBBDbhLqOeUUL8xMm81CKTRo83W1MiTRDwJHBvRjOCcwEZfkhqBzLa0+3CstCh3wSE3DO
WfDezbfII5ndEX9p1SIiFpGml2iw0UaErciL+vzhqX/63z8989pplhjWDqcMC/IbLu7V5N+eNWU5
XAbo1th7Cs5F6/sckVozgqHzaGoh3uHRDP9zD1UV7z3dKZgD/rO0mfXgmeY0sch2QCN+MzNbIA4s
Ecxubi8ZI4VFHPOFOuKmOlrLsI+YdjdC67PWSipKqhJv0ckleLHSUHfbssCNnMJK9jucbyiIl72w
yscKalqz6LPXr9hbAnpiv1C0sd078Hy509N9bpCJ423Lr/pb8Wv9Fx8qj11AJh/6XspNJd2e33GH
LbeMcb6rC/QebtauBfy93LCAjcbyx8QgrCwowcHfV38p97mZ8zelZjowLbXF7mqzgzAEFgKSPBS4
Gx4nO/C2CNoGoDuz0yxnJMep0ns0AnKHQLuN6T6b9A75czUUGkPX9Jo8pmUjp2BoB8jsJNV5lybR
hB5mfuDN4LwZ7eZk0UoI28Jwfa0G7eoORgYEx8qZAsh4qhqWRHhdPOZ/BJDwmB6pB53wtTk3/eXy
CauaVk2nho9JoVti4M1Fwttm4w3tLl0f3/Yzib6DbE4QhO02ID49XLhJkkJXeQo1chCEffnGJ2Za
rsqadlIEbjocsTe03QC9OlAdiHRcwFozlVPyBa3cF6ZUipd9Re40W5+Mi5b49OoFEymm2L/Wij/b
/ioty4IOL4Y+IUaky4b5OKtx9oeazk5uZID3Vq/BpX7kRA0x0VuihsmQpq3oRqcnDZoVrvWqB9Bm
LCkqy07Z7Yao8fN76uiXHf5JoOcG5H+xbZMuUEFISqdpwmQ0YiTzDYnI8cyF0eRWP1Tk79NOtH8n
K6HHgnJ1rjl4+vhAGRQ3j2WVhjD8uhrkLPh/mZkGoXrmU0eHZ1qOcd4Zp4FlagheBXGc/abV764v
lqyl2AQUcI8ZPbvhe4Bsv+8NeBoDdOt+IMa8BaYAS2ZLzHSJqC3RP3+BNAafWsVqJeBoFx5Z9vB9
fXH2uMOmcnGaSAnpCH+tvQCBvat5skPMl/5Ou9UiDm0L7bDhQle/lx1ZsUHDPlqdtnXjvMwkLqv1
eyb0WKOdCDtCWew+BSwcJUp4PrI+Ou0ahY1mauoZGlYdfXdRs8aKhgy6W2XS+bK/isA96sIg+Xsb
jAazhKvj5Kqr17v6Q59vM/ZYiVuWzYgg0GJpNCKgSMcVI/hMHJSzFPvk0TKplLh7rcItRW1nevSa
Nl3xFTXe5fhWhLT3eP9bydTzUkG2WECdyeNJZTjEuSJsxmp2Fo8vYDM9yNks3pPCbYxxQocKDdfO
lmprz8ur8BREqL7/k7WsVwM/FGmRsEcUXTJFU2EuSkUT4a9TgDFn434orgtL50DBDrkIYzt0rGGg
CAXPQTst6F+5d4q/UWBMKZqWSF4VLbYHAYWG6LaJBtDilKCiVezh1tXDo5ZWo4DNb0nL3GlpMYvF
WU8j8rA3RsOO6XjifcJBuyb4YRJnbLspnSFNAKGFVTp3kB6I4Y7PHWGSRhnLNJv1U2uw7mYbciyU
qEAV2GEVKB3SX4IBtEurRlaNB1YRsF/BddLTDQYuMgrhzEuBUjz2lB/CcEI9Fto0fhLGrvbNAalb
cV2i2MkFHLmXeOkxY8/LcqdIgdoDaL/zboNX8Bt7keLYfb/WmScGDp0rps6G5ca0OButUlmFVkXb
qHFz12zkZsaaU6nXAEG/jOANym4Dq7parXj6SUksteQphtp/U5pSDGkIVDGyZuPOT17KZKoG3uef
/OY7EdC7Yhf1LezdK4hGpPoMRP6UKzgr6c19ex9WCPg8ESkDn5FUjYIlcgRVpNSzSoyfItP/King
mE1+NTZJMqqkugrnLWG15aD+qK/7tIpXq8X4OVbk7bdaRfbY8vnzortmBAodUAWo3bukxZtVAhpU
pF5cdQpQDhA+jS8BaKS36dE/lF9PR7dUJC/vViKdI8QVLorlO1PgTcfkLM4WuDPdYSw7KCR3xBb4
HuIywTMdMYfhwHHmdyFa4cJBFS9CoWhTS2WpvRegS+Z/o6y26+kzuVoptZScjNL9ike2F+hVuE5W
CxlfpKNvNfR5+sVDT/ZYNjnldk6IrdvqJTb1tNp8JAedpMO4ux96nkkF+n1Up0AmmjShk7DjyXl5
ox81F9+1pf3YmvRiwSXbTD9AMNXHr6N5FTp6K/WEFFtqIr0HDh6omFbVJdEmwK+ZDQCNlQ+kqapz
CPH19guEH7Vj2knxQ6IbUjiiYkzP1QL6GgrQ90cCsY5uD4hFF8DHuZwvOyuVvaM+5kC4MH4G0+Ak
KurMEfZUf+SpeRq1CSlL7/bxffnZzkLUSakZgOc+ezRc90PtPGLvuZFwOudDS08k/vZwwHLdF0KB
semAImferEqLJzsZt1eP6atQtsJCuad/s5+Jpt+EXS4dn6Bm4OcHmRGF2HJr1NCVlckXI2xv8Vg3
978/Sn3luPwYN9Rgc0bSMDQYXXxKcXCQ3EdjHySRS4LgmbCTy+9lAZo/yuYp9sTwOWkJgX4Tp3cH
sD7u8l2US8Pq9MYTuCPfDv9gKUkBtDaQgXxVOQYk5rb6me30Zf7POulNmsrLl+qXOwoJSnEQxsi6
WvfojncDTzXSYpAT5llwAJ35WMrkPKTjG6VMBPQwJUjkBpwi4ufKtt6odPT00ovAiJg70jgBBtZ3
75GnUt0PjATS43cy7n4KdKFcJkKsbCo6oDkZx7pAkcfx69ib+vVU4HIUWBhQe/oy8LeEQAURt8r0
+wkXhm3eG6Jq0zMN8Ku2IZ3UeP/Zzit+AHoGJ9VpNVe09GOq55qCFL4vI7pjCUN5qmo2FwYq+cSB
+SrtWCGRsRTq8kHO8vFJvSoBJuFFHvKEDb8UDvpnwqYRKqQs45O6Wtx+OL/zeuwS4LlTLuK11B5y
Bt3KrlzYAvUn+VVXEXe6/7Qv+jiWMueVxR2/enijNNQnci0XCzFKEB9EoiJIdnT4YT6CL0nSgfsI
FzXXOKGIrkurSFsjRJtiZOCvk43yRyZz0MfCBXGAInaYv1839HLlJsuOfMdMFJJ6VSZTnI/CrQ+z
+3tUF0PrgZ4Xhj8KQyWDxej4UPH8jSsJ9Go6eRYJ3tyBJgenGfEXdN1Pz/MMTfK9TjRfufBYnay9
pfNPePLO+J2nLHvhxqNrABaHPOKVmSkCb8ITX0apeUwOJkaduT6732YonknyZPU3xfxoHgZQKQB8
2VInQlWfO0IAO+g4JO5NrTQGJ6jRkjJVS3jM9sSmiMmx1/dlUdGpRlCGallpGHr+EyYZ42zbmrF3
OAF/SxQxvKRhpbPEGdrFzwlEsjcoNi8epVrswRtwhjC95S/C/tu0Wz4+ijHg7ZBxMD3v8VeGYOAU
U0cmmJW8u/x4TAXryZKV8HSolhKlXM51alrYb5Ys7WaI9yTSqrsU4p5SaQ1TxU2YXEMClWDFWL5e
+s/Zn2R2+j0WSgheXJ96sEz8/gwmZcB/A8sVY4UgIHAe4q9caBlLXirq267EYD5dt9O3PFvjxcFK
iQ4/MwzeMCGGxY0VQIN0MD6Ws50pxQKfpTR3DRfhloAs0jaOqZzpchuQWpEZfztUeHEarIuZ3dnp
RLc6C5T8aslO9TkwUIymu3IryFF9miF5IfP6EyZGYhFXh+21qSvEAUZf2qULCZ20eqKmuQ0kZuXf
JQNpBEghLUiwUg7b7b1cP148y0nOZ3CabusUoAbPiLmtObjf6nXgYO0evRUbn/B0SuzjoVrBf8WM
pwjw1Yi/Zh72BlpJNX57gepPgmbgGI3hjLdEqonHog/WQ3W1ZmHZwriU8wWj0SiECvfQyexh/USh
lMuwj/BmqpIp9LF/qoRMi5YzqBDhyXN/uPWeeilPY1K4cm7o5RC+H1l6F86b5WS2VFJR1yriIwLs
2Red7ibWsGVLrxhzKVlQ8caHZSGEpmUpBO/tbOHE9dS2BAjzavUT8xRe6sxPex6530bXw/1x4hlI
DoxyxfxAGVeuRxQjyAj9MChty+/ohZGVGP/z/Oo5PCOKdFccXI/nvmvGxmof00s+Ppz5IhfqsWw1
Svjix4ApaojGq+cHVkl6zi0+aujRi5wSy2qiMmuIqL2TPPxOqz+vIZYJ1r306K1pA5rV3iadM/kD
uOrUKqo5fhEmZmziEA3P1t55b9QxnEA1tyEB2NtPB1/xg9Q2niE76A8mf+8DJpbDS7+NDwi092YV
A317+/b+Jm4AHc1g8hScHJ8PIBOBXCp5H/wkRf3BRLLmGRFMELsQ/QMC0yJOZk8tMJITw4rswvbP
JzNy8XgS2k5kTxnPGEyrMmumavwIoIBibn8A7pB+wTU9xzzuCeTG5Q9BDx1yyRQsFGtM56jm0zav
agkpNd68HV6wsDcaG6D3YWBU/BBhxpfYrqjdEzpognh/IkGNXUqtiEO6HVFprh+/teBeOWUxcS6m
BUVHu5Trqratj11Ja7RS3YTilgV8nsame8RIUVEzAEP6SZG/RUnByqJG0kblP6kg39mWp8WdLj75
xbG14Ej21lfwxePWzXTKv7/I3u6hflxvnq1q5juy6expwLgf7zh5KpZuxUSH5hNRHpLT6cT1kkW9
lWpQuLUt7wdGnxAmzsIs5wuLbwE0ph+t9IaCOWEasx1jXUFFuMij4QJ6k0CM6BVPDQaYUz3V14VL
PWAWAQUcAeGJOu3KMwtUswh3sP0JSNZ0T5UFu6v6OawdXmxTjEUQLDqTJq305asqzM2sufjl5vDP
vu+zPeQESk3pw3XL+z/+G/EnBfJMF43eGO89J2vOUFFmPWf281wdYgl97BOypGvvyLUrFVWf0dvx
XzvYWz/jhtregbMB7mtZkc/P+GDrPBCqD22hsJ/VOOfbashkpSA7wrbQOZ1QMbTvWXQACYTTtdp/
5P98D4qNaQozljSSCFiU+bTtigzoQQTSpZ8MIVRpLLzKtZIN2IdJcGPTnRUjetlkO4A6AyHrXojj
1QTOcuHKXzRUDG3gmI/uipknlrCzJKEzvoo480MKd+ChnNqdnJsVTEx6+jRsrK3/Aibfe2eRfZoM
2scPjZhy0h/0QjRCqSFGqQ/UPcusNDAc/8adkayJFAGqhGoiChPervqmudtWM+CSI5oBk8gYjgZj
+GYrWdxAXrk20509+r6VSKCr+Gwz3A+0meI4sXItJbc64BP6SEuZPxOWnpIrmLqmBPDR8oJMsQSQ
+Q15Fmkby8bsDbBjghmIAJthIKGQo8Z+W42H54g6n8C5NZsZDs65SezeaCsFFAY4r7CK/vLMFMVm
LT5I2RmpDSKr5oikGKa7FGjW1M9c+qRjbwVIYMKvxVkpuGBPvNXMHzwxvHj79QZksvSVgH9/jKRt
J7c/67dzGLpONOp+BDgzAd22DkmtvnVguGX9AcDhmEDT5Ioo2NiXXIEh6cnzr/xH135Khk7Qh3aH
1HZmg5DTrk3NkiQLtu/iolcYOlG+VRJ9qekynr/3ALvxBbyxyq0sRcMYKulTMSXT8EIT9mIr9bGq
CNUrDU39SOEWH31QC2UattIzM2zL1T2/VRkzFVsx3tXmr4+H3zYqusdA+lyUw0to4+UAA4P9oca1
PMB9ozxLK76f6qVF6cknMYHsSjh3VFX/FU+bpxD/nSYkHxnUL2Si+9cr7DLipoz9pc+NLLFH2pwh
eOyOE1pL+3OVGS8lsXXe5vbAipA7WDshROA0jwlQbGoi5TCu7r0Yw8tmmFvlT5xWXfrv5+dNdwQR
LP3oQ9l6WShcAC6LGtosFwPs7RGlUMXx7/OwvecwHcEgoRgGy2d7cKCYRWmKtwv3K2fTXBmWsoTS
/kYdAMRmiAKT3F2sIO7uKtThKfIQgwnxCg11uzlj7khA61tkljiOWBnr9vrBHZWWAHs6zIJx/RUp
m76XxvVax5eZ80OJH+2kuJxWD9yqoQ3rw2NTPU+yOo04t9slU9lL2YfKrpcyM0y4wDSmI1d/Uj7Y
gpYdYdQvoScFeLCi91peRZf4wEaeQUaCT7CuchEZ/vY8MNFS8SXx37PojZkQDq2zOdGYGf7f+TxX
kFzN5fwo2QucS2UbDdEabeWEUqml2sN8YhQwdZmcg9ALgiM3STFrnMtu9SKaRDIDAnOhF1ii6EvN
kRWYie0VGPf0kPvP0+SpV5NHh6NibwxCBNx0jyzn77K4Kigg8rCXI8yuxTnpOEV1VUn6IX9UM3Zk
tPFtvZgmRfZDymW1Umv6TYnaKDMMYhRdzXtVEcOS83e8NNLkSXPZNSpygvaro8CBAoXYnvSE0xGZ
1dbW8QIpolkGIavCxjaU1DdUB8jFnFjiJvSHbhgtspAknTYdkmX211CZrpLabIIgsOtz8BgCZGQT
fdEnwIfHYSUeU5tE8UKUImCCb4rrJGh0lqHuUFSrPdQvivB67hQxcNySC3YZ79vYuCwaM/FuM9L7
B4VTbalIe2+8euUqQBOloyY//iSBg8Bf134DsDjpnHIlQf5FhBBsT/qMjTpaZAcQpzuqHQzQGkOW
C3GXnQaQW7W4H6nWPmXth8N8kGukSXjuKSOkSRDg50pBN2QyLgPgCmzjvV4cL76eyi+nmn0t/VJg
1Y7suOtjyYA0wNTPgaPW4rADwcui+0MTudF+Fy0pOosvnirD4FmJJ+SrNhzvimsOviQWwAlZpgiz
+sCiIVV2syry0Axvqzt0QOeiHQuCJah7a5OU0C0JEZogoi4RdewJzowbImlUwir02vfX/8cGewH6
xXSHcUhkYiSlDs0QlsU720gZwZeqyy5Cm1z1LP8rzfRrOlaHqJHz+JPmHXqWacQWrPeUgRVpxk2n
DHI6fUnqJBDuUdDowZbfBjJc8htAqibweqMkaCBfpRIBVDdVyNzvRR7nI1x6aFSa+pV3CHBfAWvx
/QlSoVuBlu3b6O8dsiYhplvNwHD5APUhW/gpOHUilk2QXdurx8Uv3x9McMDZrenyv2sOWPPSM0cS
i/j0EaZEp7nC1yIPeaieaN3VoFAK8bbDH4tNrWFnmbrgfJ42UdbUMMu5bAqd4rG2pvZDtZOJLs//
ZkXzrAYE2B7VBjlgg0/WEiSgMBIx7L9d4nu6ih5PLPHnhiOIf+1fCg1Yd7JVY0Tpq8u659kU/SRl
6Nkt6yVLL3UzGxYNCn+grLSSTaxe6S5K9xXoFRfkBQpAWDdeV8Qv4wXRRJOc0rgCQCveI6dT6T2y
fF7stoJ1XQm3n+Z23xSSTD2w2VQUDDFdqvPPd6NX8/hi6O4FTEHXL+VB69Q3z+7r3dJA9nnIz7yg
rR4wR5R6VdnQKtoVQbQmqKlWiwC/hwagDgYDhtM9SlmmJjFQrqiyypQJW0/oq/jTubDaQVfe5Buy
MST3JP0nNZ2GcH+ODdnC6SopWfK/Ex0GY71ssV4Bfzgo6U+HOL2OMLpRjC+8aILHQfj15JBiKCN3
7yqQN7n3szsq3CSUBExgQAMfarl/fB6q1L/7adoKsLEpeqWPQr2z9G3ub91TbrJdB8K37EfSjgJc
CQU/q258bJEkvU8QIdnm20KFPezG1blU2Zum6Vw1NBGWmskELn6NUgSkkNuR5Av4erqSA2fwbZAf
p/KZkVEIg3Ueoel/FPKcYmgJs/kCxw40f3g/PuJwV6fa/hqpyNAdyRqlX1ZEJV4XNg9GnSRODcYQ
mdHQ6wrzGt3Myyj5aIHhI2zainrZ9MCQZbxestF7HHglLgczGZZn3pwOmfdNcFWDj4IbY3deFZ7/
z3FPMjcCTN8GYX5Px97YVHw/9HsvhvwxjMU46Ed7w9my8x8w/trcCd6Ah3qNtnMAeDmb1GuLYwnI
Pef6nWJxBtckrcgEBocyFjr88hMYI7Ergn5nHRUyHzrMAE4fyPjmqkp86EPFNh/DPJAf7Kx8vURp
Qr5cLdp2+rM02A8R0JSSHe1HpAjbdscZ+fMXjbkKbkMASjMUVxYQPRTWs1CifNQfdYjz1y8thNYX
XDVZPWxyNvemIRMTWUq311k5IY1B8Ni3FuFrJyo+DfqCqwAxjbpwApwY0uqzDR3uElS8EYUjDRCp
TzgqhABUpopsNC3a9DXnM9HNx8qpEOJ3SGKVTmV0hDkalMr3nies7s8isDgRzdr37ptLbjmkpoON
plQqR1x6+cEgVUzvCCMiYGyfafbuHqhSXtr8+/bND7a8JAkUIcd4Y5tfYpmyEUk6aKdiY9m8WL45
z02ryCQBbqQafK/NDWwFopn1UnPgfIAXId8vh6UG4woiE03v9ab9ovyY0HiUZfQYoi4nGpgwX1qG
mUA4aBZpv5KK6QPtiDGv7zohgVORHcmcBtrVwy115bIQ3AmmlSvTack+dH18u8yfQzANp1sIEdEV
O4VzqdBciasQr5ZxunVC6hHPG57Cc3NEBmMZ5aHRu4ng6llQZXWuQ5DhoKW3SppH4z+npe91F8ZB
RfYvFBIZt0iw8ppIh47puXAIBHr9QolIBXL8FKzkJMG1/LzLUH0IsNF45qbQjiBMzjk45v+ojzYj
6wpy1DG2sJ4slA917yb7bBfw1IGDTBi1GCK6QOmseN6/Frm5GxMQEgnLIvx4pmasZqdACbwC9kmk
nrOk09k9432YZg764kNB1LscBBFCrW9C1X3u6FHdBOfeXC2CJXwvZOCueDmaScH081M7ICUWWsDm
9f6O9KemRXJibOqQP10+f4KyDl2Ryq5s+aGvlL6JC0+jDWyALl6tMTRHWsL33cfTwD/q6ocLhs8A
c50EqVqS4ynmwNMiC0udCuNYZZiXycpgqYVrAANPAUDrO1M5Nu1ZTTcrJN3MlAjCQKHbEjdmUnAs
rFhkQ/g7iseg2BMBrS/PEEF4GfmrxZPfnGYcg17hLWv978T59ulbh04ySk50n6/2igkoRn6gw2nh
HFmigvP2UNnnLnX48q5fgY3Ejbg6SVGqYEO5zQVb+Ba2HlkxAbRZBGUlZhlQWZNf75JKxAW9HcHU
TJmjrA6qHmY62JpX2Fkkkk2QAJ898dtw9CgFzsymfCQWsSNnhk6ns00MQ3M6AV+eSbnDOUkauzhO
sOHSLIPkWVg9I7Xx+WbUxWfKG72ZpL7YW7iOgQNzgYXksN1eqZe6AMT95SvTCnPCkShw0av+tVk6
vnat/mJka0HkooOpFbllHrIBLqZVK4JFUcVhJkbHBJ9jO8WG2823I8YxpyY1wlVHK0NNEqq0dKVQ
ZKunW4pAUzRwiFcqZf7itDFj3PgVWJpHejHTbuwNnNn2FnJSRKT5CzkPNiUuBroH5rLHxSSbHE9G
aCbrkH4/fmy5gWSQ3kH3fAs5chiPWmRS+tbI6Yv4OeFdYGYVC1flF1tIph2FMUYzVH26BVA2jdDw
JeEUdco0lGi18FLGU/Pwbe2PP3Yk+IwejIlxntvCzohyR5hukm2FR27tQO7vMYfs/koL4qGZYg42
VqcPZXm4vXQbqBd3fWTTGsccKZEPCAAr9H4fPICtU5oaVKHX4M7EMawm11etb26nCWR+lMVc5K7i
FfEEvLJ0U5slt+qQL/ZrgdyeqL0r6DyolyPAexT/lOepWuI5uU5bTjpxeP7pLPvPzidGTN5loood
gJ7m15XqGY5XEQW+tJUB1uZiEztaO02Wa1p64s4WvYuC8+at8yqa8244/OYd38VoaUFi2mFV2YMQ
MUZe8fOwiuevGnZdPrf9w2zlo1KQ5aENqjiND2ITFTF/gkFwGD5tqjctypuiy5iBh0eZZZoePSdF
iy6JAmn210HnlExtAC8MOf0RFwJk8mB2ABLlLVBzLO7X/m8z8k/0HM0xmn8dA5esHtiAQ3PrudF8
VlrUK6ClG26WKgAKB/hxaHYlSrmYswGP4zKNMchKBuWDnC2zpCdq2VmUqXBqx4rzJvVZtM2wGvF+
7zMB/qsSu1fM0hUYR+NYdDoArIOhVBEgbyPf+4/dLUTc5Ia7E+VzWF21GUF9d5N9Zr2BKC7+rpna
CwolxDPXw2EswoNy0dxLvSnBK5a9DZ8Jx7OPstvuE2P+i3hsdsUu6qDXMMKS4TC+5cEsMIr/bqYg
Y3c3KLUb+ka0kDdr3gE3sWGCXhPAif4rPXWGBYRodE7QxA6NzCYpWH51LLNPcYByM0yDCBwiSQfq
pVhhCEw1TSjLlpkRtMXS6aIk7PyjPBrqVtfZNMHgl2PQyyp14xkvVa2zV2sLtl5viFCgxTxVa5ib
WJ2OCT1hiHdgmV/Y7SRiqkSsEKgHQG7bo9eLVMO3jAd5ps7YZ/+UMGcHsxREwYUcZsF5hHpqnk5+
nVvnfiAPD2x3CezwgoPWDnm99o8nDOyNFUQ0iTl6Do3PFL3ymUYOhIph4XdMUib3e3u2meFdKo0n
SA0Ls68ct+W4BOj1X1mAO3AN9dGxMFH88P0Ed2xCJ4T3oBUMLzD+QdixOQK/bh3hO/tZ09BSM2+7
LPOTmqvzhuvhH4kyuk1hnq8/FESD4Uh7ky/Zi21R6LPYVIrK/4K8Pqzz3SThpn66oKyGSXul+EcE
aTvqXsT5lImADKDzxpDdxHWptfOfKUmF/zfpw85JoPl+Y5Ivd/euoOIscV5xY1ssJ9l0HsRJ+9Sr
3G2aS7m9NgRd0cHT+tGyzquF9AEvxGdcHyNWwQx8Y4NbWF/ngev+WcKa0L3lX0IFkI0tya/gNsXm
NM+15DGrOm6yMri8b8naz1vGT+ZDYyd6Cui+giIgqdZ1X1IYUH0Hqwr6kFWiPtxa8onJD+DwUbj/
sluUiG31SvMu2gb9Jak6Lx4CbK5eJ3GY2mdkQnS4+68psvE63qd7qZGAwBaWBbMd4VV1f3TNGNs7
sdt9cOJYgFnBkCEh+MDeo5d2ZgwQrw8uDiQymEFCvnrCfZJno4xqh3I6zbzhRBA6ctedaOve9B4x
ZKq9qldhPW5kmkDTooD0jqYz9zhhNIgDV8JRrnr3gCVKTGSWv3ac47bYsaq9U94VWTO5EoBx4//e
x382hG6p65IVP3eV5u894pDm676bYHgR7Q0OLySHhf7MS1U92FbpVpOLlwzbXczjvp/bt3KsHAlJ
UfRQbg2MIhuU0Lhp0YVM2C59Qs5CWk2O6hCeidUzfh2Rn6LISWF8GIzi3MN3zFfsHcyEF5w/3xwB
+3gb6K6KssdG55VjSEiUhkEWA3zF8jMu8XUI6wAVoH2saCSW6LvaHE/kc3+QqiOQBTOqTIU2GaiP
PysEg2Gq3XoucdxOllZyykNw8IUC6bNZ8itKrwF+Kv0/dxm4aY+ZXgnGiZUzdJ22nhIcSyI6vOfP
QCLJgdYtmqh9gk5S8UZFLZfhf+udAuYaVOEg1JMDkSw2+xBcjBNktzpjp0y7xujqzzZ3Ndoe7dHN
mUErrGMd6iVsifMfMf4jqGswXinaGJxWL2edtmNgAQKdvYwex8p+133KtyIe6PD8Tbvdga5lZYQH
8hTJeQXWuLpIHbrDqvEOZM5vJrQghcE4C2C+JZzS9RgeT6FRavaDp6FgOuSwk58Si0B8i4Rn1Y/6
k0sqBQuHl2i8WTbOBV4mkglNIHeo/sYGKlScnKZc9TmGYnA4pnLjJoHGRpBOXCG/z849zh0LGBKB
V0kW2HRs8vLU/Il11jkYud+Ez/0PepDj/j3AN7vZhhYvjddSnqToLbgPPrKtu0ViA+VnM2IqqQLq
0ejS21AqBdDYVOCrJI61oxmqoqJ0xCd9ejyvhkAaV2L71BsoWU4i1FYXJLoCEnxctnfOoQ2uL2Vl
Z3iPSdDBM7/0XLawYa68JcnXW4XzEaz5avjH59A8RB9cRVx9NZhF4alZj0W7B4UHURZdWrpOY2ED
YP6uLT+IKwYaYx+ge/9Ng3Z9UNLxWR35aIIRqTPV+7XP0IVHy3dTzpsPaYyW9bZZw3CPxsPZfTdI
jBCisVLWDBwloeH2S42ToGicVP84llROiOSI7UxfeY7Pz58pVtVZMmGDrhIUPfNduF6S28aSQObj
gVmOqjiCrGGrhN3MEsb/UTYFFGNOjgShWYSVFPySqxaRxZ26jxJHh9amENAdC2QjQ9m6ZTdBM+XU
MZYVvefkaVXrddy5b9WgaSbECsxk0mKv/KsaydMzY8GlcUarb62jDRoLT7r2SaOyl0FhwjghH2o4
iu6uwpHyRbU/k7VoMMeYoeMIMdlSGOvEjub4/eJ8qxbI01/y3a4kjc+g4xaB/2dgeAV8RJPak4I5
dMI1RhPfwVzZjP0m7bzoVxtqwiPL0BeaDQ37osYu2NX8i+I8JgpmhTHX9dUx6oAFWOqZDwWBwAaL
ZG2eHyFsbve5+apstRrYgNCSYNp/VVL4EKfEOVSVN3l79vEmwm5vEeV0hIOKYrOaRGf6dGV4rBBH
Y1QvMGiRu3sbUGJp9CFLRmBjSdPWwkqZg9lBeN0jRIxnyQIbnzYsOEn8hTTWnsW/REhk+LS+wFy0
w7L3ZdGTH6ZDTzLrEdCEGeck9DeddhwtdPBe7/IWo10NoBeKykYPlP6k66J92wTlVKbMTRnWMlgP
bCR36wHXJgWjOkDUP+zhnpHiLchF5BIW4SELZpUAf8z/RnWqiTbZqhfUQC0h708gcQ42A0nmoncA
mSLT9mLU8x/slFqFC7kklXcYoByRPQHc/eET/dKwngnc1UePDL8H3WT1UmzCBJ0iXOhRYiGL4a0F
i1Y2eW2dLBVrgnBO+7XaRRPDSzp6Pj3HhUSnfBvA6A77IhCfQ2OL07YxzkNraqBGHxxu+SBlC9rc
uaqLGqW0wAxEHHXDujjn3DJmwbcz11cAuYukw9A/xa64LUl5S4iJEQ7g89DMyDG0FJZsEtLAtvPh
DSlkIAP6n2YMDWG4/NU4dTGWpT/8uaiuKBq3y12Xv6FDkrvhSwzQR30NJ6/NtVdH/2xkMxxGXkhp
5UbqjksCUTOPQs/+oBJlj/NQWi/YwxglzWVxfU01NoTj1B/Wwj6QCLjclIex+2V2ZQFoVt8VdPUn
9RxIDVstWwc+EFqpLXcaL4gyNUY5AL59q5k5mlFaUm48SN1U0vi39THyX4Vslcmn5JvV3huCcDIs
raWRorp74kXNQvn44/c1xv1g6zG0VctavEvZX2imF+IxjevJG9QYZWIUjj4NQ4VlLLx3NFTkncoe
/GxJwwVL6RmygUnVkxfkPY+xGZR4jKVN+9MmNeseCC9vUSIXDkkRLVFVWoop2yZ5W0VVowd+znoP
6Z55xeIP+ZuPwhINP38qw4qLLic6hIffB1YNvnpTYGznCnUfMX5D2M/MeemDKShft2g59DLwUTOe
/OudQ6vyKq2Akv7pmKWTsvWjUJmo1D+y6U7HfdkeCc9cUDLix50whJJWWKNofvxCHIlaV/HavJL0
9NlKCGfPTznvPfJS8LCuYpIo5DmZMKbFtTBlBk41iRG2UHwukyovBQ6wZAFNHqYHYsUruD7OMqy/
QE7vKVMnMPQNVioCIycHqm66shCzCziC4sqC9X5wN7kkp48UvBdPdKXwubrbnuutGCx+q4gLa3+4
YC9ISZl6/nhngsclr6Il4lDaqaSuR4M0ZMp4zsrqHEbJ62a5eA7T4hFFdegxXG+8SmKgkROWQHUj
o9uCj0WqLi6nfsVbVpqHI1NbM/HZeUSy4QZO0uB1VeOrnPKvJSEpTW3Jc4uAcVRC0UmJmCiUYd+g
QqieWky0m6alWzTVfbIXoOijhiBKUfvQmDGG5AP6uZxhWLik4JLhjVUNmDMEyp3/FXJQ7FPUGRH5
K263mDReazr0eCgWdKfUM3mHMa36VPSl+n+vxuaZEJIU+l2Gfz6Eo25zWOaus84demVSKX0v+HVz
8FE64Be9F9KaJoI/SjSeXGZzJekr83Ohd9/Xf0ZB+DYt+TV32Cd5ZW4P8Mw6gGI1KARj74It1gQP
MtS+VeVaGGBZ0wRItVKSj3HcnUcMcIwyAUqJoFZsIL5P1XzVEYadB3cjU2FE/CrKPBH8kx9JQQZ+
52NXa5uRiBjGHoDdy8MlB6cGGLvFSvfZqzqgaa2tf0Q0pWfn30OuEBE7OjRyvPtsdsIZ35QIwvk1
/cdCnJYGahH+7mba8st+RKEhW3GKDPxH15yW9+HnSAOfoxTnz20nokPEMJvNO9NvO8mB7tv4y7aO
8BUe2UyqZHC7FIUYIs+vSnft6utGj8b7HAe8rtaSj03iE6l16qjy5aW0GUtlER/a/ifVJ8nUQNfW
rOuoILfta2TkPL7Xa1lTHsX0EP7le2M0xBm3zmTFZVi9AcBmpxUiNfBXou/0kYWQcsaRCTQ8tFLU
USxgRjeS5VZvCIcikg8c9A+lqzhJ4Dm1AjmlH6jX46bEKFE8JVjNKEvbnFnAMGYMN0zyGMHvsl3U
cQ75VHkK7EvCqO2/K7pjPhfip07i1jaOKAsHoaoNFHQw7FJT9HCHx8gHdbTx1dpjmWVtqzp9lrmp
w8ZYW1CR7+FjgPG88YaNuOr9mj0hUocUZD+5IhHi8jQ/VwJXFoVk7gaPwpyRTdrwCkmDY22UJEwR
Qrfmttgax6fD9l+Sw7fLG1kOfIBBHUE/eKGWxNKSOTSLPFQD5rFR4yX09X/mnU0zq3g966XbLkHe
7+dGBvQRmRPnwfsEyt6qTlxH14timAXhZ8qb9CGggAKJreQ5Yz/97xliM7mtzuRx4uBQxl3S4pKO
7MglDrcFCirnmvsYrvtlSk3KuK6ZrYnb2hl30o6qeEG14hUIJBvmNsDWsBfbGvIdPRyEHdb8reW2
6Kgaul/krR0yKnk96lebIwaUagtBx+gOPc81pv0GQsE4Lz3pxOs2Wy2obiaQ7S+JulDcQTjvkyhF
QDzT0OlQLi/J1Y0CrXQsN03uP3w1IpGvpnpd1auO/e5keiIhwsME1AxR2Yb6LRXf+IJYjirfqFhb
XXi+MggKO9fRHA+gsl4KfksFErHzjPXByxx4tGAgp5SQYBIILeyA6WozVFpt2Uyu8BDrv7ClNRlG
BvB1RSP14bbzd6b3o1voqnV5NhU+8jGunxRYAlquFfM0CM9WWDp6ZsUeeBsv06Y9xCjbmq9yvfhP
bo3qS+wT70fZ+pwYrIr5ig+YxQqW0XxB8ePsTCEDmfl1lNZdYrHn3yFN3+Pujb8WutNLebnkAtyD
16gUSAl16EByoD/yKaxiDzSeuHA3F7mj3JiN8evVIO5B4SKGthSoDpzGuVM/vFExb8qZ9W2Xatd3
TTyZPcyoYFzED9bmsQ9ihZg3xyVdIgaeV7+U3y7xNRofe41uv5KwgCZa1VdlKQWuOagP6xYZb3UY
YtgrVs1Qw3Gr4+j7W/Dge/V/T9kRwAQCtgesPwmSFpZUOz32FxxPopek4R0fsnZYQL/PlZ/0/ZdO
wc6px+pb/5b7S89+1I41zYvxu6lw/Ib5Ty4nKeUZCqqkFJBHzDWYp20aA6bU5hxPh917pjEsE2mZ
FbGLgkSL6LjomD8aJbjLptlJw5ECCMddL+WL5RXRy8UiWWRT9G16HJ6FWvbi1GvGbbrnGachOWwB
s0fL7SZc1PyJ0wBGp3MJN+VQuP3ssNryozHibni9FldvJaI13p2C+fOMX+O4pHs+OhxvueE/b//O
KXvuiN+k/ExtyNZypgak75DXcBGf09VZmGpL4MLeo3SggK6Ohr3gW964VxGTiqUR5SlSS893nrTX
n34CnuWJ1fEAdg6GyGAwV9K+XHqNVlPJkmCGFDC3e1ZllaSQOANfGuUCh3kDXW3DXTGBQUejtvOS
hFgVgaOlzTzY8t6dIpbTemlahFt97DewSOsr7gyjhZHI8m7v2UOQ0xxT4aVzjb6++QwrConUCRvu
YSYaVqBOdX6uEUH6ICTgczNUUo5tUmhm8j18CxtY3lQ4I5SAtLlwt6IviUGQpOUlvoyIz067BhNC
wBxwj3XfMWsHWLpko1Yducqmp3TvterjImWTdy/DmrlIqedXqN3u6Edmtabpdym+lU5GmqwV6InZ
DbA4dWRra7BiiXAbFV10n829w4c9zsAEbiTNPKmcuw73xJp049cYB24C9QDUVkgU3X+yTBNrs4Ed
CaGClPdboQGdZMJosJFkIpkmdS6HhOCIJzs0hl0srTboL7xeLLk/hHCLq0rYD6c4CY7M46pgtlur
47t5B+cF7Co9kR00ZMMVL8GYnXqsqNkydPmAexyoLD1MA0f/L7Mcue4A1vlEi1L5yTnGLAqabhM8
OL/jk9+Nfs9ahu3FoqLTh7Yt1aYey9/EItABfzeqQzVcVXn1ia2W/5108/wvnkGUB2+bxTAxyrme
bDlwfUv7iM9do9obzmTLjOX7Dyyg+Xr6eDHiZME7h5BGls8+mXWeRJiM95bPlINwEnBnkPfa8Ctb
begSyZ7b7uf37enlhnGaoEoTWO2zae2mYR+iYCLYa3sJt+CKP/LdxtbcV2Iy7hsBa9AzmbRN/KDf
ZQ5lBk2YAHVyFVTFZ8t8l6gsnA8/SpyEfwwDg2HZ8SCdh0Ddrghcdq0e9IDDFSrYr7xAUoqx3ETS
paAnOcBOLLPsO/4om51DAWO0n2TKfe+B5366KIkUOdULSXXcHP/saaWN/nQ89Zc7/IDPD1x6MU9t
2aXo4ECKq66FlOOoRBrRnahHVHkrmgbHgIVIexOTJEunUn+/tdE5aRV3T/M9FNMXm4ui6cuZOjuN
+C4neGiRWBJ4gKc7FwLK1OGZ7Y2Op8q+6SKOppwo1qepXdCuBq3Ls00w+IXmqRhrMyfsJsFX2LVc
JEuqhcoOOgX3JCGK3UmFTzTrLVMCpP+Tr1a9k1T7FhpROL2n7v2a8jblS7Lr6zqCLuCJ+JN6REct
y3gR2HKLmM4wlcoGwOFSXNNOY4PNkmVnucOOgeUQGBQkxiCiFIFuvvZt9PKxdcKA5u/rffT6PMLR
aUlXR6LDgzc1648yxQ/ypRHtf4AhfdMu5P6xDshrCnzyQ3N/XMpi4DnTTvfOrI1bSEOxLcn2t9VW
8IuXFTE2iaULpyvZTx4UOUchXCqBBazitF38I1XaHzWks1BoOZFk3uDSmppFndGYh6slcQ4JFxqv
XbHePhCBxUl/FQI7sdj256uysS2jvC22XmpGDxsrfH5ZKShEudJotJKSG/YJCc+DMrtsb4uyKrDk
07MFZxjFct0uSKvvNWXNCA4ZaFFaLMglt4YYhZoqWmkAq70Xwb0rNbysjYblUvrYv/KBfalkkeOH
XonJuK8IGppHEzR1xpcEXxZQSMN3Dtr1uznLsySe6tfrJE7o++4CBdwCTCNeGX5yJ+a6weYPNpPi
t3F5NPKjBB6KOrkBafIhlhLEe/LPsm4nxv1FGue1vVa6unA1+/PEKjOvh9ENRRVfq2AvFxYGoBdH
VxQbNnQiBogZQS8UNrUsPOysMIPYcqo2IhG6/DN/ASODrReZiHwquebem/2O/fTVyH22Z3htpsN2
cYHVPe4vrkaehcCWBbTCUhBB2Q05UpridfaW7I3d3gfte5bzfjCjDMK25Uzd4CnOUd4EgvKYuhWK
KjApwqPTEjBDeHiq0Q3dkawOfOXrdrS3zmnGZXWTjfSJGM2Uz2Pdz6YK3xFbwVt/bkUyX4d0KxHD
zjTvPDQDFzK+GQ+tnK8bd7od40YHyuxtfu65IEKmVehKP45foVf2pIiiZP79veLVLabxtbVSNuzN
EELn5oZqe6gPUGigyUk7oMxKIKumU0llOOy+6/BAJ8ICgf/3JOnSpSh3ofWkEPzmAZoW7v9IbAvU
BKU5DWIFW9J5D8IjzFtiuKM6ixjcK3ZSiFtVQdeTD3hesV8xmlj9MicIhQp0G2lgUj77YZa8t12y
D6mIQsxKXqVpSVEwLGibHE31krSd/s7vpiHTMSACH0NBGGM1XoloJjbOU9rhEL8V6Nmc9+3oVEQk
TcVpS/yvHcIWxe43dErzXCEm9ku9s22xWvETHJ3JU1QAcVh+7exQruz7WtD7D3lWsmSqrWi29VVn
zTNgw9NoOcMpdSB+X1QKjgM03jewxuJ2HNfrAzbGX8Lk4xJ1ubVbnWeJSwUn6YEEEugIRMy23yWT
ENU3wosUjd44W682au2yYHnF6h/XL18tJ+ooofZ2fQgNqhP7tewvpV5w3q21MsrJuqhwcTMBVguW
kpCx4MAVubtrKyQg3LnAWW2kUlBZEatXVRIzDBS630DfMIIcc+fEUFYGj96PTZVhrHsMjqOiEtR5
YteQOn2tibdOEj0soNhDw+Dby1z//0X7ebRJQeyDxlVmDZ883U8p07KqDB+dT/x6bFlFWwrh+zMj
cRu/1znLQTh+8wgTj5gc3CNTKEEowYm37xCG2JaPh+iWM8j9+WDgBUkuN/2gcZ2gUtosNpfFxhDg
azSAW+cYZ4FkQUNTYvctM6v4u9IsU4wY+IyLNN8oKtI9vRg3MO05OtRehA+Wl1fMLDZSVY/Bo6x6
D3eB3QhpYpzX8LbklCNZsKJEULwE6t0lg41freJcfTL4NxxqfPYmRokK22NoTn13+bQUp+a0/B8Z
+WhzoocEP0RfCIdMyj52cTe+pRrw5800hpyz5tWpSiye9ikt+bKnGmsO7Cz+YR4UtWGXFOCUhVEg
wSX/soXlim8lP3deB/eB8VoLfUpW+1T7bhosfpOFgk6xslCBIKQsj74NwIs+0gx+R3nnzOlO6FIT
9wjplVpf4zt+3mLYLkTwdvLD3n1mF86d8qSSi8RGHnihm8WlbBuggDbX7JZYWGzwobQ5s86rJjU9
rIT1NZYKgLCnLVwknjdJnPXM/IDUIBgBY8A/TNmW8Ygnc7CcnTa77eRS1ehd1ps+DiX+em43GKSP
ifdq500c5CPAZzEyZBZkaVswv3SGzjDfuSNqt11z2/YbsuDSBvhazGBouRU1CJaucC9NdYYJexOI
mdE+2T95Gj94LpO6LuZLqFqt69E7oq5Ox3FH+ON+wSSxWebMONBYvzqQ9oKSlk1Kd0wzBfiNXMhX
BYbjhgrOEzkXKWPn2tJTtDjvMMGG/GSuD/SuFDW2Tu58X6mJYc3HOw2WDUAIrscXJqi5hqKQbN3G
4+wa1U6iIijmkb5zhG7Q9TiHYi7uHU6+GR6TMloRMxdLHpLmYrE+h3w/KDbQe3e6xYaDXpe30G0V
lghmUHOTj5AufitMaKcWIMwvl8NvO5hAtSQvfJEMdBIctVAiKvAyryTYx6ZsNqV5KwWZqW2AifYh
UPXX1PwIm/9kmM6gQgAQrxN7/XCFQtFqcHjV/437125g31tlbXSZrhLu6g/UedT1Cvja/W6dk1vm
JgUzlaMKImzia87CN+IKNsquzqSiIT8ycPr22PhBardePOTCAW71wGUezaU/Erfr4fE59yrlYlI1
dKAwN0xeACWdAT5RCUn+MjF3whImhA7J8HS4FsBS57EE5uvBQ12iEE3HlO8DH5t4rHyc/JxE9lPq
3Tvghjf3YCzH8ThVklIBdIu3LFSAXeyPoFGeIrZWWPmOPVMxd+5K+lmUO+bsul69vSRUv3ykRQFP
AeJLFLl16wxy6nd+AxXhQnoVQcmY9AqOtM1XQoj+RGMLURPfnztqxG+ajASyiLywH7PHkFoSB3cH
Yq/Aaok//n81ACQT12z8MTFh5C6BrQyfdXcFoEfEAx0cRvN2HpOufYvCsZrKISnvboGiN5H8JRLw
S6GPDHHhyCHIoJpEB6N6M1SPOGZFk15rGOaODyIrTFunDgI60Hot+MWIg6FOJ2BYGf23weYxgOdV
VlGIPftkhQ3/MQNqYsDGqzT7pe3yZnjIeqHwrH03lf8xRT6AR75GgKg8+8886ikhTVsD6WJD2koN
IY7JKOSPIlUtdqv53ttUUfUUc7E235IWnOYXLBCPPpWaWT/pyO0A7slR8pJT+7Ize9UJVCxFrBHB
RzaOvsJIpxqxltlUqQdhY3XMlQsE3x5MbTV8E5wZHdndv1UlMZI5yB/d5x+8jId200BWJsKvXBmO
Lti5OufdqgONVCWRinPEId6I0YPJdLsDtHkqDZ6XddJ7Uibkr8NdLZyuoCQKd2yi0hVRxWFvTVeg
BVu71NzDyHmtiA3/9Xwdgs7CTFjWsxU7SnvsQfJzwxQKr862w8elvo7Puo9krl6lIYiYEO7P5j2U
xz+6ZlPxVHYPmJbTUboDBj4C7Fhfq/a/SxG2xuQBJtFU5Fc7VOiWIETmkmdypXp3cOejvQobCK59
XROc6PWjdpHHa7EyHDq6B0C81tFMPCxeptp9v3ZQRC02hFqQoyV+U8KKjpYKONRr1UQ7fPVeIPKC
UDKIEO8Mqw+xc85dOuSziycu97yjBa3j3CiNCKdXnB6e724PEiJMYX01M0umYSTWjKnO7B/8+IY9
GbV/w51cTiRTsrR3mUs0aGrV9rjIYVuFkR0sxoDg6hIylSiH749nBpHHcsSBt6tmtNZUTjGIy21r
uFS+7TacJmRTc8ofRH0c++cuEjiQQKiSQuSoyUYAZMN4fXU8iBlUQFCXWMuH7VxA608by+ua7wFa
b409aZHLppHJ8mfswfvbpVzAvdPs44kSKNzaCNNCb80NLaCjPX/naDCint6UnIEVIzcQDj/u/sj8
T7a+4UNU4nZOo2/Hck9dEhU3nJJ18ew9+jfu2dAYapgS8hz+yDrVdmcg776S2lYQrFag+PrCHaMu
Vpswn+6wggc23lqujshsB4H5Ly2J1fTn2cNNXNYMInJbHwR4a52SfL1jdxGIFqYNbZST1GoKl2yS
6ppAfhvvsf7PjIEg+INXa6yY+YV1FOpSUhh0A/WlOn/aEuhqHSAujr8rl61aZim8JnN9BwcU9/bY
dIc4ttSwri1Qa+UlKr9dQytYwl8l8oJXnwOstx5Z/4f5QAimnQyVbZFgo3XndfHhg1pyY8VvnihS
tqTtsrppm2ZsU7EepV983K6ioe7X8OTveOB5fG6dRBrvPhFvTkmmwcb69If1EGlBE9lo6jLEmqw8
pQ5X8lns6oFlZHSck4zeFEItQbYjC9e19Sk5F7k9bnxSx/wtfSE4e391tXMa9EJR+Lb8Rj4qzJHq
M6mgvH/jPJaefYFBuZeOlf+PU7shJb8rpN1hM9bklRjylDhNIGFOS2csvvBQKsXk1z7smyI4YyJj
Z5rxdLftkS+ukzEdbqubQnqnaXLPSpH1OFpgawpvgfQ+Hn/U1H9/Xp0QFlVuVzCSwp7K117UIF1a
m4p31VmmGXnAkidBhYJw3VIS2ZwLVOASSTi/r8hjKWdqdOyuPCRd5InEjtt/yfiAYLa/0iQbFd+v
apJB1Ta6AYGfNxg2eUJuMD2d6HcKIlGqirSlnu9E0ei3XBsyQYN9qGTi3dstd3Yz1DZdeEG4Bxlu
HNv+t8+gfSKUaBwnkwkEqZU23YfsuyGCcQ74KiKHV51RgmMuMmLj2tuxNqSX1+oCWlCzFurqHbdg
SuczV8Ep38qOOmALTkhFSM2kUHEhazCr8m3C4ebf7Va0yJoIRNRHGOBZmAwAYVFeiXONV/gU1YWY
N3v4/RWzKP+JYZc1XHziTIH/Z2nnjlWrT1NuPPt4XGNJTRL9Bv3R3VGF2rbjBXKJ0PQqvSaSMsAl
idl12inqBP0oZrkO8CIRX1utpPkiobH4aJ2WUXG9tAByHhZMm67nnm1ekSulQLpgQyjPqxxOcmxz
UZC7mj+Alz0HicpxLmlbcQ/9/nbI6xv/lwO4FqFA8Lbwj57l1VOt7JVr+YLv6/zZvIwmE+KV04vd
z9EtOls9Hp+W+MpvmyQfi9bOSY7uiOvr9c+esZu3/cqGy9P1S0QfJJGoOETqA6JNPCueHkzhe2Ht
RGdHmLajJuR6O3wugsf22k+dxNFD4qWGMfk6HxXa4gXULGfhdUKaNkL/bjzFK+mhWtcbh3w3Z7+k
Q3onJHF56KfPBhzIiTw98+GpeZ17V1mJbs68kcDeW7pqNhWtCu4qLokaWCKJ4z4Nbkdb6HJ/g8ih
jDqkVB02o3zwkThNmJmUL5q6u0u+Vq5iT+q9RF30eX+yMM71gvxsRp4FJP7qYwBX717FKtJhIpha
wphtKVMZlUHwhFI7VRLo0v+n4H2K/IDxxh9R2RKEpypeZ0hpYD5Pz2D5Mv+JL7UeinGykA29HlK6
x55WZV0lUk5lBXyw+SFzUsxuejYrliorh+8sd8dqBGY6FQKM1Ax+jkrw69z2wNMrpqBS2XDHKLWu
H7cuG6QyfDiCIWtA7M5LpWb6bgR4PGunM7+bi2GcZAzvjg0p9qwZiXCOcn4kx2LFAEIdNoweUXzn
VvtD9IEkGYg10h96CmNS4LwQFyJiDUHZjMkyh1P54fFqtbqFwlYR3ZL5SVn6ESmNhCrzpHr+kI7R
AzboAU/3iFNdzMx03Gl69q6QGe0jwRem1nHojrKfDIvBJsOaS59HTM1MXFwl7J1Jm5q+9BzXQ7yz
7bnhrHLN2IGZig8y4DNpXTqudHHNgWt8IVbq1wN99/lh0bskFtu/98eqLzvWm90I8tGYbVXTEoPu
WC9LQkMIhbelhqKcp9/yu1YqDLeufzeKYaeM14KG4xl2o+sZclcDFI/mu/cjISx4iV8MsAEW0nDd
XfivvmGbYPQiM7Fb2eW/h4kJK2d4aHddost8RUO8lKsZp8/k3I3Lk6se4/88NN4MtLLfkAzrMcxy
KSuwr6cKmsPP6GyaZaXN3zp6zJz/KoWm+r1/2uCvbB2Fi8Fb1u1hOpCEPE+eUzGVXaoI6sHg1WsI
B2RrGJgQV7OVKxkkZQz6zLMjI8wp/Qxo+HOpd2evNw5+Bf62+NQGo5vD43Fya+h37TF58MvcwRqd
PfZCTS7hfGaolzWUX8hnhnH4kQ+lAeAzDImsihjG6G4i/HvNoRhU3kU8DKrCONDok1FjBue5Y9IJ
IgQksqGa14XgZsY9g46JYyQd2WNJXTWVl+vMZGzgEXuqV3D8vURdyqnUE7/8nATJD+6aIUM2NymT
ZkpmGodMVjufg55KgF5RyTxSwgoUAlv1dURhOAfa2SyDp9qkWrlwWE1SxN7Vav5Wacgg22HIvoqj
lDHiH/id5+iqnaOYY/7fbC6QUHdFFEM8HPbT6EwThRLLzl/UHaClMb4gUJ8qwRxNGK2kiaj9yopM
YCIqETGYS252m1pXNF/JjhVl2GJl24N0BpHJwi0ijAQW5v30hauJpKWQEzQh8WTYpJWV7zimG1ss
WpCCQqrY+r3/WHMSlaaqcDcO9izHjBWlPVaCyojHvHN69t/Yp8UsdODuHrg1fFTpA7RbQaew4rSY
HxvvG9+ELJShdZ2QPjo07zBsMmQfCb2jLAcXWnMSvbC5a/mURiNU+aNsZClO912M+8czopFSArgj
jgkZbxAY59+w16xuNUvTNuRY2omciawM4kDVBYbWvw6bIWvCv20zsLCg4wSMfSbu/kJrlPVOWm9n
sHCIrS4wSRhvuWxQjGYh+HUXh/UzD21rIGR9wE7kNKoVJFUeB9QmtrXXxOSWG/M69+hAz6M++WrO
2x1BdXUKUnxg6+XRDSmkTw9J5dcHgE9sLvRDh0AqI4t4NG9qaHG17n1hrfS+druCsCImhYO4cJ2n
dUhMvpE7kDFuIk0x1koRCVUUEUBbFFQQlScvVszxYbF6Vx5+bIiwgi1dTXTKiL/X+ECRMZmcHshH
lwjAxpLSyWO5FjkLbLS9Mpu1VilcAocw2u/4CZ5vJGE3Je6GS+/YRQ+TO2W/xN5wuvr/pBzpecC5
X7jgvgsYEaNpHPr7ZK7/BCpvcXFZp17OWTwL0MrMB3qEKnBfb9I73GUamkL5y/qfxODNyVXbV3vo
H4OO+awOZaHL5Eh4bnOSW6mPaENTHB3+VTNO2IsEYOw1/r1xWAtSvQ9Ek/iQSCxcRmBo8O8MkSkw
xmwSYZ6Tjm3b8SKF0FA0b5X2zTax5LfIQ0cC6OTeL0ZqizgXcTN94nDyFQGYQtj9rijZVz73W42j
16puoNmyb8kuZp33IfttWZY6lTcXFKMwBXAs0jRiw76BrgLVhIY/U4J+QjlDLYa6H+vxhzxlWi69
fxr+qR0saHSl6jD5OSCstpuy6mylEJ7VKr0O1V87NpqAgWPUpRR72mDvtVXf1MadmHZPq4DcCi+O
6UUBF0ZYCbKARga3tyZ2WkZwjF7p9GpEAT4sl3hBuyNF/JOKZ0aQIomAxhz+H3eE+ZAGjuMGdO0Y
IzEAdFooYuXycGBGFg3DiTmrvroAD096IlzACcABCVYTkFbybecE2j6LGfR8Tch5Uz6F58GyqoDo
WmiM58onUSb512nKM2Q0mkfdZyDydtLtT0ItaUCAeDGPJWUBYxqnGGHu4cIdUc36+VN9/bnRD5zM
PF7dTW9FXT9iqyYFLLAS+8QZDMYtvtMQcdo4Z+H9LG9mePujRParQHgtqR1jqm2AI/xEo+gx6fK7
crQ2Z5B6BLZU86qspZ8M+KnJJwc13ptrMnNCFd2RBtBNXbA9XEYtoSM2WmCFIKVbCEW6LjY9KomT
02/BTMF0vRIvIBJleuasp2jgFF0tjzn8iyVcoMq6Jo7o0eCGPitgJr0mp0vbqHh1Q5fB73lXKD+a
qc6vQ6GfjXnA4ltu4NmpGMU4YLbEv3rLLbSr4cDuOonO8mgwYDxW+hI+rO6SAQSjH1TX76x3yDWn
7rjDltjHEixdfa2iow8+04OGfnjV/F2XQPmS8SS/f7lgklr4scjK9oU7ZWTuj/cM/qarbxY/NvFd
uVltiwVHfyRfQC1ElwfY2msiTXOly7DWEsicYC+i0f//z4IBk0nxeb3gvlCF/rJpePKo4nEItY+3
IAo+ovAZfibp0JlocRjapGCVEbnEFEM/5OkRw+2otB/aN830OPStzj03b4p4kJyUiM56ExPhp2Oz
XBz5TbHRu5d55uG6f/nlWQJ1gapbbdGsoyJ2UqivcYGjAGmGOyyV/QKHsQCeGsVpfDqp0nlyXep3
1Y3KAfsGMy3d7hqSdQIBDvNMozHpR/4DDnqV8OWKQpTIKV5N/uSyICB+HJtDx5QDlseAKL6mUdnE
ReUJIe0jDKTQdc7irw7goFjJ1ML7YqO7r8IMMHFrptmG1yQW/l9x4S7FJdF0t7gfI5e4SxciZ3ar
HM9lX9TP1qR4xTz/3+1Lol65vmGsY1z4/kpEBH398B4ceU746+9FQa/f8cju+RGZLcJNhahHVF6X
wDfmQQLQrN4MLkLAopHAFQTQh2TKi9AHCI5+E+5+UhJim/itTPWxeCxEAN0DUcgVXx4GRFJ8wcBi
jS8iv/pbfddv2xIBNCpLyRQrGCZ6ETzt5segXBPKw4fxIs1kPQmvtvHHQ+w8Q8xRjFBiVdIvms7B
Jd1PoIQEhn7qE0FnZuMr49KnZ/OoUamByC9wUqZPrMVLGMx9T6uWdnsnniy1Dwb0qJat1sYAxfDJ
57Q58aIdbJdgHjXLTJdyH0zB3P6zXVdE4s7iMfE9KtKf+qUP0JGU0HmZ1ivM05S4CmJL4W56Fi+k
klZzU9NwEB5BIlT2TVUuwopKn3GUDMuydM535bKZoTaQpYzUWK9wccuQULSEzoFQssCPu39wjs+y
DhaQyWF4R3Z+UhZT4sOqM0dwXRb5kCMZ8e0tBMl5Ci0iXxrOZXIrT0iwR2coPVRVOOXvO3C5I6m4
yS/7n92xnjcoygv0VcO0IZzv9yDr9AxvQR2A/Mvc3yeSastDfMeo77yRp4ankoxyr9fxmlurcCUo
NWHRKoP1yJD+G485d/GIUEoCMHCgUdoe3IVI07HR0MrpRNInJ//m5AUjHpgB8SqOomBwowhb+ht8
GlPM1PkGzZ88Al6ic6czAHMfkxE9efF+ZB4C1LnrjmZmkoyJhktCNGgKZKECxPPas4ju9j+mU3SK
ZE3SjKqGAGOSGL4wFbSCWF1yeB8G9gMq9rj+6yYmnnjtkkEYN+PRm3KcJNGb6ulN1UAdZk3eNetE
OpVC1tzghveU1HrDSvElqj5LVdsVXs7bAafIptyQdcSc9Tb3d0wMva9EdIbUjWLXnSgLV4nlXF0O
fXaO90NQKqm8V/5IICAsUoKMHlhOAhEK6a8CFebDCqGYPLhE4cN0pnMK05QuxUwPUtNmKYwi24yV
Ks2u1ENH1/H0GgGNG6px8CJAY5MqksAEhxk1dsWLM8iSSLZOjneqwcN690ChAXhk9dGwyZ2UHZ+6
PSEQuovrBIGUAtTOruOPJKK+jpWSB8iBmmDUSISNr0qyKF4oHTitvDf0tYkk97IILp34i85TV61w
2bZdQvX/FKWOJPM+aVqS2YJjfiJLfjkkYVb/c5L95sBQvXtKVp3clanJIIw6eFnYI95bX92SaM6G
aukf5ZUpXY/dNOvjF8CXkA1dP9xY3XmPZXwgQ+dfrDj5GFHrrUQo4UCFipMVv5yV868wez1kml9/
rL1owmSqbUkEftyFcLAU/Z6AqAB2TS/rSwsH5gHmvOd3qJAqUW8pCqL+Hq26/SJJ9kXQ3U1ruIjx
7FI4EQ9gJ/KSghCFcc3B5m2frSDwODH67nLFkpSQqYytGxUF5hpmpggqRpmpffCJGuv/ZzQpZbVy
J3EAkiq0l4rYhllb6qI17QP3oghOKjRed6zbkAQDGNbTCmoyVgA5xDtU3uCbkKKi0rd9OLPu4wLI
TEgbWSmaxB9G7YA66i471vMEP1ulplSNRghTWtS6OwU0e5IlTfGMeMbWJya7qwyo8Uh2XS2vjrjz
0Q62+ZRS7IR5/+QYnk3uGpvqVlgA8whnDoeXutFy0Fpjm7TheY56gP1zXQlNzXFNlHvHop8ej3k0
bZpHmTITXjTJYHoNc8JTufBRtO/Vxn9Ml5752N2soK+7vbQdZYnoLyd9va7vXgPO5neBkje4z71h
7vggwVxf4wI5fGus6Kn1PdigTxalminDlJaf6xZ1JGL827jjk4sygdqgprgXHL5ynDwREjicMtOC
I7RSSN0fMjZ5m6DwXO+gctwP/jTkeIG7NAIV7YNoRVfA23P0xZeuq94XhUP8yGpnjkOUBwQkqICC
nivj0drWslpnzRqZuL1Tds64/Q84aHSb2Puqkz1FEdSy/GxGhZoYAPjuOK8ik771MccVLjE4Ine+
C1gpBPXAi0wkq5ynpMZl+greYWfPxSitYu9OlQV/jTjPCGXuOOe8HtrnRyGQQQl3mT7ZpgoO5I3c
G7XErRclRkc+JSiRa9eLViVH5egawEcXCPConVj8KquKyBvCiwRQTE0XUIet1XEBZHgo+hLlE8Vu
qRguXYPkr+2VUBwUqch6IK90BSIQEF+EM5AHa2A+Hq3rbUxePlHsjqx7j22Y/flO4RH5wIQE3i1t
mhIi/3ZjW4x2pAACQNESpJB8gVPtYrYbkdKyFqh4Pu7b+g+PpfrPxsSELMgey2kHydxW6UTSSSxt
MbOxMjhMXmtcLWvaf8e+vcVwyBK/DfxvCGHi5HfFnebwmp6suJ+xVbfqQG1BNj8KIITRLR4dhRt/
Bw1+1ngivun2b3RJBl5+j8gV9WCwic9xJANF/bZM2/YEl7xXKkpQLtmDJHBSDo/RtB40lHfk75eH
0o45pbFE+Gqbm/nZSSVcQZPXBfgW5QF+dnU0KKDCkursl5XwZ5GhLuUnKMQ9XcqegjZjMHlG2WrI
34gtS/UGD9YlU0ixRAt+b84cQhZWud1+FWwQIctXvqPHIVvL7Q0g9NlvoSZYglgSWsjJsBCfzN7M
Wnsl7tFAnjhnnHX0PkOw0KsyFbcUcyf00cXI22bADwWSz/cf9+exoqVjrzD04IW4pCDCMhZr/m5M
cLaGl/y6A4/OjEFobCIzXW3ZpYjhiaev7rE+shp5jQvwNa2gtjfkz2/5OijV7Dx6ldjdKB6e4eoK
itpyBIFZfCeIL0lW/+n2e5T19k8ZTmNgmH+HALN/asTYtaV6crMSHshvFSVabXEgsuuxXZ7HPZZt
CNyfthZHHF4U3DO18KWL3aa3o/ecWl7WrhMnHYVMwS3w84yF1NqXjwfHanKhN85y59eEj4iqdc+j
vOwEmNe/cWiLPhs8INAKb0Do9N/WYcsYRDxkZA3izkCoQ8agcMY3OpYgViKZ0NSK3HMOqZiU5KCg
GZFxIx2PWA+9RjpY0xddKmTgKJqnztPG0p+aPRoSWPXkylqK2Pt6O45NPZb4WUGDx6Wvu50O4eFe
8QDRNIN5eOZLD6/9c5WUr0YkWLgX9lf0YBPea/Nx7r1z6YVVil4TyRUplrMfTOn/9TmwOrFyn1cH
G6hE2LYd9kCDBh1f5r9vnvi7V1ZwXyO51euVWDfQmMBCSbVldycBojCqxOC3eiLpdEUvIi2rzQCh
c7+dj5KVRgGJ+Wdl9s+Gr3c0cAv3eAjNhIxO69UWF41cveUwhDvVHfraTbOCmR2EGyXcIfXvQA6C
jTW0Iiu8nHWkYqtordJiXzyUldRdjL0yTb2/UmeNFodcM1lvT091+w6iVBCrSCZwHyQUJhrbEXSS
gkHjtxrNZdysSiWzf+nHyb/40xw9M7C9nHCUq1ts0bnF/hzk7TQw3FR2iyJiySD4N5BDeUx1Y5VG
mMZg8aX7zRn2FliYonJfG8C9FBrNzkTEBmVa8hxU1tEx+FkvtojcnuzUs/24vVqDS13/QK1WYkwS
zTxPETdD1i89u4XIedKQHjY5kOG7ZvB7LVRD/ShRDq8K5aycL6/lym9Jsa6bf75yP1NAO89G4y/6
AAfQSNEY833e89UoFPUGkjSW3jgwwnNagwU4YJJHKFzDRGNQ242gYSMigvOld39hbKOboP/inv0M
UUNvHVccAlc6FBLBj5V0jWPJi6R7CZuArMX2UVrfSHpcTJwHBoDqB5GnyPbUaQ+CIykiVAhjGRtu
uXAkEmQvBBut35H9SXZUCEVjOOGES4dJnOfPkKCcATY/AEnAT8RtGCj+8tnopFxe/5sqRxDBHwJ4
sR9Hvu9cNm9FI1wVU/RUjh0DsIEUP25u8Q36ro4g+nqvMMA9NtmAXnnZs2qDeHLzmhVjSmxfrqgm
2kTLqgAPONDS4/TCMywbnllzdNMAl2JI3U6uBukYml4alVTRuxwUWlScKd2loq9rf87u9DYEoR0Y
7qFR6I018Bysj/ZYNTuMcjL4KLfgOLLDS25O+gHeBsiMFRITv2n9t+dcSNpjodWXS643WLXmovhP
+Y/IDni/D/W2fLx8Xv7ChrV8Jl6flq31Gj0DNXJum+HCTcrWValZjZRkzIPSV/q7vHl+LT2gbWTr
bY8tHaDyspq5sOpdmKX/rrsSFRLnNYPLS3qTnu2hw7qIKlbj0LKBmqxkT3NW+5a4Hpv6tfwHdrWi
lojNEzJz3K+fGw4Ix0UiV6YXPZu410KVTNLP0wXu4p0vqLC0TSRtdjON1O3EdZZcV23LxMDbpYbu
+ylI6Bsa7omqlnjcm8n1hOHbDoHGmHWGz22LpdHdhCoiNpbHIXRBzzu2WWSdMtNxCQX12lwQJg/1
K/TZ+MaTjWhAe/fld8gx2uxYNcVNohS43VdF1WLXX4wypKw2/r3K9txBrFEVHla3jleKfXbM9SwB
JoL9T+h8sAK1+T9sgPrA8E6SeT5cy+GtSSQTSJWymliIcoidqYWrGkhwUTEL97sP8pZz/3fFwfAE
jyMCc9mafTEcdY/mlRELAbJuuaupfhXfCBUkYAhZaYiXNJsptYoGkEuUBfZ3CsUSs55Ss7fvCMiO
fDoqlBUEesOy45uzJLFlJHz5GIfVT/XRO+bQxflui4Loa+axsENlVyYxk2q+BnMoT8RkBUHndkzp
6s/fdJXOMvIazUlFNPX/5kYQIje1eF9eZqVxHWKYv8a6IFeLQrX1jhHyDjw3wRuDPj3KdJqXOzl4
lrkte28Ko2r4N0x7+K2OryEP7jtUDlXcHtsaXFvEsfOUQ6S8B7ywW/usj2BqlBxSDjNDly6TjNnM
1Djb/tnIB7v4zLjIFyUaJm2nxSEXJUJ96VA15IhRo71AjdW0/4UyV2FXz8QVA6oFNcFTnzZ7H1sl
vxMUk01Dp4IujZ0NokY3gr5HzSAVqIeSowmRrIOT7OCSEJqe0b+50IUe2tMCd30SQCAiyimpGr1k
gYkNRlfz/fg4bL+rdptg9YTycwYpQXlwitzeDHtFw8moqNlpZkrSZjI3aKiMrvn1leqKcpBxa8ku
Ld0ZfmDBofx4ZLZiBVygIv734R+zcv++Wr9naVKb5oBYP9G0YHaOeq6+9SSdVUj9gPfsHQccItbH
BZZZ0j8IyqOoomFxBEcigj0Shuc2HLiPBn/BKg0p4ww6UA0X0qBF5wvHtt+tZpZ0y80JhQS7cv7h
EkTI5mhxKImgyQEyM+lfg3J+qG4Aoa/2MAobYy3/y9A41NetYFl++xIzmIdfULn0uaOHH0FI6k9U
Ms57pq6jRqzjkythpDIjJV9GZ9vGTD8HEL1olME99cyGxLWTcZdMpUso+5fcUGEcLyaOGJ1q9h+2
WSUegIrzaoOZEF8XY8iEtvfBGj7oEhQP53SvZCb7O8xc9eN4cjGA45Sc/smW/y56/Xh97v0zjXKG
DQx/sg5qPLjTwkiuMmt/dv6POF05ebzopo3e7z6yTR3Mjlu2czoP53Q0hl1vY0aRF+6boiUiZbX9
ubh+K6HHtJ2XLMJh7FTpmbMYnKeMQB9qpLxTmwehuhWQsNTGXnngjvwg6q49oPlhjDclu4vGSAfe
o5Bt5phZzT6rGi0ZUNVoba7l+bJUmG0xEJe7NWsRF0y2jkZxTNIvREbX/uE5tKCQNrrOTQJiXGiE
kk9wnFt6ox6kzu12FqrZg2NqgS+5LKpw2aejMLdQIQTcD2NxZSaYc1pgq5H268tolUfPh35vLV7O
LUTGLwLvz4lXwmSDIS+1HMEnmucf6D+W4M53HLH5DXnQ1G50h6JQ1WUeQVHmArg6AAPfGdgGF2yT
Bmeu8UZCipP5nA636zyQjtGiWKRXsB6V4u3oAQ2A2KwbmrKs++mRbJKTpVApyBHOylRIrqPb4cWY
eyitpv/tYaaU/LrXphrm5ARdK6VEGxr5MBWXJfrqrLPfs93GsHcaravLrksostAxu/+i+0JtLttt
yiY7brgJ1z/66jMxzmpJIzUE5ybNAk9++5AHFsA3wYcAXwXsT1ba0FizPZmM7BxV/4zTbDCvQk/s
jiIoxBd8h4RTVzgTfETDCfA/8uP7xK7KUggBo7kG7l8Qe08ZWHK9OOgc8Qn4rAqQt3sa5XIEJlS9
jwjojTJFTW8+UPgm+PMWFOz14iVCUPdTsVYdrzUvjoaeUTEuVWUiu1nmq5THAbWu/PMGAFJgjdF/
SZXxav1aURbezEsYD6xo5NY4ihCka1GGhSZyFhGPxLY9tMvVrP7cbtkiu8M7GSj/KZNP8q4WRUCP
lxsFbAeyD1j0MKByxre4JoXTnTmpvrSegauyT8wWUfwGbtr2m500k7XK8kzQrvpx1zNy4kHW+piU
i5wr2UV58DJQoTLQ4y1ggGEd9H+o1eDg3M+MpPJTJQkL/dTmRBeg0lc8M/LPIxaa52C0SA0uDaLV
kz4stWxv5jvEta6TrCHoe9MCO9UIkovjbKkEH4QOq7QzYAmjeLKPJpSVGC9Lqqu1/mwW/lGrX+Tc
rrqNirzfdCBQTeYDaRgLkb+Q1RTjBeggio0ysd2DKORlwXPua0fCMU/EmDv4wlJY8I/aa9FS+e52
dNidMXH4ngr6/6x41m1ZmFqc8aDat010a9/vkkjxoXV61PI43/agiZWKcrAyawbybthJcG9tVYmY
xKTktgESe1bPO6ZLOmxyqCwnTpfN7S19WxuwPvbs/W5gIpOQ/qlLdyTmjn3xQ40uPFpW9GfYgStT
+Wf1qZcQW31UV1JdE53J8JKHrE2/Klf2v4T4URC0JewyI/RxQQr9vptVcAWHp3GePKY+mO8g9EgN
jDj8mDVJnbrnEwTNsQINLimKhwIpw0Ge2TTw4p2Pew/4DqZ/9ysUhURiu12jaX43ySiVsfyw4YNx
V55XfOqS0X4ie/USEod+rbgfwuuknboGvNc+W+FjmkKxOLKKqB0Fhl0xPw5FWyDodaFMBYs0AoPR
dIxJBooaPKWQgjXatFJSKzjFwWzuspC36LAXCA11URejKwTSAsiYHNg1dqR8xeyvW5Sx0f165biJ
xZ0bGhay48TEE2odpvTv56bYZVNSH3hhZDMRzWKYhaURUMqhhwbhPo10RDzYYQ9tlvjSsmfmbm3z
aXLwzbCfTaXRCQW0IwBAYrX/aWmVGRmwr2iTTLkTgI3yFAy626yKvHBWrnwbjfIFwhtM+S5Fi47W
J7/idKJ1V/EQM/1J3Lwvt5emext0JmmigP8NKkQPJSALIXP58iJWbgdMl49Vk99m/bKSN+tF7qxb
bjOw9/+M7gvq42xRtQ1KlQ+h9tsbt3v9PG/d6La9WEi+vWP9sMdZnlmbcDDqyds0AEVMz3ixbKVY
Q+6TJrZZJmxUXfl0MI94VOBVEGU+M7E2BWS+yjZoxgBWU4Ibs6uQq6vMLZacAF7KIVPfvHrT5QpA
J88s+d60tKoXequWLFVKN4SlCyExJjk/roB0QrNQFnGNMmvtCdHvzjPJXz26YF3ggZ/cDd20SrRQ
48YUAiZHPW/8H3ydM2wRU0c3hpwhl9z4u9BDoXpxgxkK8EWH1lxQk1yXViWG+Tmz0KzuaAySmQHt
3YhQBunBahxAis0n/ia5670R2G1h5fAU1WzozQ4vGi/LLSQLPwd4MIRnx0T9BrOkYCzDOMWIrbNO
v5uOtpRyN51clpcC1nsFXOCzH5Wjx1acWptT1p4dAhIeMYAbwLWceiya7VdELbnkvCV0HELcexdn
tTtXrQ5Pu6OF8WRQITRb7PIwDaREaUui6JmCbcSU46Rvn82CXYrKPBr8mibv0PzBD7Ygm7Gvv+8Q
1imL6WXmQxro7tUrGLB3RV6iDL72fGTyNDgMOoT1hddAdkzSU5pG9r+1PkF0k5B7ej5A9VDqeakq
a5PlXmk60CJ3FhqDRXj1bMkgO4lN77/GOe55MOkS0eyMnLcG69uwQ8cKoEj+MK2Wmcsp2gdivOSo
jO3gbZhgxk33TUYb/SxKT54Rfgdgss7L4oWRDRuAtoSleLBu+BerNRQ/J7M8FaUa8h8bvfgxv+Pf
8/pLdI1hNQUMGEVHt/+35bRHwnJfNMljk68bckTx/vUJhQEUKaIk1ZmDkoyN7yNS6t6V1iulbpEw
1F7J7IR3YkRl+vY1o1kK4x6lrsvqZM/s2D8P2ya1GXhLCUFmAKR4y8ayIR0fSCgH8vOw1ZFB0s6k
c7xxpL6rBqq7L8ajgMD6r2s/aCBESU40dpM2hg+GExUICD1lkPscnvtGw88tHhMeHAewNC2PanFT
pnDsSyNuqeIKOu4LVkz5R/9mk7ghh3tYJjVW3vt2uSl8PW4uR9pT6M3Ys69fmjOJweUUzQhtHSdI
3W4tLqXEUGq7VI8djhs0L7Xwx9UVgexEz6UN3ZlMofFCFBiCwlWWC/E1R/4nkR0MgHH2/b0x4/VR
N1dl6WDhW2/ypykRK5ujSFmjczlRfObdYG9Xm6OMb7/cRnLH/F0JeFzYBG/siDMfiDtFxq0mi+9J
gprQ09vTIMYCSRjT5wOvtxkTtprrHGgpibZVBm1md61DneqmNfhtu7vfuIRmUOhzk180T+Memiwl
SHz+4/PijIJNjIf08IqeB5XvXVAOiQ0vTJXLs21ooG/oRuCbvvkab4yJ1AksGr7mMSo1Y6FBUNbB
bYNmbStY+9VEIeGuh2s5myIC2txoAvR9YpT4x9O0P8jSlK76Wzor4djM1HRVht/uNp7d1kM5eP23
jC1IuHlc4BkDBM+QAEiEAHMdGw/98Tq8ep7TGUr954zMWLjmkyrqDOeHVZBDknTsP8PYpIQjgD8n
vowsbTe/dj3t1Ziu490ew1ZFwaSs6Rg3CVOZT0aLK+AbdjeSAsnRLLzrmecAu4XumPa6m3wwsymm
m5TmZ+sxRP+P+lYlrLTvQj2KKitJO2r8l9gJ+sI0m6KlXn8Dg4ExDadO3jAXQMeavUdxrKKf04cQ
xtGQOd/F+ofGG3dgdcfmVv+tCrSekEpKRNB0J9iQlNthK4nPm9lnBpSYB8mMuxRVFQDqjw2nmq78
LhK6weE5fMmTtd84saBTgI4DvU2/8d7Cbe3D7bT6mktcpAOpi6mJKWZ8rG40c/bqLh+sZ75A3Suc
OkNCCeVpdAlpLIBKGkoMW046S+Ml9k7gRDy8RHKc7VZyZNlnVRcqxLXMPKnwN8MI06uDM2DtQTHp
b+vN5kc0W2UIo8IRj9B0dhdEtf6uyrisPZj/+Z0CDtkJkbEoYHS3x3RhWwp3nxV8L72B13wGdkL4
BXDUJj3smYlDHkkGDbHkDVFJxFBAmq9MB5+1JdBw92wGHCyaMDvmIbunSrIhdaQ8ZEj66QxljifG
qGUxUbFHEt8Cvo7qo2w/mSxPXAz4TgDPXketKpDY98E7nPfl4gq6Qi45pAupl06xBQUDDBZfwzwX
wq3PPpK4Yvpxm/NIz3W1RXRT1/lo1TGhzW/J9S9Gpr/AC9hI4hr0yXQERaKGPWI4JykWPPTqNd3V
v4K9okfN2gV/rxVwrQSEbBdrtgUvsq7T8aJ5rYaWk5tnPTpTGhxWPRqSthRsctOuWpfEBCLFvSYU
B9lzaezFUssD94V7vmbI0DXjsZAhlXMFDI7jBF4sH9K/7cGeeR2ZDQD/v9ZkJIw6aL4eC/7HHA0f
ObhEuWVZblejjRFylyJAqrm6qOhM5Tehd0ZlBo6CLcuIxH/s4a6orXM2J+5++4k66ly/ttAPIW19
mUwRvWSayCjVjetjOKOUM3RsfDhpvrB3GnTBGmoWVbgFQv2eVqErY24fp08nqIZZ1vvjxuaJ6fsB
rg1e3Wdz0FXCTAgQbYZV4G1WOfdJTPou47PbBsZqL7Sm943A+aRa7VWrHAX3rm1/J2d9iJMM8/z2
0STCiKoWePWicHaQ4cm60aygvahGB19gIWUDWAEDIEDkzhaP0+wOVixcN6q2voe1aa25ugvxl/U2
ezxkE/xkOhcPJrPs/HTY9QxP2hPSmPGGQ1u+OXkNCRe7jwoTEiTsEfLsruj4yxbMLCYjurP22ddM
XktHQ5pviyMeIbxF8tNaFo+eTe+jikOa2QVKtaPQ1zgurUzjQDxw2+2AqIzr+Jqrzd01o4UMJOdN
fJ5j5p4ZwaB17YZTD1FZP3optOA45XTagqpTgviS85SZEoZ9bAti/LO2xq/mbkOo3HDwHJkZ08iy
itjcr48PDZboPYFnubnkALi5bOMcWyUUQUyZ2XFTSzvy/MeHNO99+Hk0LGw2oBembd/TEcj3QXz0
Vld0gp4xo8z4W7RyKnvb8+KP3BDNXZpke/hn4Ytc2IoVRSa+FK+OogQDKp3s+fRF04rnuqjWh77n
g0S/zBCQkxiZpRC2h07fexyzvVFomtncXyK4yPXKlcnDqwa0co3txKWTPqLD+KnhqHzoJk4XPC3A
W2k9hR3oGcJ7suNhLXjUc/h4w62h8IJkFbKD64ExT98qVREkAbhoeHSgODmYpQIZfdVo6ctS5PvQ
QvkfgrwZAwMVzqaZUbOr/2fo/POjYacr8ISd++nzzSpkevj+l/gjw/vW0hky9W/jzcOpINb+gv+T
cO5g78qFTg5to4ptijLbOv9mDJDritEGNJVEePYAa9YgCNSsuLrvhTjw8iV7dk55/dQ4saAkJ7r6
AI+6S1F6URscFgixT8+Oi6TwdlImuoSJy1pEN6J/gpI3ZLSJPyalezmsYIefevE6GKQ69twTq/6y
ylj+1FRS3FfD/OfbgoW/7ubOr+OfxdEHyq8vFQYuozmP4pDQDlreQ3xDMhDzfgcN7ls70LE/Z6Jx
D/doMwNhFRUTUUSHp2LhYiBDwjyLG4zyLjELFYtI5vv7KKTaobHEJdzTyC6tx5a8PZYAN4j3loHS
ORhNv+CbkcEG3/dpetI1bMpaU0TNUxiT3/V8wb5wjcsnDeYd3sdI8j7a0YZWq9TN2pcRq1Nk/D81
V8dsCqIrEC/r/C6hBjAD+uBI5WYq0GNRmftaoOWiHXDffRPzfs8qqZYsoWioPgOWnY11c//xP64f
N49iUtKm5Z00Y11aNjbAvVm8gfj/80R2TqMQ3fATcunTJFEscU+a1dGy/ix/JXcdOqXcXTZUfFKY
5B3+yXzkAdjEVVPexY4bi0kkkG7rwqs9aULk7MkEO9hoNq7XnQojadHsj/sz8L/RpvSrjMwHk/s6
3AxGZ4s5ABb79+rnxgEVNQblKnceEXMhy1LPyBD9NGXAz1UTIST1yC1wZ0Ps10SZR+lzsWRk2jB5
y1gLEvfzKNbVXlEf0xvH4jeOTwy+TbhA7BiwD4HPj/gguBmnaEpFfOzxz84WdhY/jYgbqPwvIv0k
eAgoFqzn21dT0cVFSXXP2UTGC3P7wnrlnLF7fuA3GgDrA6WxVRne1lSFkfcSnWI9smclyfCDMByy
qzCdDpsFr3NmvoEpCIbE7u6dry7b20jcY+dxSqdV5duf/Bm74EoMtogrZqcegoYCFyA5wKJ2GhIT
9HxRoyG/XNN7F6gW9vg89XsRhIDQ4hbcqOJ66HL6WCeFlEcvxcNrrue/F7rgOyteVop+yx1Lvzdn
vH8bagfKdvmNaaeOMf/XhaFVD5WC6TNcCD7DwVLAlD3NEAN8ijRLA7dCnmP+J+jcHYSObxcdtC7d
A+FeE2NI+2nLuoKCiGb1aD2Ai6sloqSVf5FFBtFWViNGx2/IFutwhMHHXi/sC/9uqWabBs5wkunS
t7DQdEzBT9IZNeIJG2jD3tXtrLtDPoavXkBXryzl4BztBETgxTbreGFKkJ7Pj682Al1XWGsHcXi0
Ep8bE7wHLNG783QfCsZCBQApPYTEg9eJdyFczfRCPogqJ5Sup8rUUZvpzYrL0bWCsO9p8vffmoUs
5e7pHz4RKaVnB3JvEsBxp+7MGM4giLUAiiPTyAmG5MXi2YlAA9uPePq4Wz5T4Qb/SH3cT8LxrjL/
bOWvoYrb6IQV+wAiQb3n4rsrVFGhgYuqYycaUwLBC2BU/4ZuTUO4PR3G1skYkgETNnMt+L9vhG7M
G5s+q+ikIdhbTfvsew5Pcsvme1YwnXdjgQL252oPmfd8nCXo0drTp/6+8Lq5B7HGBTz06mI6DPOD
jDBr9ovRLP0ymFyl97HnFC3vulBd0FrAhSrfNXzgG59U29rK/7mYiYQkuSr5zNMSxhNpPuyDgEIw
N828jsoxNAebY1zTb0hhUNyH7C3138rPsboq0f6+pghh+wBbMf68y/wTWPtZX8QJR8jU0h5zOHPy
1IsgIw1A+xHU966P5/sdS1De2NHdiDPWYynL/IvS6+Im6jX3BhrDqZhXl5fMrSVHYuIn+fJxGxh3
sN7riG/DiCn3ZJ6VNsAQFWYQ1LqjGAnT4VKRt52h3GHwhRh24A0zoMkQpuusVae1Zk8Whfh9HIvx
tmqZeFn2C+V3aTAiVzpT5+YqF84/4N/NYPi8RaItBH7x+HAbLlKIhOQV8OI3h7ezRj3OZNclsHeW
Pqu7fIxxzZFXMQGZrxRDiaW8MYtoiksvK0JtfQh0VkPlFxReJVH6fpA2AwJazfo3tYWN8CRMSIYU
dharjnRq5WurZD/0gO2zeFIIPzmULKLb7xIfzdaFuyXHkkPZhjMSFcXknXYBZqjNNGYXDW7Qhzf0
iWyZvHLOQBmmhz0pNvmkr7MCKo5hQaB3SrsQCQ1Grm/LMhKrKTkK8g1FqH8CW4WSYcKhv5xkfV47
FG4751ap26FU/trsdy79rMI2qRIMRB+5gPHkB9RjVf3gz7K0eTq56CwGc7uVgKyU1UYhRhh77yfr
JFUKizmTmb49iARIUFABtvximRLIys2+wCZxAOilHglD4ctfod/MlyUhvui7zqe15C6g8Mxuos3H
bFinOPuVpojl1K7cTsZyXfwcQZDyHmwdxf0OsAJzMQ/2tloU1IRp6aFn8PzUgZpEd8eVUsFaZ2DN
Kg+g9hJ+E79OLeaTEen2gN8K09W2mCFQT7uwpMDA4OygXEhQiP6utLrbP8TvB41p4YTtmL06GI8U
PH9ggfKg3yrgXDlc7daTAcEkN8BwNjp86qrZteodbtzKPDMZZr3fyPyPZhQzMiaek90xC/D5NsoN
I8FVCUyp+R0LoEf5iLJ7O9or4U8Oumub5TAMz1jWVTUYlkBA7tE5tiOECILnFwE4wsn+3nqpdFK8
swu6rWn7mqmmTOshE7leu/rT5ILCwMWLeJr8bIXkXYIiigaQrR888MUXekx2KI3E7db+KJiUKd1m
cTBp/RSF1gr2Aw9WK596KZuEmTmFDgdyWyooBM6BPTBe3NnBOz2mXVs5SlOft4qEF/k53paK77QR
qOrv14joYa2c0LBsU1NeusMJXsDCpLjfRX+0RHipITPiOpCrMrR5FLotCGaeLNNjuiNGh7v9wcr4
d73QOoUhePoxv/oZ+By1Gc5IxraVPsR63K2My3oPiMF0zLL1tzY4T9GOoyLlslXalSj6Cnmwjui2
ONyYXnAP/vK+tWKHcTwGSo+VqOI3YdlKbwClNrtAvwY3lxv6fh4sbNKc8blBW2pgt5tp+ZvgmEm6
iKFwFq9UrYEksDS3Bh6Yo7+grJrEyG7PxM2pJEbSSQnDjrdP/sF47TtdFqB8dZTjV8xrDL7QBaLY
1WpHaM+jPgSGP9+JX1TXh5mEtf/4Rdlua43Zrx/cwTOSPFF6epmjYWM/51ng4OZ+RCjz+lguUtzT
NMKK48pjgKOZr7IT6Tg5fTN2QOYm+rM9+6ouYXZDK7OI6Wr0G+/HqYXxAK+H2uedq6myOdfQ24dT
P1s9tc6C762l0zVgmbxfMZk9Vhi8tIT8dmWpLIXDZ29o7giCXiQ3+qjH5IqN3gQm4S0J3tTH7prE
+6L/xc1poGqiJeWi66XUVs7beu0OrT+yjxj/RQAzOaK7mF1wRGZguy+WBL1LtEMDmkZ3qzFzfj/d
KfdYOgCSwl6OqTwcvyhgNWgwB+7fKMjvWcO4Si578uD7I5GaBHXFAMzb3Rr8Alst/yfhVJrGwlbI
87FSw/02DPO0Xz6BgEo5zuj5N3NyZnHvXMAHY/4T/I9yKw7DXdFb7HB5DSAASUTmOALJybqeJWnU
Ca1iRVPc7TmuEyMtPuSp1uEJj1CuLzpvWQ39Tp0pN2aiSkOfuBeN4e97quzWGfQlvZSmz2ZckQhg
S3va1l6ebfMvWKglgkujNzDoskeuFS5WKszKhLtsXOKjxMDijSHb+7CcwxkiMh8ESIm/6huX6WR9
hnNw+saD9SR3wx4WIshnH4I/A1x/K1K/WxLgoW9upbmmGX+/Tp42P9KtFwGU7GpKTAg4fvj4+9sC
jQAe5oyXnQS9FmAuj9+NZ8aW+xUv0Q2PSwKJgpVRfNrUhtkOy9pW6Lyf4Byd5BGF0+waFJfG9Yxb
PNy5WbrOdiaEKA2wpwLYq9032SSbugWLFEeUpU/QrJD44oYBZt3Pkz/WV5FMgRwQ5D2ivRrEQ9VR
lnLNYkQfQA3euVQaXNsZAzyyg6P3jVyyqpg3mc7qg1WkkYvVYN8E4ZGvvLQSBP+iMdEZbidRxS4a
5O74dpgL8VfTH2xoLImXkpKqrhOqwTw/kTDlLplpbxiHGJOkTMXfAljvqXZwPIBah61BbDM7mDUw
WNbfI5Y28tuW5g/lBa5Cyn3RF7Q4xx8S0+dadJTn1nNeWjhmSSQYFoMMyeAjUVoFJhW2FQzlZIHB
nNRWFbsKgwcy/LLXCP8/K6/95Jyq2fyqdXLRuqckM/nFju8L8FHcjerQ4F+GTyyHD06+xuSBmesw
NLbtjz3pfgLG9dAMLiI8kvJ5NdwP4Z/iFmfTcMvntp29OpKLH0HuV8VmZb7gQA1pEMnTRLDFm3MO
3eBWoNXKOFgcmutzgnMx9ZykXma3IZAwu0Qhpb1PU5l96/5jP2WDW7FKL+ZdEvJ2rQBoWYsQFq66
dDXmEfY1vgA+xX8QhX7HV/jR4LAy15fJDMmxB4dp0M2rFZz4NfYi9lr6tbuje4Bn9ya1xFQFWhw9
5oTvAZ38c+6EVHNqhW+3uT4+YXmaCIhnGc9SoiX4CuL67+t0mMAcF4Fg/9j5F3oAs+lOGRVYxvVG
AtaVt0Fo6fvheCjsWBmN1u6C72LsNBxw2z5s8LmBWr6DIaMw+8QdAWeAiW3FDlbW1Fj7AqKg/lsF
fWGEaQfgI7ll9nKGUQ+6yZnTTlfFKDjf4SHuEPZhN+0T5R9nAKEdPBHxWAzEfsspZFtSj77wVjH+
xJKJhDM6d6pkD3VzRC0jyPHyCXXGWFkXb4e20Yp8Vz4fHYt+aX3CJaScQYCHct5UVB9PD4ANrUH1
pGhoxjp+IBk2UwgV+YTmd98Coh2vVPIUu8jwcaMwbkP/y4kjO7eDAKUYhw8CBMy6Hm/KyPnSycfE
VGKLvQ2h00isoHJ04YCJMacQI7PAp5thNuP2021xresFhW+1OfN2smMbnSOmyr3By9qNiMR85IBd
PIKAnYbbLJ7E2a9BhGI02cnqlEf3UW75cf+Uwp68IsEXfBB8FLUKfjh2ZIEBdpvgZyJClKhHkcEj
l8kYxx0J3Hwlj01W49K2kK+Oi30CEszAxZi1X8hhI0o/zOUU+7eBgFr8MDZu7CwzCb7RoCxeWNKp
5tnV4LCvsqxAzRXkl+0kxxeeDFD5k3gpQjkvFUDb4Mlj7WDTDfbIDCugVC7a+/9Vm/S7r+ekXFDp
QXg3aMCnMjf1n2JEWT8muj8Hu1cW0thR7gJFU6HUUqQ3h/P0SnKpCheVFMK/7hLV+dEXhRnfWYmi
mWv2CkSScCOdChTiNFhPt2sEDZOzpARm+pilb7Vt2XZIEIEyUDtiGIyneEwo7obw1wTT4GBYqIQ9
h6v+WT0Xrde0EpEFLRfFWr8MtPku20Ipo5I/Cl5/KJVkgp5VyEXZHrNsw0kHBNmzWcev6d6E9pb7
1JdxWeshM/nfbGF7HX02dBjG4AoKJrAO18HXo0589xhtL6s4oEBlwBsGF5gbL2Yj8LRfEhuAMr9r
PTrdGO3u+kkbKpfulFFGCP7L48kSI1zQtovmDy8dr+rqdG6oRyJCK1dCapJwFp+O6FGt2pdM/6BD
jgpH2EU4CPIfxsWNJ0o1Rx9zHWeDPVAPXNBL+V/HXOwQADNXZ9yQtSI4Rl2/xQlDDP8fr2U5nKzM
Od5U1SlwI8ToB37+1ewGCp3HGlkXn/lzThsGc5FWJWj3l7f6ABt5qN1cJ2tTxSfCi58l3m7M6dVe
EtlYyxNdaDymjbu5rOqMiFqFS46c3QgzGGALegDvaec5yVohL47KbZBLGn36zA5LRtgkVI+uXlSv
Vpy06wcSbQGsnwl+sPJRZuTA+egFQ9LP9HpYHhLTSxavZKpCVUL6X1eR+rV/Oc8RV2EvbQpGyqJu
usnA+esAeENK11dM15xOOMsXKc3eE+IHGWibKlSS15uSlYWqACrmy02WTA4ONriseeDhVsvsxw3L
8Qw+0sO2IXJf4lv2dZR1fVKtEfbT5E4LM+CivvPsuZ7azHSboSdijkjuxdn/Uqthcjbm863nCY0o
eDkctWW4S6+iSN2z9tTwUOlBw21PZjohyVREShbFd6SrgxSiv88VpXyyaPsqx0svT7q/rVx8/CcF
yBZd1UzvcV6OzroZpBbUIRGivodAclAmlnCKT/cc1INlbppWuAlqctvGUt2w9Ny0YeV85HPP0XOY
bnYvMoe3hd71wkvx57SVR410YSO6FldMQlu1hSFXWVaTK0XJAM76jaKkq2/fGnweBc0nPcZviDm1
qtMNpEZzPTT/u1Q2ct4qAT630tjVW6Tbak9+ikECO4x4gKrX2AcHSXArRlpEItWSL7U9hJa+yczV
b4n5ZI52ZmZSwcnmWRVHRnkoVZviLxzTAikTzWSRm6RNhu37lUa9bjLDiyi/Hhb4P0ZhQ7kkhZAL
e8g+7/JnDbwjTy/Pjj5TCYBa5QKNiU3frel/Sm8sCEVgdADeoZfYsy0reYPfS7MXIVC0AVugJ58z
e5s2hotWoHyefCQmsFKbI+IhWDGuKxLlAvVDmepwGC/VYyjWt3OqO/a7ZrwZ4E38t8p9l2aw6sXz
w5WeZK3hdaX6kvi3wnZFPHk/BlX7VsJXVKm+jsnrSTdF+uzddJdTGJ3jMDWfWgOeOmyVLy3BvyEu
oy+QFp/2pX2FTq5j5xRdFvyo+quu7y2HGL70Ni73NKZ6tILR76dqxoNiSR4osFoG2kTdKsmQ6p27
Erp1zhsVChJhMKgcm/ZwGgFkaqXjSNFPKPHwPm1ZsTsy+cl8H5TzpOeKAjQcq+uZvrGwdOtBSdTY
1IHPGYqqI8AfN7tuZnKRJXqb1QAEoiL2vvisPwfqdv7pZ4O8ZwjLZsP09uPOWUU+QY6PpfVY2q4D
VyTGLQ51n7AY6wqKo95rFfSUV06//mezWiG5q0zDwW86yJYgZV+6ZxGPU56S49FMfMCiqA9vzl5O
YotbiWWJcojdp2SM9UwxJAOjN4QUESm6ln06b6GulreIqYmL/K2rgJQqbs2roybWA4uahsFm8sTE
ZYrstf8Xh6X5jJrArnssv8ZYpd5pI8SkqGrd6WUtosX46DmTNAFv5y+ItgKyfwo+TcDQEyGKk9Y4
jR23NhkKPVazDqO7TQRJ1gaGNov9O8nPm6Tt+lgMXChu4jwaqOYJnHrD0eGG/rGtsvKadm4DvcdK
WsnLig3ZV8sm9qrJYnczXJGTubxVMvURj3A6kJ4GiB24xx8b1MdliapMF/XFN6L1mGGWj2ao3HEU
6vCf9q+Omie5uszSsW3DTu/Fnbry6opQ3QR1h17LXclGmCOPRbRfwAK8R3cQwkTwcfBJcXjXlwA3
/6zZp3AG3uCMm16r6c/QFQueyfRfkyIPYyfKdwvWhhbOyYOZKHrA0sIMVsxTwGNK2CmdatMOjyni
u836CGifzy225vqzkTE7nvDnQTT8i2WvXieMiCv5T718TYoQi7MHv7qdkfCwV5jxxS60X1UglGyZ
/YeiqN8GPLmw6hX/LLHAXafPAQsRG00wOBjHJRtYjYWz1N5ppuv/Vp9RDwhWZy7aQKjstoO6yMHP
4TpW8kDITync4FkNPoitMeQZ7Uzm8uY8KKOB+ULiwOgqhr9be7NxjFw661jN8hPVnDnsZgWhQixb
IJ9stcqXXnjELlWAGD7RiCxWkI6eZnSMBQ/jzh2YklObnaZKh106H/XpIeBLoIJ9oNfaX0c5g35e
I2omr7WAln6ZENampqR87+QJr3PcVnJjZneaD3KdB4eUd1FuHiq531/Pav77ZCKdzjuY4LCdMFoW
3fERLz4v5S8j4wyJXnyQqLurX+Zbh0ADg0Et8UflXEnlJU6mro9EOBrwoMIYQH7kInOQhlgc2m1i
x9aHOEKHyDJyEvhJP7n2mmsNR9cv4sSdn01nLUCRVIOTu44qZQ9w88bp3RBuwd1vztGM3rxSL+Z/
WsNGfoIVFxYsRCaEMu0TT03EtxqzoSFQJKGg2KGi0ufO9eYVsjOzIHxgxpuJYbbk9m/Y2uLc6oHx
4j5yhKWPYXxv0amAuQ+6AJebn9x7q4s0lay9+Vqeu7dKj9lKkFhtwiQI3isE5ggSYRe22OytBOfa
nSdUI6WvnBYtKtpIROx8Smxq7ZDUVbek3hUDSxCscr3rPHqlSPF+I2NKp+dQ0+V9Pb9RZdoQkPdI
P8aZ64sDDSJa0nRfv5+nnwxEqIWREdCRPEXk7b5TOu22g+QdM6tZwOb+t1PONq5lAxzZP1ymY1Cl
EC45kVmNiq6cp7Bj0LSYoMR9bI/pZUbnu2kc3PVran/jlmhYc3YPRucjD2aHc7fhoqPookU5GzQJ
frdZ6O+mlRebK8f+VDPO3WSRiatuWRkrq93X8b7LGZZdOQE8pEkMyJBBqNpxbjoWAd/VTgA1Iv6b
ioJVH9sDl9AwfQ0fITczGuoj9j4mUo+uIkZjSgeFH7fSmKBud78VbF9OCloeuqHSLTYGJPeMRfya
Sq2gBRvl0dePWB+7lYmbBZkRaHxDJjV2J+vqmflCNQA1WQj7YobV649eR7uuUeqkfcGfmUrg/CKN
IBUUp6vv1Eh+lATcJZqJx8OslF0S+dUqZOWItEbtEyxY72gVto5ehVkEdG6Lj8XSCGJjBMoFVwhK
OnvI3d4utCksoClQj7cNSJhoHa33dYYFNQKjFM/aBBJSp58f41Coabwz+AN1y6q5Wv6PoOgSo/b9
0F5dlNaGfIu4sK95lDw3RtLdnlYscNWFVX+Z1sDAbOQpM1NnGpy+CqD2NpU5VElJb0UEDgn+cNqD
n6b9T6u967dwQg18Oq7MH+9ZtLWKUC8mwI9ksYMl0G/HBiWn98z9jYvgE2UlF3Ec0CSsuOmSzmRH
8L+NW9NM8R8t2cAks1I1RMsPQB+m+GBHdiyB0jkZCdnTvZNDXUgcII+HuvJL3USjlDmmrnhS8dVA
hFuoCZrnGN1O+sMlVGOSPnxM4um+Eaoyy0w/ldoJiRt0nWF1iwxB2izYpEoXL2QSDxaypKy7/W56
zgUJ4yYNI9bIz4ovgbCdv1Mpzs9QZZK38ska8YiuP4tFapaUE18xBD1qkN/4QmoZbuh4pO1IWMY9
G4kESw29qRtmUEdejoeRNDugteehpGlqYr2PdAC6Lifn7CZqeZ5wCJGMHFzBTLTE2GDo5AUeezKH
VzEjbVd7UQ8KU3k7axFsy63NWji/E4SxzrRwph7tTQs+hdmzHw5TebDQzdOO8fGZ0pwd2n1mUAf5
8K2Zhm7iwiewkFztHie/oc2cJjcR3QB69VcjlFj0lEM7nr55DWTjb6+d2WMAxcf9PffvhXzRmCrf
5RY5qESVIgxHEBTMvFPdhQpDu0r8nJb9D/qpRQ44lrMMLRVXUItHOEuLk+6jmKpL6F7+OLO3TmUn
QvgaSJ2z9V1+aw4RdF+81L18JX1t/k84pePuxBjg5fGupxvz75fYq73LT2LbVAAy9R2R3AeF1G9a
5MkEYCGr4IeWLZ3hsKA0QAZqwZcK/crqWwVI1eFyhbmZKw8kFsJdminlyFLJMYZ07pnDFV8neDRV
TsjyP359DjwUJaMDtfbgiKHbQaA2C+8aVt7MJmFrVWL3LAHUF4EJzZPsab3tVucl/OK4ZgkQ6ngj
QlgxfBDo4X+swVDOLoGVQWxoyv/f2nDKRI44PL4TZpka6Dkn5z7P4fbVVcI5M1N1RxdJN/42xj2b
P3js2SMJZcBIbRiIsT7lU7xAsD6zlO4uwI0Tz1w7VrAZ5mZqB/YjFWqBbAT//TWvA2HYLi63awVe
/8/teZeFf/Ewql/7n2LXlopbjivx+z060hIVpMWT4jC6bxClJcE/XWLS8zCTS1BEPrsxlG0hOmfD
/IxWPkNEUkXiosE9JRnrKZOTDCK6zS3jc+iQ58GSIIAbe+swNsvKdivaJmhp1mRoIFghacXiPgnw
v/ry/fIvgAWs6Xcq+PjYHZy0K5VVdBW7cRPlcI5+yJqfybL4CubuHCuRKplXDD0kInC7J2QA2epM
/32wS648G2rIB5ITdH/UIA6QLUWgt5GF/UOw84/9Qqi1y+fkbhe2Ny4+jdyghrbn8qub6SeW1ZKD
xuQThodGRswfhUxQ7TxjUDAmfkqRbE24SWiX5rkuNXpYp7GC1/BPgnAich+azEtt+PIx8z+cwqhv
ByADMnl81MUnjq8KtUWvKiWXec67BlPLVePReeu/xU80J5MHJJN0G/IPpexiLXz41j3LoxMUFDPc
4H2tgrutPLaBMr1qX6otV0LWe6ikxf/oIyVorU+I0KtSPovE/KkSwssO9+qhzUEj9sAT1b4mXKvs
WEKsZok3k9o4i9AZCHTryNVZ4hr0s8ylY0josHrP9N3Ywosd4/sf5+xm9yOnB5AADCH7JSiy/iw+
9y5lOBY1GKFSr8z+8ECShrjYbKRB/bbUXhaVKbrRdZf6lcA2dlN1CV5z0PPEIsS7o1P+aHiEYkqV
wZ+e4iHQZsiSpVINVB4T+mZv43dxJ1Hr/EJa8bXlMlb2EcObO6hXFismRd+sYmhurclOWDvZJ8q3
NPoOW2rLD09Y/vi8Kqe+2w4oxLdQ+IFnnJy2Iz9t+yaN19kVUc4uw3z8PDYAotXeoMbRaTBWvT9U
Zok+7egP+hd+QJNf/mf97c9Qp8x63CUX2IJdom0ZcBS5H1bcgvDVlN4MIkB6X2o6uvXwv+q42bFY
RkXk5tC9YFmhVvlAf2l7UbRIg29uGVUPzK7wCSBtWsEsMDMvxgY99WX9iwhUVnH35zPFY5tgs167
NbScCnzHXkRFHszimvGtcS1dgSKBm+q7LYeJAP4o4ytHRAya4FpNDTsZENq3Y4hI4uKQPOODow81
DfRDtg5F6LPXP5hymlPtP9NWR/s0Al6Bruy4QX3X+zsZN8EeeTDWhSJYQF+uY42ipWgye68mtTOc
6jhEj/G+OThqxfhw97BgkJ9zLIoH5fmreGzVq9fdhgfhSLuBpp3FAmosqheioJdCFGzs6gNVyZTg
OZg5X5iAzDAnqBG4oKnpiyZCMNjVqwXKch8s6/DPuQvjymgFOAi1Ha7l2FtL1QEgmlV5XXXva1y6
wXx+2ITdZggcf+uRjBy1LSEHmkQm5cymGlYzA4KTzO6vGrSRlqF1MlJcb6gtPyvxQ3+YoxTW7nyl
U58vfPh8DDxOYmfcVPnGRWG+aASAkAanHrm9u68LrkjaQqQIlEQynTIQHRlLCQU0kAbgKGN27g+h
aN/5CWMFEecqTcn6TmouY6iGAVv1ysJ+JfQoakQA2M6e+S2GWfD9miklCxMwaOUdx/5kwHK+BUF0
fv60gnrwadYt5CqiuEAMbv6WVBhpv7iFekQ0p9rorTUONgbmWHIkHDy9Fr1gr/JDBLF9IH0ubwQ/
yJLeu/YLxinVjD6JX5xgph1S4XNrRTEFXDvr2mF5/1LiCCP7J5jfjiR5veLmmQgOSYiw7oFL7CBk
4c2yz7OH/pyaCL3sfFXXKpomhevFU02Tq++qpGBkmMpoaBoYnbaeKZxpTX3G1YqE4+yFrbFWxwqc
VRz5zNryHv83HtOB5pO1guPV1yIJewIkUSH/ZMZI7iI3cGofjQ0IQQpsblcaxxN+4gSizHiqWSfB
/o021oyz16iPy+lGjc/Wp9mtrKbaNFinxbqJ6uJ+27GKxQIc0lg4mMdkjAECdAnvwUXlomJoIfDs
tjtxcmy3wd7AEycI0gHs1dTWNd2dsyrFaz9fpaaYy+gcAAJyZmFh5Ur3WCBQRgoxzz5Lutdx2Vso
ve7iADT1M5yrJ1gDU/8wetduvjkHfgE3myhBbs/6IIUuc3g20jbOwacovH4ptjE59ab8Q9/DV+H7
ZJwcBXH845S4kguwm9rAuv1LAqPsLSNgi3uX/DHOu8Uae57+3NdWU/cyxjVEA0Beu2QLzmHuUu1H
6YLMChYNxpmbOZ3xTocIbaJhNwXZgopqX8Cjr9UkgMKxj+7bCK7hkU88IRw7LcjkFTtAj4tfCii8
lMxnnUonqGQ8IXKgBr2EDUMpFf6UEevuKx4V3F2fD1YQ5omsW2k2blkubrOhyW25/NuV5eKukg8E
zVJAyYTv84s/Q6S7B44LYVhV19Wl+Ba/vg0vKkin25vyTzykjb6CiGhcBfjKRcdXrGHhCsa8xEos
25EQosj1MFXF1hJ7vJL49QWqmuaDlN0ebPumhqe9RnOIeRAqBHik1hde6J8KXrcIjbEXcA2Bxmn+
YVADIi+J7a7LFZTT0ObdJLLZXgr3ti0MnAeZgX4oIWItwRN4QpoUrrvwJUGK4F80H+6kqBB87E6F
EC3+9NKoyOWkwA5JgjuDEw2u+d7w3PESDH1JgVc4Q0r3RJ9rzVkAm8RzkWOT+eIKTiaXtEBNzs1W
O+lZoIdo5ll/fAhnJxMKv+gKr3FdFAMML1Y538tMByshOsQXFsLsSsBKFUvaMn7qb41fBOuChEAS
UEMrBBSCeNfGSufqqD3pVlFL9elu8FhkN4xYcUqMB18uhPacERMEqU1W7bJdQAJ1EkCtDL31LRwE
L642nEJRE14mir7/PijqJEPPClK0hwGAsxYXQlWotLTIv1HMa6g2MvNp9/baVDFXhXaNEnw24tIN
LpCpNBtFLKtXS3s9iHsoEQ3w6o03AA8uHMXv7aXRe3fr+hgVuEsP2s7OGyHfiZqjln0Rm8RdDFEF
sqoxE1WXQtEQVN0Wk0D1f81MwcIY2kMV3JlN2jXuZldCh4hPED3NsRb0IpXbc3NJ91lG0fsFLYFm
mZw/xIpA+35VFE/1iVRgpvpD5FQoPBoXuP7PJgiOygN75MBs+nfruvAOi19tKuzYXKpc5JaXAdZ3
Ti5EKwtLxwmoTmP8zf/3GDJHez8t0zgI2jxJgrCOh72UaiEC632Ghq6ukDtadXJWAVMMU11bTGdv
/4gecazcd7zFlLB3Z5YcU6X3ix77l75lJipVUIhh1eFSKkfAJQ/XAhpXxg+uEaZq5bLj+F15TKeG
hnGGJJt+t0I4JzWfXxHSqJj9lrsFsGXBCJvjTxl9pM6x06lg4GhoWXSKOa5StidOJ4zRSb2vF4RH
0s5qNkDKWNv7VXl3CRo6Cp8LcFsZXHIThla2ZeV+hA5lJoJDluT1+AsnZDC1ElF0LDISVzH1Li0P
I2kSOCApHsQXcP/fu0Qb6rSQ4OJk5vn/svWA5jzUtTXD1NyFN9IiTF83/J6IfG3es1bRsCJIEvf6
gKFVEXp3Z0smaqIMPI9jG144jo8q60GWoyF3JMn5NGtYBhlwUFMG7QTMNlmPpXj+3wnkxDH5OW15
bEg3sSpfjh2zfVK/RAmMvkrtf1fbqWTkZq1zD+/mWIXcIW7Bo2q+jxkOyhFqJGLOReLwDksYIOfp
gDnaN+KyC6tMTBE6DcCI5lgGI/DWW/NV7sNus9LtYHEBjDLb0alNnuTf320R2baTDLi0T5wH9C8a
P6FFwJW7pdr/DORy3mt9f9SrsJ329BuRCqmFn5meRoYE+xQAjH8J5yZHcpXViE3CO1VQ/ffJI7lc
ZhJZp1UZJi+yVE5wXn7m6YrQkrlHaHFNsfZ72BZhSdHoBdDsNjjc1EBXDU8laWSn5VYv/hAdabu8
YV/a1uWAvIsjMDFVE4yOE7H6R4g7Nc2QAnrxFIoKp3MumZrq5vCaD1mWF3QDwAbkn6Krh1gxcJDH
1UNBzAnbzOqZraVLWIbig6AavS0YQk4nHz7pI9RV3t9DRA9AoQCzSbv1kHaL7bcyRjihcnNXp4tK
n+esqdIBZNC8CrcTO8F5clOzHkfU+UBJbL0IW7xP8iSqrKckCBlzWNuvzN9J9EyuH00jzcGeoeUf
UG+SVlyfKP6/NSJ2JE0UoA888/VbY0mOhtBM6UIkX93LacPrgR8pDM+OowIBSlbkZr0EakJ0mZkJ
TszNAwAM7eyhlfCdhn1ilpv+RB0vPD93fVBCAcB/HcAcMYuIcWbQeeanlPd/EdrhZvButpqVzScE
VqSNgc7o4+UYaEq9T0ezd2FChvRmIBfh5si/jR5aVyJR651XbM0xYCLqbmuU1E5spEkq7JNAdj1i
DABUzuNYUvGLOO2+vdav9cBIt/MRJEPaB770A4yRQck7CNsUItSbBcwyWkCIWaDXTEwKtjhiGD0r
Ac3p8CJXTHhevh5daR22de/UmrhPuGw71slNn8m2v31ar3B2T9F8vKU0lfgSzBOtg2jgEeQqL6Om
v4qK5QSvMDLXX38/hIyVsGvXjqlEMOkcOsu/XYHLu5KqpCuBSE9f3e2ZvzasjfrDA4M2VL0kbwh9
P8dYz9cYIAPrhbuh1+g3l5QRcesmb+tsl9omP/ke/4ItQQR3Nxa7oohPjVV2o8wQFV0Yn/PJ7EZY
+DP2kdYhAKsSAh0pk+wxZX63k7c8pVFh0AXm6X/IkzShaM7juWJr5jgyWjoucb5ehjW4A8qtlnY2
sxFRtr/2atnUPhxSbucW+Y1lYrG2TSmj20vFStlahz/VGJROgvxC5HIWJL3B/Kvw6fWBvsrHdGPY
c6fmYvNMJIePPFr3gP+hLm401o4sT/ZlrEZ2veDZXj68NNFfkS8vaB6X3pDjW1a2eeu99cRUvUSD
naEtGZ6TqmCVBn1I1FUksjvutlhmxyATslHpmzdrxwmd2zAJ06jTfAGVsWa5gVJT6xJeA3cbnFLB
Wru8FK/Su86LWMv8ikecCMb28y0CHIsxFHPkDIW5vaO4Ry7sN7Gk55cHCBzGBLzrbZ8y/ewf1sWZ
PI68gJuqptYqO59yGw0EiF8kuecZes0PM8DYxAuk0/ecPWnOx+xlCZdVVDbx+Tda9g/j4WUgLukF
EI6UIClMf0IB0pFoCZWI60DyZzB2mX+/nPLapKDjdVboCfq1nBTxKz8pqTR2KBM4ieAX3ewqxutl
7n0teMYCjRAozSdn/Vq8mTyNogP1lkE3htCBMvTIc3qTQv+WDuW0GY+mwv1aE+OyBxmn+T8SrsnJ
x8/m9gpuJDYAaNDBDXrH0G2+mQbUCspiQlyHzpbpB0CiFZdSwePDa0AUTx+tsw9y6BWT1206f+6G
QSzfhwtx1f+q10+X48boqgamVbPTN4b2qgq8+RgIY81Tap1wi9K/41GlDtvBajfPbmORMoQKMVR4
psScy1Mg6MUZkEGc6s+pxJSqXdKuw4IjZNEFfic7KG3I1+yClv+6uj7RSQiqKtKqyeQ5BSwBZSJ/
Vs4wTphSujuDbErzO1S1z2FxIe0brZpMrqNjLB+7HsociLAGAwLl4aw3CNkc3D0PiQNdx9Qzjigr
In7O0nisctPyPwlJqGlkcn9shQemXZ6SoI8LzQEPVvOB6PzIRJTKGJc6APWCh8gBfhJKFNzREFV0
QJdx8ImsWub8RXmma3seogMweYTUXluQ5ibY80w+OZI0XdNoAunUNBxX3RUyYuD8KFALiACbe+ot
I1I5HJOEtZnVnUiAt8a/9SBVGhDXvdDycQDkV9D4qOKRCMDZrSVrPk2volywjAikemJtYGulVe0e
kPTSq9hm/pjgj6fCHhfWG9Dh4kT0Q1wh7PSDbpWkvSKy+xbA7RPgEpdmJ5XRTD+5kfihFjoXrdLe
YYLSFB2jrA3qGTBWW1ov9HblzbQoX8gUbmDJZzWjHMUBSHHk09Lq6VudG6XYgkWrnGhTMWGfirpP
HJ0k31hGKGKVDBMybRl6+YdYRXgCskEIEt7YUVaBD86usNrrn2SPXGkzik5VTXJkCi80a66jFxjy
5MtQvvmvttFNE50pBxTmt0KtG5uIEHgtE2aqn8kwiIu1hd4Yx5I5z6WqcG4UCnXVbOj+U1e4G42F
nNQJGoJXhBpqbYSbP9i3V5KiZUfvYfWHATBLzhyqi6iHhEMqN2H9ROZDAts5UxNZTzQ2zqzQvBD7
5zODdkw5Dl45GvWrWqnIXfIhpmcCpQTJvVmpAo3dpRzvFKZeuWwt/PMx9a2ES4mDQwzZCPIic6M9
C74YWC+Btc7kO/auuIz8Cj7dEX3sHOIiD27QQHayjD66R+HtA08PZaKJMOM0rbFMWs3dsxJBwNI9
GrvIrQBUluChjS+sp/oHpCJMoq3DmHqrg/IfHpcoy93EEpORqqXVSiUPj6U6WuHKpIFNDfri2Jnq
CSjN5b3IxFvCbLH9odO4axq0AMHtdP7V6lW759Pa/0rlr6Y4POOfuOA+J8cEWMxj79C8WkJuAskI
EKuU9pMSu6I1tuIZL3FsItUTppxK1Fo/mOiQPTeh/kqH3QuCpBfJm4oInnaNM13EB9W7UmNktco8
AIsZ/Bdcj7BJmPA5nHsYy1CJlCrqi2pulBgyoXeaE4X1Cro9PZTh5ryupzQLWhufk4zTbTPyPX3s
SpcxdJCvslev2JJVojCVk7qq8VgW+ifmXovMOfJ0vYDOqEYzUjHYuKVn3bbmF++YDVuKhEV+nBa9
rGddqfbQZKQtedD+3jtIyvJu5aGZTqJaSU1nJlmQyR6c3IK8IJYndvqkWFDyoVbT+QR2yxpfOuXq
Rjljt/5nRiGSkRd1HXyaBF499mYqmuB3CNYfYmXLIANHo1tcfpKeJQ8hcWD4i6AgEaHY5wq35MiS
/EoLmRnMNZO7B6Ic1b7UDWtB+0MKZJkjgFMT92SqABZC7PeldMOmKygKrv9yAAmcjEnFlpJu39bx
iHJ7DTbkwapL+dT14/eKY77AC+B7GgdjhTYBmNY/YZPxcP2y4WUu23F6YNZ/yrNAZ+LvRFpI8ilb
ptcwbgv7RHTYxkjU0dst0K60kDJ0JJRXHMFrtWNZMXxEjyWmPIseVZv8F8Fwu3QeotluTH38cZ6c
fY1uKdAt/1q92DlWaN0FcQAUBKKzaRmkZBbZFayff+UbvI91zcOJYMvV54GB+rhFNSH81fHCkk7S
swHGLQNBRYxoOSdRApsP/O2t0DIVTNuquCvwngApnNU3nsLS7fGIFXcqqbGecNiOVtJa3fJIDsLQ
/D8i2tpF71sXP8qoLu4T8lt1BVFCOj5xTg+mnGUeqmifMsNFXAXVGXjN5QmIhmFZUn54FsfMaGQ3
AD5UNYC/jdtuGonTsVLUojsSd73yO5u5yi5m8YF4/mpxAImC7Xgut20pxJ4GS/JJ//TPbW+nirIe
8KoHOPAoj+w3JJJ0fqGSNmoDU/xAe2rFliXe5ak/fbFBLJRMutaYu/vNJd8Gx0CWIfheZvfHnV8p
HL95MyhWfC5TdjHmZxS/iSmxTOGV+mawYZI9210kypAhnF8aDPr2cl80OHdwQov/IYOApkqaBVuL
HQ73L3zvvXmuBXx8j6kanPAh7F+EhgInSfFAtwcVRPjYMNaLq4a1aWOnF0ujrHbNKnIfoFM8HfSj
Bkh4W0d0ZCwQpKAaLANlZm5g2vJiDZCdUPeold1+QRAtyf4KxGA6ArZ7cwDt+VDX6l2VZUnt7b2f
V6xjXUelYZbYKMfk7yZufhtHg1QeZnjX4QYE26HwjCN7MTe/opV4A2str0Maixr5bsCIt+9jRZ4k
EmKpZDwu8tPEHEpzV1b4AmjBach2GblBZjbKPGI/VCZ+PBcn4UO1c/jSfOA70jhD8Boj6j43ayCL
EpTXjtVeZhpDvXGy7IbUuigluAKkGsHgcp6ULj00DfVXPmeH114kcroEPg5GINAUulMMx17RNdoj
FPrwZeFx8mudUTxvnVn+pCNpDfbPQMRNbKuM2FwJX1n5FZ6Zo0pou1cXCXz7VE5DBUgnGrEakHyb
AniOtjeMBRiENqRBrP78hDLDazTSEL38Kfu+/wq1shjjzEeeRUPnQpaj1HOrGbxLv3JgSL8PTwLs
ocMY5lblmx/FmrXxcFhcUvRKvVmLa72eiHUn5zp4p8fQjQYcq+S0x/kiQWtmkslayXOW9zDu/QyA
ogBJO9oHmLhQOVvwA5YsPMmzuzczGDsvkxO7LNpMj5JyIaIB4O3zjIcyXDSRBGyhXfYlTEB9u6nZ
I/dg77uNmQ3nHMCY0dKX0st5BB4EgTXrmcNb2BnXN/JBGt4O3BRYhXPaefkhAfYbxSOx/FU+xeTe
AnD8Iu/CaXu3kUUe+8C0JUo7YbLTZGE5RvUB1pjUKQs0qF6jantkwV3C+S/yVlZFehekdaJxM8aT
2QhSruwj5S4TlrbvgPkSOfljcYTtK3/HCa2s+XSEimYl9aSiZyn6E2GIo0oC0rmV8zy/au8KzQt6
1V0PYJZFkgQ6pvDjUcA5u94VewVHVpyWC4N7YLzm+oLdmpyPn23oOGRR2qBQO0qtWP4twybaqPrc
PoGUXrssZgQ/vQl52vlx74tJ3RBMTT9ZJ/7kN7OGooy+NVaAWoaMKu9WacaK4dCkkI0Jl9+0VO9q
KkYxx4ImCasyuhGXoDBb/rY8/H4TtXBkP/5+qn+Vo++GJFXCBDR+nrBaDg4g3zyLd4tDzDMHE0UF
6De2nPgvSpXjEQltogpvnC7GSP30k8yu99f78riYLUMG58M/D7r/HKAwISfwoACk7AgpIlzsnTAT
3gMe0mZUhZvuuZOcjG1/fHnb2ZyEdBBRTnYOEXMu2PhtY+ZnJglOlqUt5jmYGE68FejeqmHnfstE
qqpEZhZ5IjOZwtSW7m8u/tqr3pnZNr25+PLjjySe15NAVRZeyY4+ipBXIezKp0/tHjRlqW2CVq23
T5A93iRv754gZ6IAT9IYzWMvp+obqaoWg8WMS9zTzmoduOV61rXpJv/VGUL6cH4wj4y0BwhHQShW
pxF/Hu/cDvjKxt4O/NVVlxTs9FowbDxfF3EfrnKkHbEYEKagE286aWfhFXiKji3w1MSCuVynUjvQ
8zyF5zdGR3H2Uw9ejZfjXkJBPRFlwzjChd/73V00IrZPUUV+kZmsL+ZzKok0ThUvMMu+p02rBLkk
KK613ZPkSnOmx4olqyDdUjvX9BJgOwmWNea3CC3J4zQgvRw7PqVSVwX/QP7feyjWbHC9ix+asDCx
N+SqBDoEEYzh6OCPhwNKuBKpgrzsCvzytL8O7k/A6Fg5sLc81J5NJldVoJqPlDeTGzAZ4GqxWGGp
eidypYXIYP0LQhCGoow1nzEhEdLTAbnWBQXEixoY0qpEYalM3NKCm2cBCmQA5Gz6VkLVeKC0z9qb
pEbv7Rzvw8N7I8FCt9skyipaIIfMRZsedPxtQJxs8f69FxoFINK9nK0eR0Z9cY71B2mey83PEgJK
qfq2Uy2gLmrOUduzLlhadhHbmljWi1s3Z26il9UoNlfhR4j+pAVvOdCnPp4fELaMxgVmFC6agB2H
DtrtVU6NFgF5QiqXBMonWd7uPmuXW8YUpuAbPLvy9CFQhKmvRYM4d1UgSuNO0z/p6UFzuRM0W7wJ
2KSAAKWqHa/9mWek/E5b/blDoOKGIKrdHbADrr0wUh51PSVz7H/AeojDl5EZumBlp9aD43jyAMNL
rvHRpa7/6prIBD+EngrPf7ezGMgKiKjgvmflPUUTZNi+/YcXehpFJCF34QLZ9ENB5KxCR8K102Lu
AoQnR50s36LCq5S2Zo7huiTt67PSckDHTRESHhHxOT8mJX6woClnc3fs0U5dB5oRVSoaPtrWFOl7
ZB2MZ5gYRoWm/bN8epCwm9duGlAI9TzNfijSHSTFInIpKYMNxZTMsml4eDLlZFOjfOnb8J7q748/
RqVcc2BdfEbYf7uA5pCY8M+AcyjuGFiIsDIN1o0m6gPykzLXgczF0428uh34twnFtALAokfBaV8Q
jKiTvypz+k0TQjtFmUCJrnQlCz9ETP2Y8XxoKgd8Y1Vs1TVCb6kyPLWn4eSwLe+xX54I3zUqHHlr
vih2JqdAkUcH97N9k0NEqDBfJbIlMPU6hYxotlQJqjz9DH/c7yW1axKPnTtmxtLpitTe5p7lRhfU
Vb3lM019fv5i2AYM3+nesBN+W8QMNP4+rrt3WAHMcEfMOeIWaZH4/EwNzxJ9Wdr408GJ2HHGYFcj
k/ep0MExen9T/bSP9iGfd593oDKoq48sakRLgkeGJbqDH/WOTdV4NqlJmhGkqCDcVrgwrDgvYB+Y
53whO06mtuIugwpqNOmFYUIptYTYQO9o5LRkKF63mDh+z/2HfN38C9cuumGnzHikb1ewr8rf/MGX
rLQjtl0iRJb2FfyMdw+dGJwSdjcKiUdkdHus+UWZeE7IZn7TKVdJh8Cg+XA6aVQvSW8RvhzeCSf0
kCURQjBYGDIkXOlRC4It/wofn1YljVbUZfGSzWLlC0FSFyZYJlzZccScLpTqI0qS10BjIQHOhqSb
6PLI4i+uDKnWogLq2AFhlkPFFxeIGpEKBCHebFot/V4iKTtZtlT5HGL4N8RCdt2vlpZrZD2XMhXF
26bE5+8uTn/5ue5AHACwPvrp9KYGQSezpgAw9oYekD5+GWD1zE59fVX4/i8eWF8Ox4lVHc22m/Uo
pqoMs3PYjh8VSZUiHU5hrdOOf1sHLgu+rnQKFiuHh7iroAGh5RfyECWBAlXf73vv/OiFuDFz+lIA
zye8lF5ooXv6Azl5IlQrAYF8Ro90vD8VlBYzK/xx8TAsjA7zO2L7sHIPURoXYCewxY3V9XXu+EdC
OfIr8rdauhTVIA8cN97vRM6l6/hzuRGzjn54BrmJ+pvqJz7wo6XmjWkaY1NQfHBQEwdfzo3ShaMq
QzWP5xQBsr70y5CGoPOxu25j1YOhty7xYUEdoPBJiOjCsjHqXWUv2WMl340mr4uhs6vW5/SBh9f+
5YAefLu4Te8+bsgHW5NvI0Ih+G8IGP1oB1Pt4xy781ah+d3Rad6hiLnN/NH5OwJmgk433Dksy9yM
Nym0p5KTom4UU4ZTXjXu4Imtx3okBk6XWiCc9T1EfJWhDoo9t/g1NFthSvpoGPus55DOcKxJ6Yyl
F64fMP3Ak0xAx/pels8nCz8ObAk0QfXL7GymThDO8264gBJhbvZk5MC7RS/M8TatgUBxMmX8pdUK
jizNLumpCyBMd2FWTB94GU4F/qOzdYQOhCSkrQ6bn9tTdasQ8wasrq8BGKVeeD9X3h0xh5wXxDWI
PI8sr1GzcGPcbkiDXElr2wgFxeif1VWNAGaXvAg9MIqdgJ90L841tH5YNqsyiz8UjexO6Vp75RaW
tc5KKvHGs5zosgGNdzEUGxT+tf19I5MlFM1tU2S9Smc1tHrnT1sVCYxqbt3uOnkeXq1iKh1adZZF
xYQQC7yWmXSIOtqcsMFSTPpG+Vsa6wN+uWgI/yx6NSlLQYMg59IOnXZCHN7CrpHTlPRonOogIbj1
d3DWtEfnmqhfIcp3QfJj/RbPgbPg8ltP4qcPuxwbsI4T3KgePcC0DX48OaxdNmlVrKxclp4awYuX
KNiN/sQ1QhVdeoIngzUYbUWihYWjCF32FyFRrT+32393lBXkQ/dgkq/h1uxia3c45+47mYhidWeX
7iQIpTog6e5P0lmEVcphBdmv55stSjbSDzoPzlBdke3vV185YpBW4XLD5f0dwz5J2Tvoj7ScRmTr
mP8KWRNpTmnnv/YT4G+Bd4d/EJ/QwOdIXBsqBvPVmWuoZod0vWNrMxaJ+W/1ufdyYge162tOm5HA
VMZ3dAhWAQxWLVB2j84quo1JOQeGRN1Ilv/4cHDgQvueQDscCLsMDdKmA6HOWe25nWwKLWYZH9Fs
BT3IcJw4KUwBEiT1xXQ19WDGAwD/n0WXp32YUvhJE8CxOE2lnzQ13IhuJks408O/7yGrS+2RSJB8
bop50+azuodykIp8p3LYhGKGpvj+xrqselA0hJcpzziPLtYMN2DD6eted9tbHeTWZjCyCganI+5k
EoXlAhOZvSUFONP2hxzcbuvvG7CgXim2LT5bb1WtfxfJiq3d0KuRzfwMbQZTAbzDyVKl0UrP0ulA
I2c3YNbK8Ha84PXXqy7jrWT1V/FEpCxCPh0VwZNnixlvIy5QoV7aaC3oF7XGtnsH2NlpnZqiPMx6
zohcc1N1qXp31TwW+gJYbb5gal7xFM5ztx2YMg7jR6IZaWo7fe65wGTG7xwlOQH72mMYV3HhT4aZ
0t/GZeU86zrOcJeA5Acv/A+qPkqiRnsqTfwuExUPMo+/QtYxoNHIyNBt6sC/CpxVu3wnK6fQV8mP
zvHQG/kuS16iFYFDXmnUqJhLGNP0b0qnwB1uHAWXX7NdhdGi3gOz8Y3SCT1cr/qQ7EDvZ1T9oOSv
8qdHDgEs63MsHkV0ZiM42fZ2uYX9HwmRMOxSvGZtF4+MLbFboQw97yhRJWeFFkUHfCTGg5Ah35qD
KkdN68krX+gPypo1uR2jgdLIY1PzJ9fbbKDdYf+SFgl68v+ieDMs9GV/QzfNxnIB8Gz/6LOzClFf
HfFWN0Fuc/8OqEUmpPT1r4E9y6kK1Wwtx/oh4wbHmBqeUT096mDWJVM7Xqes8jcp18uzUEYUWUTs
sATJOGczHp3Y89/ulJtUJ83njlKH+bYl18DiuP6SaXq80yILHR9wFZKi4BaP2OZ/DIanfrikDwPK
Uihc9H4hOrgbPmCjrEXoK4lhPV6v2bTPSfD+nN+Zb0PzIego+JNHeEqxKAYSx8taUkYVQI5niT5+
pVOY1wzYkJYvdArQVYYWjHRGoyijRGlyl1PHKbNN0m/9Y7pXDJEd85GViFcGT6JqVV9KoW7xbawH
A/nQOKlnu1yltIawzo7PWVktSbiSxl2ztPi/Pe66HtFisFbRZEjMSryK4B3pFW83McZWpf8KCpNB
SNSmS9Rh0ph7TsdEI17v8J/0UbUeIQBt4ZwMQGQ/lWMawZGdqfu4/0WEvp/QT72ft0A95yH0Ru0H
PiLuyS63WAy1Zl97XXiduLQ/dQpLwXOnTDXYunA1KVGMPPEgR2D6u/UEphBWpAOKBNKAfsnykUyq
/8z6fesq1bgN3U4ZcJt/rkAjTGRpDb3rLRWckcKQ2x+W5xLBBsUJlUDEm/KqVDrAWAqbPQ7j9aB5
GR6WMKM8u0kxT6XAUNwnq8iHGttZTMdNhQWt9IloP7CXU4JQIHCRVL6f5ydyp9JIUh30G20n/ZwG
PDJIvAmiv5T9fbEC1YRSqCzaT4yGZUiaCYGD5DuRuKX+LmIgTHONxNFFDORv6vfK+YO3BsBMVFVB
IO8BFI0pIdxycHiZ9BfkzfhZfCy1rg2qrLxD8CaTqh3xC2n5cVjJfeyoJ8MvyZYd2aPX0HXEHC1Z
lSTpR4NxV+rimj4dA5h7uZKwVR6QrlLSEh4lnpBEzcr6ysSCiGbxv0G3Dzs8F/K6jiEN2t5paBwd
uRQJVZEJlEpm67Svh7nuXGRquna3fkqICbmKdGpIOSahrQEbaulQPNuL0UYEezos+zWDCMdN8Hxt
hhtMvHeQkYL+oqM0Q+K04zYNHBxcSiMdQG1qbf3i+RbxjxbvBcU9Exgq85+5kLQLAEcy02gH6gU/
3uETypczZbrqoWQl0O57yIZEe9GAEJUNY4LnuCtAoKIDcRtHVCg9BB5UoaCPNU2AePp+YihqIekh
CXiYNvoRN6E19y5oPlH4b4pMITcUFi5ZvYth2Q7up18R2/wV97wNNumhqx/mRIZ2/tL17oQhHnCN
+4yKIcKfcp4x6RqrFYyPYfO8X8cgJCcIgVHmLkaIFcLH9zD2S+QCuvvMNmgtXEzDzpdjXViqGse6
K8T3PYTJvGoACThBV1TXZxJRqx2UGhaZU2WcgkIgk7KAUq3IZdQYuG/UuY8OdLZKw2ssPvSepC0e
WYssSBfxxYxi8UNDfZiUO2HBNDbBsWfrwZKnYUJiyPVWJ9VRaiBCP+2h92NQa3qYr+Bpf7NolV9S
5JDd6jPJPhAM4NYutCE33TASYTM6fsRtWGscdSkx237eeDhItn1P2LvF8mQGJyzjaxlHQlX0LGd/
7vwU37Pzaca3mJU320HMqqqqd6bmT4hKc4ynf0sZ/7ax/u8bZeQ/qYhM0/+Xa7AW4fbXoRYRAbwP
La116ZurHB/QJsX7FHvSQhMRrFqyeNnTrE3GjznWTXRBwtVn8lBpW/EyGsWJf5Eg7xrRaoQsf2wm
LVzcwdeOUdhMFQE9wphoyzenDH80h04hox4xQoHHWr4tmZCZP69tFnt1OLfabAdJHbBfD+6D0Qtt
0v8wrMDWKGM/A3bHoofcZFNEf1p9vvwhXf9iTQn7heFPtY9SzvUZPgbgMFhGry0Viw2njUN1KRGs
u2nefrAZPkz98ehFk21z1sSkDt5rC5dZ2gOuuuWJRS9ev357J0PK9gaWLqYoQ9TdFqOTOMZZOLGC
AmOZtKawZ8KR7PCMhOfGOn7KSAh5Mr2x1DK9q4rdP02eS0ZbsCekoAQy8Y0bIzS1aS2KqWBG/Sjy
xFABaOAZ3OqydL5jy3yazEeli3cXIJ1d1LOkxyvysG/3HjLPhfhi7M+wPwOLf2Eog4Bz/7Na3IzI
QgEyzyjnb7UhUObHgo3e7jc62rGI2VfHxVi7aYVBTk+ScWnoCCxWYKsvku2SjQe/pS35ECxUlfzu
BkDF81IVm15ovY24ji58grSee431iKzm+VteOkFwAhVpG4LRNWzHSxbl9S9hFIoZFr//kZviunkB
bhYh3bf0ctm/UpL9exXue/R8AymBus5JChI8sE0oHb9kYbNvSoCuGWrPNYQPfv3iPYIXAK4uQVOg
BA1eaUHH8p9FzFidXGQAKkeMbVxC/KKF4B2fgcUwJLcfi7laBxQmTMnNrdH8bJE2q1sVL2vCfMYk
vVwICF5UZgs7wB1UFVlS8mPuwUB6rVVb/6TggZ6CpSeJbex8Mryae65TKIU0v2ZCIAwTAz3BVIc2
POwEpE/59hSI1ES4+Vnbjs+fGw7phx1OAwdZqG3dsz4LHj2oZn5VFf+gSTVRrNOEsuC3bZ6vgo+N
qye+76xHp7PSeR8ettJB2cEp2Uw+H+fQ3iYwcDIyLYXg9EBOEbDiRyz/pFSol4T9ym/OwfZtssDB
BBk/65b0y4rPehOEvVPnyNlayV4ykZ/z/EVgl0xzYtFYK7or/p5NaGDSVmX+hVPeM82TwVgEjPJE
Ng5Qy54XuBJ4e2yKXKUq1B/cPvx3gS9o1ehcvWlbpNlzNezkpoUc9Xv3NEZ9+diZDUbUsx0eeB6v
58gCOkLxkEs9kqQWiMDwCq8O76ifmixTsDEGCxf12/X635Ah/FXm6csnSYXu0AD84/gxaKZazFqs
v2TuK7ZBlR+t74tblIaT3jzaVaLoezbRmZwEeNiyeRewidnCRGwTe2miicar9OXZAvFsPiLE6xaf
dH2NMrsS5skJ6KGcn8stfz3FGzpvVWOfUkenwYpYGPcNg9HgnHt2iftxHTtENjTreKkyNCxHqo/j
SZHldGTHWWA+HtR9d6ncO2Z/1OZcgNOzbzsliqhGKoRmAaGmuLhzoT4ZkEqEi5GL26XZLkIiQuDn
4zBFvsNlLZcoXQ+RdllkF4AdkkdGNH8tkkqcwDzd6+U2khUB8/QIbNmXuG6p5hJqIAy19S9b1G8s
mFn+1sj1TrbARCQmxUiB5Cnr/IK6tW/EpVP4OkLIb//+NCBQf9tQyHW8XBo65OTfDdKYHWIzLT7i
n6aJjpXl9yoG6UiIpROltePW9PMM8W0RKHOwiNazhYFy7V/6lgLm3rQ9vcxteBOcZG6g3iJJcDpW
KTSK11GjGQVQsbLRfkc4xcLFTpz07brG+HYt132z2aVwd/wmSfHK2GBv0uCEM7+J0i4roJObGdwe
CDIxDBPR8fMJUILp88WwN17aMu4xrwLwsYewYp0e/i0o4EQxzfVUysUHj7VQKy46fNLjpuVe4sGx
bSafANZqhIpE1IQn4+BGqyxeC3oY60bpvWpN+rsMx6JmEPagtk5GOliH1WEEHT121qvSGQ5RvmO/
dBStm2Pxk4pcLgtL9X1O8tG7o5MfUsq6b97aIqOX1N+BFMd+EFYAYQ4T1WK/795K51RU59tSrGju
kYzUT0QiOTHPjI0J5DbLiCr6iQ7SQPwEnfQP+kKXXrSKwVkKuszJ8d9h9zv1xRbLjCTbT+ye3hH+
5A1mOEvzvYxvJmW4cLUJYR5GRJqRUvYypPmFb0dO87NSLx8vekw3MFEvo8BgvZFAPq4r3vMbnfr+
0KzvLeBU0PaqzOUpKBr3gIG53V1F2NwgBmvnWhq5fF+QTrUcYv7QIvvcLJL8IgYfQ0bMQlU0Wai7
J4fY2yh8C3IvZBlhGRkFcrS82PZxm0iEJgymd6Riy2nqlWa8NFkaqBIrQLuAX+x0IvFTO1Vgs06n
Wo2sELvyMUKOJOdtP0aeJ3lT8QRQYlaBcXw6o0+sQndOo7i6G/I9RAf+Gc0UZq4ieFMiZRML6HPE
bBWJjDsGGcGXwa5LgSL/JgMtDTOTDbRjxgt3ClwGVwFrOA07QzTKa47bIsaqL8UUC7G3B+E0bcBu
Wf9OqE/OuYVVWQVPReDE00EDIzJYIXEPnk0ED1I4C6k5WBUIv+FSLLMIIu3VfOUdwnkPoPMvQffW
NEiY8JvaWd6TyTTd1sv+KKXKfkLPzLOXyp0Htm43YajnrQF49ZvbNpL4LAWHqFLnu/8lNiPnFeia
rX+JPWv466FXysWgkQQWr8Mnvz90y9KRbzugk/LDMCTavg9b5AD2FJO2Y6XvfXgy2PjDM6yLsKgK
vGEp1KUZJ46COAcvMQPe10VzoYjfTgEwIy6nc/3qBFpjHgGxQ3+P2Gzwms9aPKuBIbdzSObHYhna
lLOC7Y4nkKJ+M0RZio4T3FN2+cKWQkENyB/Ztj4G9SgcAl4RuaLdErovpQimYsjF2IVej23g/CR5
EFFd+ScvHE1JrsgbFvqOkEnRcdTSdMY87H78Mqgrj8YKBpWtMBFDW5cXU3kLwPM3T4clSJLGlSe5
8hJWAfrjdrVsB2Y2ah+JJUKgC7e6Ehn+eVFjXeMgHDzMBuNBHvoTRnl1JAYwRfsytTcDjoACFnXU
EwqoOvTo/spbMbDk5Jof/2yl5inSvm7fE8QjTge4UWEquOiAuPk8b6lQv2Cnnf6YmCbTwao7edWU
fOpGEUjhv8jjnKtXi9qz+uyPQT7kgccFX9mVtSF5mFFs/mNK3w4DsV9Eq37tcALWyZlpfJailLx6
qC1F71zAgUEYDwYX+xlUPgDqafxwOO4d2mFsgpRFLAWrRHuSFsZa74vxY1adMBkV+elYElCu516X
QRURCQKoIFEpPdda9e6490trpqdIizh881NLEz4fHunjSdUsBpSL96K5I1RajkEXlYeWbK8c/7YF
O02+AKGruJQjoi9j2b/zLD1+wYoKZI60gSluIJYBcjTTrkcEDbvaG2L2Tvf8dCRWcIiBdSAgiqLg
BdJf2tCDhq5V5+INm2NM7A+Jof998cEvXM5tskYi802TEjhdE0gTqc/2v4wZXGbZ98whN9iU7kv6
xJf+Bdrb1mZf2pmU6bXsHkXKKmNHKGkM7l+wAGnQOz6O9AgpKCXU5PsI80qonj7uXiM/E2AXxQwy
GvQipRwSo8d0HLibBgym5t15EX3zC1Dd7gpMUdVY3KUZTc1NAMqCE9aUKLbtnIqHVnDeUVD1A5lc
XJqj2dVSkzD0ID7x7CdFkmyyErJAha7HPD/k4E2uufxpx2gKkrnk8ST6+3AjjPYsJ5WOiZaYvCh+
9PJv3LBowom+8w14o6vKq7T4u9QIJ48THTNqgM0XYkeBD1jmSKLFBZaIcw0wvXCy6t2tU+AUgRr3
VbZhVfhHhZG9H8xQTVKj9ZRQnCBtXVNwTrf2dug8hG2bD/aORlQnqCx+p5BGhY0OEdQGBIMavlbG
wK+bUwPr6gSGXvne9bw/wyYnEK1nrZqRz/hz4CCMTAroMf1plquB9FLp21DHyfbvjBklFkACk/S1
t4dKm5qnVFRI147SdPPlduSIL7F0/3tTO6MhmKkaKcgQDlYTgZVrobJkpAwvCwndemQ389ywNUe3
REe036VNx9bDaLTwrbwWoEJ4bafzJB0D18foP1KFKBZCU4f2KXn4QGVsillkUg/DTArDH5o/IZO3
rbQJSffuYsJmJAJXY4Ah9DQ79MfQeGlIAFy+izpQ23573pwVBa4m1A/t50BpmJUVV9Tql+ux23ac
yXXhT5PW6heU59ykV8IRPtUKJGXMFjgqy09KOzz6Ec9tLEF9wZpJdWkMYa5JrXGA6XoxSEhpDNFE
VH2ZfHD4nyl9lEmtbJUYSyRw+U/1VUup3pRh/sU9w4XaEhi7Vfg2pvT4ioU8Wd0zraT6FetgUpOR
b8kW1SLTh3cYlqseTtXv6627+eSfyrYYDJyr9ZgVRWhBruCtD0sdElDGwYhRTYNiYuWDDPSJkhFt
HWLfXd/r4aUsXCXrS1uaor6Ffu/s0cUuR5F1+ce1bZi8gdwE3fzDk78v2fOZWHAJW01NzX+jLGL0
S6r2mdjStIDR509XYZTWM9fTpwSmCQLldXSFNHaoXDH8m9P7JC/yAhQTonxcOg3NHIFRhdN70m+y
1SckqB36/0dXdpRA8NKDuNQTWK3WbRnz7yDIYrbmHb8dxjRCdBnnL/QADE+JN0eaKQ7K9r2Ql3rc
mklhp7VLVoyd4rFo6lCebckWOyq8faATXJgJutBptO9BjCKtG1rAAc5xfShmFQkjKGnr0nuqHGQl
EfwAsTYxZVj3nzQZ8R3nO9skUPMClUI1rrEetw8KTyvAwroNa2g4hdMrfpvmGEiHMU7Els69NRrx
B72+PH2iWOx+wIeMVqR1KNkuebVE/XVjFLAlh7qfcipYEvqxq4DkL610ogIrnF4kC0UWvw00Uzd4
/NOsSqVfwcfdI7mmsT/3jAmE/piW8nKOwPHGEkn8/sQMbX5jcpy4w5Tb9uiBxjFFGMTrksel5inc
FuH1bc/jqU7p7cqiPdOA9xfDi83SofK9ANMra/yj+2F3lJXNmWInsTlW5uoqtFkDxnZh+3i/0XKF
TTzcw9vbIUAgFbcD5m6h0t2Bv2THesdIE2K4Da/bk0FHBwo87Lheh9eax33igbUBl9BoSNP2zqNE
9EdaLF/HpiGkTuGXD/ZWSSHEOxvo1rID+tiNzbNFJ3pnadkFX3T2eRH6RZ5NFoeuGzl1qZhSnXkr
sdwJaRLGrO3ujBElepRREw73H8zys6n+UV6akO/Oa9iKe5owA1VM+oxwieI9/pRQuWxc7ARy15m4
H0s9nDUwmH3JCutJyzd3oq/14gQuJKlAUcZeeTYUYWffewZ1QcQl8uwhq1ARHHFbE+WRNe0R7w/x
6uDLe/h1uXsZXsOb4rUZValTGCijHkmAjc6aZmU/xx8ng8FwSxLLyQv7/rQlFMO6J6dwHElTdja4
dnF+ZyoDEzLSaPtNu0GNW9T0bQ7IgLjpkZUZ0MN9VUnknGPjcP7WNPtn+aga48VxBly9S3iJhwYW
6LdMhC3jhS4kNKJgmpSuNQK3Oqd8MNFKhnAk4YqvBgo73VU2ejJ9D77hgS7BNQohEwiXPGjKOgU6
Aw8vLUezTgH5X2W+j90EpItmYi8zRgkc8mI2gMTjR4S3j4tj7eTPsxCC/mHxuk0sCPH/f12kU+2G
2MOOIbgtrKaU/UTmZW5amfjm+JJYTy4T/sn0wA5Ni/5UF0YKwGpxVjUE5qYDD50MEKmCgEU2TLiF
Da6DXkoganVqLooLNE8hWQABSLY+n/VA5hXJ4FE2mCmg8+jKDSN2IMuYVpU5wkY1YghcxKo0pYwy
4IM/vX9UYVGXsKxsErUT8CHcPk88AkycwT9reU+pYq0Q9jlFOdp2xt/gEnBxA+0lXfLKNMJMsLNH
chZzJy0ZuYyrkieVEmzIUsQGufpPIcKnu2oCwHZ/DTxaHVGPc95FKAszLBW2kTlu6fOmIFLBgZAG
aioFHYylv/Nx/udLnzYVw2yJKlu/loPkHNjeDAWfUclxkSj3mAZ6u34muGQ4bAgA4BLOBW+OrFA+
Se12gRSvfrcYBIGsszA270jViKXOZz/YfzGlBF4prGfv/spcmFJwfdbhB5z6eL6A2o1T7G2thE7M
IXmGyPf6t+lSNo7lL5DeLrQrtihvyWgLtMvhGthoc1wh9aRdUvgK8JYF07InNkYb1rhIWRVRlYYk
VwciePWTxpZtLEVxQhXugZiKbiX9IDz/19b4lgs/wHekYbu+0RR3+8hbBLHArgbycH8wCT7ZPwYj
2JX0gPZfw/nG9cgaLw3VUpIh3vFZWj93+yzDnY+6WTg182ER8FXyV5c81ltzWg+LPwOSlLcbGSO0
pPaCkRXyiCYNEfYAdNkK2driPgT/b5g0k6IjU2BuNC/6wIIVGSORqHKR4yZtooXGFCfuEbidvQ21
H5y1V/lH5erlVxXItrp9LtSC6J9j2rItT1uXz6Oc0iVfdwf58Rs98P2kcXxQ1d4MtoSlec/GYrVv
FdHH9fgFu4yGc4Srv6ADXKSt/lvl8H0/FqA40ycy9eNHxA374gYdgKZIQStMSOzXwnrJc8h7m00l
cTYYyCWb/zXfV4OKF/hnNLhu3SjPe7dlAHjUXyAJyfItss5ZJgLsNOMHPzfqhiBdkqkcVaC78biv
k419iRaD/a0MVvaI4zULKRLDXsxaBkj8spNmbuhEkRvFpEkg2sti/Z50sT+xgE0yWgg2rr1ZRWkp
b0z893QI+icFf+DS4d6d1uRr1+W6RAYy2lzDiWjXQtkrH+a9MX6mge3C+CqrQmjYyowCufvy2Ues
AsuyQOKhSkA1iYLoi1u/MKbGTKTdZ3B7Y7cabv9o2ovvwZzdANvdgfKEl3y3oVIwIjN0+PAi3erN
uIPtmkrg9dht2lcb9JgQwkDHz5rlhBLD0M+/2V6sOvT+FasztEdd9jKfREch8f2em1Ch+CZTmoxe
E01yxpFrk5l13jeqxRmyE9TzBp38bcI624ZH1nPF+1yT8Hj2SJtukrZmdlZtyMvOdC3wKw9Tom7t
DRXT6vBu0RACKc9ULMXEQkqaIDOG8ZbjbR2D3nTXuYvF5XJ717G2SuJJRbYYgbDraImES5h5Kn/Z
BcwrjO5w6iIX1xiluV0YmCT8PkexTcQbwLbU3UBGrOsIE84Rl8AtroxvmSN8wBeCSUENPStnNSXu
RjPXDggHVefDFP6pFaYvyMzFqX8dmy80gfBl8f8h4QXDKOblzMwjt+DdU14nR6SYEN0UC3T08iBe
6tW0uPlWQTMLwvvNovkpf2o9Vf3u2fKb27GlpuJF43rSPWE5Bec1VAvvryjojWrTbRuNluE8zCtH
k97JGARRWB/QzUp9TdR19P6eCdfKGk63NtrvmsnTtx6f/rliD5JzfA5XWZSOulQ8smGkFXrw7Rh6
qcLF1d6lHSwt+CSQkqw1414zkyy+gTjF2Q1QlWaWDHfSnWXjlyPnByQA3l9bp5Wp7dTIWML5wHcR
stO5lVVl08uEMRNLpvsg352ihdBTzWb9mTe7wEOprhqiP2Gfin26MSQuWe/5c+qCPhs1/Oa61xJo
1uxMNQEz9mfusOruNWuz+J46apaqUaW8ankKy69jc5MId79H6Znr6KLaUYx+CxZQz4Nf3yHO7zLB
PY7lTV2VmcCnHmd+3mGvevcRJ/OF5OX4AU/99HmHAQ2HNzh5Z2MNUWSgxS8ZERowH5y2rWTRq/Y7
IIR1T+oTY9006pQQNhMUDKoP0T99Q2xCJMrVojo397CI1Rjn17P8vVq99ZZ++fo5O6LBZyAkUQWf
+5fxyzTu3r7G+0h8T48OGbMTr1JlpqdkO524FeFv94bns8t4x0rDUJ92nfjYG9PC9fhICo38fGbK
fES2J3d2mq3mzRsI2Qyc31Qb7GpshTPjdqyz7cyUsQPtCqlx5qbmAdjmZv4xh0khJrxTTbNXk90h
5Zi4ysDf0CEnVP5lswhxDn+H5UFRn7ZoJd1A8cuOH3T11CGvwAiSZA8ug4XyALu2Nh9YCd1oczl9
m2tv63yA1qepY+MQ4Eh39aQ0UpImjMnnUdWsmWRVxsto/cl5zdkDJy6EosMToTOyo4aUdJLdWqMB
J2rjhqfMaauA9uVmWephhips5VEk6gT8AS0JVsm/f/J4Cfzp+uUpX/re88+XouRvIZPUC76OgztN
JCl631atOlJaVyGhTol6ORU+vIVkLnWKhZduOa/++ovW010uegZ2vYfJ0QdD9H/XtM6g/Yr5gdDe
7VdcNy3Ybg+VulcFFgVvkmIArQF10VsQVyXbupYhLkYOvnw/Sgcb7gHbGIm0WJ214tJ2BLN1BcC+
m8umE3uYtL1ZMudERUym8qYI6ZqyuXPCfeHGxwIs2sUDfLAFxG6th8uJb0C9y22DTHufSgKjMaGe
pIJ/VIybps6K0SKKrN42xHK8ttO+JlljV3UBts6KbqbYFUJ3v6U7U998o3z7eLAi8xz8vELH51LZ
e67PMOkHE7mTI6p1lB+WQdtLHE6FwbncKdAL66hHFcx/Mid9NgfzfrztqqLPoFqdjuUIf3TKQsju
MvU7EzL8X/vQY9txVBHWHypM4K8wEJbiZm7Gai2cskeNr4Dvcef5hwpMDcne9PMBQndpi2vXhE2L
uxmTKZ/Z8gQ1BUTc1ONc016jLp5Deqg1iuKuXwbZ42em8O5ZP/yropZ/mF+hYG4jGgpy0yVqy/kq
M7zyr1uYvkyLyiGzV1//hAE40LKSK3QccLPg3Pv23g7i0YozVQMu9p9ElMfralyz2fsfCMWY9z8g
4XW3FAQrpdV31RgevRdjgO+ZWa8dOxFp/ARZK36ja4WUL3JFOi5JlGE1yyhahIqt5gtUn7nKVtD8
JiRJc2EMvvmd+Na02nrEOYenVm4QpwWKQOgbBYYaAbSj6VJAiSC2d3Jj5taObHDYAV9H8pLR+mbW
JewHakbtPBxAv1IWh9Lpe6IvGhBrbwch9qs3HvHxx/yds5DLcFo8OfaFd5mCz13ZNcdbBTgOGhM4
LjW4s3cTkr7s2hJnlQsMhgaJkiRJGDQQMhvC6cewW7MyTJW9zkssYJnR6dzFITKiZ5bNC7OWe2rV
LBwcdzmYRrBXe6160DVAMJFJ3MxIEGFqSAguAhAfsyDaMzqf39OTvhN0nOaqzJRaWg51Q8rUIBQS
s/guTJaxW+sTgA6BUvyghTpiOVUrRPTmTk7re6wkUd5LnwUbSsfE9aBkOZeIdcN+o8C7s/Yiirin
nt8MErOM/lLQR7SJioaUQKhK1fCAgd4cXdZz2LbZ5soWIEHNiEl5UN8rrljkpcNfEbKKNQHq93Fs
qB6bsOy+Hn3OGSn1Ays99c3mdFWsYLPe7rNVUj7kYf4JnfBtsG4xKlBtFV4q8peaMA+Pt6FTTkqx
BR8C7ur2BzJcRf18tl/vbhvR3vPcEiLfZkj8nzoOp88AeqaJb33Op1uPR3szxFUfbR1ir/W9ss3w
3IZKR2iISeTtrV8aeuvAo+GBPLtdvVTGrIfa+TNfEeyoejXrDSJFJ5/iRo16iaJ5C+qERYjkR/Xr
EFzRe26SknG7i0/Bod86aBzrF+OL2nmGSn/J1KO4eQnkxSwUMAYOK7ywUIVKiXlqzw7m27cFTyp3
z3zHz2Pje5CbUFQU2zBpbK3jJFFVrWsSP3Zq8n2gqpYLxfZiblpT6NcygzgJYC/rHBr71Jaept/U
3NB6N3Yeh5bJX4p1kdwLBuajfhxbE9vBh+vVGYWmPxTlefUkS39ymV3E4s2Y3Cu59jAnxrP8WBu1
wKHKpWlAdQfMuzELSzXC3lkwUm3TJWhWYm8rYCe22sk/B8UbbYeSZIUGH0xaPZN3W3HyHQ+bcJ/R
WXAzyrvKqk8CMhHOBLtlxhAM2XcCvw6wt2SQ6FpZTTSKIuIkT2o3Fjnct7okqBOBIVC63wvCJneO
TJI0MsHCinkyq8S2RMuOiuu7cWhlte/FzESZOTpbooHt3MVFC/FqEZKr05Z0bAzaiBcJd1gNokQX
rWmSS92q6G6BagNdlWV/cD+LYk3lGnjTto37sXA9/9uA/jPaIR7Tw/QUsyCtcHD7ZxRu9g72VnPH
vLwdXbJcrPADhPgopTJC7MCKGvNo/zC4D/Pv0NLrv+2gxysH6QB1oALZdgrhcB6orMddzrADS1b/
69l9dJlKalpI7Qw3pK985+QE798qUYd910qAGCKXP/Z69AZIWCX2rE9S4lEBVNySYQh9ZGPkpco8
ntigKgRVsmOY7zZ2dktfhT09Qt8E9IgfRpFSBGtSj5PvrNsjqwxRhZ1Dyunaifd3+CpwMaQOG7FS
1g3vFe/coImwq0r8qJuJvItrvpOIlu/u0d44citRbxPzEbAq07aN8u2OheRUB3CMvCy5lbvncSwz
U9BF2ZsOe1+0f65mk+udfAX3POkiuvLzROrbi3kKpuVkNKRuftFseqianAOhQ2TIbLlV72iHbk+t
ObBKDhsWdWHdEfEGDjapCjPBz5ClYpzYMXxfSWHYVsL8i/R59p0JTWmzLoi4EYFA3Zwfz1hnO1eV
+lNJ3+TrNg8b2rO35/hqB7OVdgairgoJsXj2c46gqG3Z1mvtknpCTMmU5N5w9HuETYrC4A2qU4Zx
7EUVajVWxZv2AGr17NUFoyRtjR49gge7cMMKgBhBrHmVw6n203TyD1yIhbdSNYvA64OGKlxicP6m
aVDxClmLZooaoMDpkL9R3je4Su67pEPTEML41KkvHOBhnnwtkJsu0yv208Z/YRbeaqwth//W68p0
Efz4mOKkA7wsw9K7hHM7LjiqA7RKc52R1kqKKbtTyY3pmf202yuI+qlrOOF3gfk6/1dJrgDQkjDP
RIM1ZGjYb8zrJzl7fGiSojoaH6FTtd2wRz2Y4KsV8ZCH+vkMDw1h/AZvgOwFAyKJh8lh7NTIJVzi
nqiHStagGeuHgCukZW37fu0x6eQFLkCELc8xoJaWMzmq6OKbJQshhmWqmTqze0sksusr/R5VvRyq
bazpbROCbhDT6NVuevgcatGV0BoeahWMs533V6xlXhtkBoeYu3/kxEFJoEzDKD22AVJMuPLeOpZO
fA4v9532vHHFQ+bJfxyClqxmK9tkw7udkA4dyPH0okWl7X+Gm/MZpZtkh8mbYKt1dp04K+zFp9QX
T95ix28t8LRW35GOMQW5CvIUwg5CQpLNnuqkevivzCL482qN4ag444RyRG8pZ7dfzWhxjWr9v0A3
Rze0Mb/lMa5EPhgbTduyDM/GbFhPAOcI1wbofotCcVIsgecyz2sevJZHZGZA5m3t31H+jfLi3nF3
gtINmh1xdOwXye9NGZXnjxijxpS/rvrqx+8QqWnCylfyTImTra0Ofg+cyqFZTQxZDFHuk/uM0nfE
dvMfq3L0WGtQOSR4+s76m9UYBQsArRG1S0Q4q3oGcTOZlOdYs+i30tJdKZr0QRVCBxLLFVPuQ/i7
ORm4S9cssiJh015u5ADoPnESu/psJ07CgvZf03AJbpwPCleQydZUhS0cvhbT9/AUAUuKV8oB/wQP
rYnEpxiWg9j7CTqUNqohRSUf2BHYoZ+fuuKBCWXyiwbNuvSOylR7GL6rGzWnngNGI2Qz656/wVxk
4HIQ4dlntq9tdZUkmK600BepGiE6rpJWwiLVxqFBsU7IA5ySrwaCyHOWDW4ZYLyjhKxkUZ2OZhGr
5m+k0s4wMACiF6BkSCS4IsX5bG+D/CmFoLDQf4kqaHPUT5SwbvHRoU9+kgk35vZhymhvYJoLGC9a
X//kxORAbqk4elMULHw/+/jQVsS0SRQpEpTm9+78DadjnfwLpH9TWHtB+nQeOIkSHKpbrUwt/6MD
5Qu08Fwaaz0QeebRblafLETNkXppqOySykuSNl2Z15xEyfLLU8eLusKjUS8vtD3j7OOV4qAFIrUe
iw/attJGYLSACOwYCHf7klNvgKTLVzAl2xNqKu1j1AGQ4HpONzM9RgMinZl3VmyxktHR8zEnw0cm
rLDobk4bkTgZpeRGn7Q2g3VHYF8ronWC0RtP6XxIwRaAUk2ApOBNjYPB1qsJoGl+jTAcd+9GdxEb
k3dhDhCJbWVIpRdLolx04FQ+v0G8UqOWyBDAQsQ9ULVtVSzvAVc4qFNXgA4vIX/ddZwPhK2LnDgR
k7dYsecBxbnvrSqe0uBxIcmnc0EC3Eo1Mh/vjKNhft8FElWfIKYVYAX03KYRJTcVE/p2+ts6zFh0
63wEpyDCXHaNyNwvi9tWslgrLhaJ7Jjx0V2gVJyTzxt/01xyKZD9Qu2WRU2GAcIcHwZ+BKGq1ljV
ijAPdYTrPJHXMoF3/KLlPsYX3QUAY1Au1GGKHZVo6CfQCdOyyCqKkUpZghYaTICE5TCqrufa0T2q
kIi+G6NM6WNoT+P31Gh68UDbtK20IUfG3JdjVTF9KJBnzZZIWjaQAXeW7aNGJjbC3MhzGXN9Et62
gt0Qscx4XzSP48/L/kwDP+d1h6jfiyukyp4Loi6bkT9p9URhz/3y3GnU4RaGKMetsJ3rN2CWgAu/
Cel7nXWmKRiZk6RiOWYMpweaEAyrRch0X5uzjIs1MRWGw4ibkFyr8yYlIYeIH0wiUdJtaaXpAZm4
Jd2Wr6HDkddFf7QGm9gCtAWZwxRf70QAEqub7rs+WPsGgJNB3+wZSno8Ceb0aqQ9dx7cNVe+s+xH
T0vkkmM5WAr3fiGjugzycJ9VotFtZaqpmeiGxHXKSrpfcE0nhzIWLR6nH26hX7w8UfOT+lOLG3Mr
K9GpPyCHYIwiRGG0TDUa9RD0AQyGzrXsM4CQp/r7DT2iq+5Fkwuf0UGpA4SZJQvYShmY2LtZtL/t
vMV8+BQVDAfOrWS6JRluiXeBdiceuv1r/zG+0V9ZDBfFIfkDeF3dv8JAn3NeKXRMXEBTwTnULzcy
x3Vd/88kuQXKEPz6viOs5tpTd4yGuaSHGxs8spJzivrK4u7unl7nEfHBhM7gHYzSNfNA4B/c9aIh
8GdxcAVHMVw6MB0m1qbdg1g/eqg3qxWDAxgRDXUxR06288dgi/Ecy+eDzMezpGRhoY74/fZSMh8A
W5ljH9qriVOAGJBQaSLtXNYNOO3XpovUTNA+2okE6oxLWpMWC/FCyIlrlLVV3J8K1mpYOM9AF69a
mdZ6/HT8Y2prvSP3fLokOxm0d58N+Qqc4xliUrgkc0TkoAfeSDWmoGG2b8IJShKOYdVHh5V4uQXL
E1pUIBcbY7DezE5yYn0BI674XElI3HtaLHbzvjFXIDQZ8uq5ux+WCE5rHDTEtYDb5aq+o7T5YfBW
QgQ8xUTzDjkoyKLSYA+0rAoRuPd6kbB030DpqVlfnywj0DIcTnfVrvfWpc2sn7TmZ19x8FspngPG
YZcNkvr1s1lf2ACMwE9hdH8VlXq9H0SJXuYxpF/K4DgNFC4OIohuI4tN3Cxvr2lYUz2gZCfdVy6o
PXzrXeAsZ2LxFEY0lEWBaWNJlQyd24V+A3HsxDvDun1vi3mxVdgqFLeLqxqrZHk+UYSB+Maoi4HC
wyadzlrtWKSgs50guRlut18Ex5ne0i8L0BOpLrlA5DEzxLaZkDejSOWE43hiof+lAosd7TU63unK
maVz4UWr1Vu+zvWDzkg7vDvO4KqaQARgi+roSTgapFFNmBE3pxaOrxGHWtn2aOEwxpz6Kz89ARs1
0KfcN5pe7YXAnzkM09M1nLScXxKGsDolbaS0CJOmmX+lO0jx97yoOR/VbGlXmD4Qp8QPGQ2dcshe
YGxzLhuq3glUYPejKGoVMSeiONZa6DZz2GNO1fiLTyTipFHwJ8F1zQZYpIj+ImbZv9l0xrWH7jK1
ZSZWGo5abL79GmTTq0c8mnlvYt9u8HLsurqkRuIdbnL1DNG8IVUOOh6ZkrT04/LUMqTfJJsJU9Z9
pMnnok1nepm9huYjKoCaFu9K0uZ0PF+T0Kq42KiF2N1wImPpnAeL0R4h6RCv0ghqPKPJK0pzy/Qq
0huTIOAc7R49EW0280s8G/uSHGMKU6xQT+8OrU0O8Vmei4d2g+Rd6upnnj+tc8H2qMWnQWbulb3J
qPtfyRGO7NqJ8zM6iPMHpMs0kqISM4b7+JOuzkMou7PmRlmZHleHHPbz5CUUFh2dolUkNWdHCaT0
K+ZVYFs28e9VCSJGBEALILym0hY/+jDJHM+6k8UQzVRCPB7SCB64zaWwJ8nAkikEm3PwpVwp7f6h
aprysUF4ZCNMly0liy/4tKNOXp/dPHV2AjdRLlROSLpWIN32Hug3HZuvXV3BATjpbQNMuJoh37WX
BJtEUx2SUVDtDxHFwb8XVJa+eqztd4Ksj4u2pBOU413+PI+ASxXElUSmX6oZHMptOO/9inTNi64n
uOFn7UYSxnvfNVnyzBXCR2q7RXk8MguESRjzVH0tYr0qOp5YI7Y4VuAvp0c0gPAT/cAk0713w/hV
rfWdlVKoIgc1XOfFAhHmFAdpj7hB/bD2aIa27ZPoHzORrKX4aG9YUUwDJLzR06fjYTn/o9tJ070N
VhxUF42KPVSG7RnsS+M96ddvMXfnn3gKg7Vx2hg5aR8iaBMJ/acPo3qfmkJHwKa9ZpjcWZylwzlO
H0Yu7dqs2c67Qsc8idhb7LTKiDrzu6/2Asv4hnn9+LDZOv7dtJyAYveXZyoPw18sJ18QYIiOWmsB
b8PpmO2BFH7pDgDxhbL9U4j06mZLl3vu6g7eWw+VmVnoXBD6vutm4uKkxeQFoDbHjRjNf6JPWsih
fcuF3YcCr9kHm1rVm5DPCHy41aDCHmWarh8lFeLHE0ZAl/bE2NcAtHsGYLbQ0YFsYno2czFmu2nZ
dmlc3C3OFvTVUlEUZA5Sff6eICk+TIiUKnHuaJtYRSAjfwxYbO1dMD9+xKNk/FggJHoCVp6efdBM
0jelhvwAr75t2MCS401n0OTEvKJNL3I4voobhaYNpC6xOhasJFvCHXb536VllrBMbVmd8kVBh3ID
9betO5r1D1yaYEJ+pSpLHfFIV/qoBtuoebq6hunIUKZjeoNDQRC9rOP1xhiS9UU9qSxBcHkpjuR/
Y6CCTyqlyS4NbmeBlfKuK9yqoCaG7Y1iejrHF3bsQQ/pi37rjjCZBkfOmV5wNNebZEluDJCZRiYV
EtGY14safhsRKveTVVm35UYyY3zyC9qoVzq7cwtkd3qvZMUJonI9jswR3/Z2jzqMFwCluz4NIsVh
ZhSOxVdTAAm8BwJLH56gnYmGYLmuTaTmz8iXJXEdQUzMRa9Pv4r9RfqZOM/ff6BBf8jCLLdSJP8o
vdNKNxftw7X0p3t82v7ULb7Iyx114HnMoB3lZBKquKkZpTzLFw47uADMzqgbssNqNQ/dY5Py7SKN
EAo00GQzm/g8Vn3jg5qGdbcIuERe5BJ1/GZPs/q+fcPeYGKr/MAWDval0hHXRIwVJCCeUzMFYJ+h
5AVtreWqlyrsECMwqV13x8KXSjWwdqLYSYtnyttvATaLzyKeBl8GiS5Uup23Imzjyy78trg1Mmnf
egHwCURS5WBq8eefsEs6bbScAQinrvuq9XWiq94Go0zg/4o0L4qyNhQJ+jkqkXs0HEuJ48M4TYF/
/4pb5AIc0h9a+QKeNhvFvblIwUMsNRxneBDoY8tV0ULfwAXWm6Lx9/FXVW3iDwkNO5SVFrouPtt5
M+wDQ0AWbGez1qmCCkSCWSqaGRFI2mpm8y6qr07SDTKOsyOx0Lx/jk2GQeSn182JL5YWt8hH6n3N
VPWxzL8enj5zO9cbE1+eiaghNg3N6rGjSYLtOmrL+0+aUy0hnkjaAy7xIHbiXKZkFO2dIooG4lci
eCNbuXYYRxaZ6nVpW84aRARfEYx2rMZhKAXvphXbzr2TdLHwQzR1glRAH23/OMK4imwXBaK4XM0X
orksNBA8a08Mob22ce6dqEioJVZXlNJudoB2BqKPda5AXFu4mgZ2p7IF/DQP/uGgXLbENRZ1Uoxt
I1jaV2YP1Thbln0n9PcIvMqPl0rEW8dr7fjtQ4dfxsZjOOupx+IGVHxc50d3Wcq9Bj55eCFyA4l7
5UiK2oKeJZiQVv3CjQ+Gjb6h2inelPyRZ75O9PYqsFYc1aadp+ZyDqPT+uXECWDK7n/GbMrwNmVn
33KUtpO7Tmd6JQrAIQYYdOTWDE4LXS/gIn6SkKKTO/U9XtZ1hCNk3rX5RoYQteqESfE30JzULAD3
Bx2CCE7Q1PgYXpHmeCCGbsbTXWMeY31EkEEMebDsnqOZirzP1BbR0DcKmlqBnWl+kVejNZUp2Ct2
DPLtz58+Cjzy9rcACNMKBFExkMv/XjTYPic3kQJ3dmVWT0V2+fHnxHLTBncFEQWECu37kH3YfdyJ
/iaT5DJQt3ep7oIrU8rd5NCov4mO4O8slh/loA7mxYTH1yBWQGEso3JMNhLwZ5H+9XD1qmhuTkTK
agsJmDFlCPy67MlkMSOmBDLu+RWuQTh+bYL5Hr0Tcx/vv20d8jWrABdpbM3sRDYqMKoiCpG0R3ju
XNj9NyMHwWk65wq6TFZxKRdNWSAmlZvlnShO/76BhmN/N/I+td4GUVOSlMI/YCdMkS+cpxpv0tfy
L6S2ei3Y5TzdCjDUDfXnvJMJA+nRboajC2nSYDmpSCyph3dXNi5jsuq2oIsO5+89VrOuaN5fekyP
lRKGQzC4uZl+2r3rwqjDFe07OpDGLYEXwYAjVSjBHKH7RZg0tqBAwsGHX6TxadzJPnITE1D/2qh2
V+JV5KHUvjlMAPqBYao3q2FXaT7gHD5WKV5nuQPPuGCvtDMIz6US3Us9gbZMtMVOxvsj0vMsLRma
RuIrLEnptbhgLl17suhYUh0hOZkJNjFMgRAnnS0sKmIPMdinY9yNrMApzAldjiYicfnZqPQXowcK
x78ZUPlxHjsPPa+1g49HuBGdyTAzKK62K9wmLEheDPRT6ecg+GU1Pd9S7bz0kAekybxnEjRISo47
byxrU2KuPDXwCTFQwhuWiQ7NaVtES+wYn3xUGOyCbjKjnKooi+WJ0S/NT/W5HX7oVxHT4tcmKFxb
2PhEBpBRKRaadkNppwvEm1CkZKnSY+v55CdM5M14f1CvUTzbrVaywdOUzvy9pQA7NhnqmaqhTmZB
NVYjEQZpyJZI+71lUH/piqCXjDW80njrY2xQQdCNYJ6O4HJ/TMk1ezb8kgINbZnAZV9jMO80kESv
8boJ1rBd4CWrSc0yt8yaBnHhtDJu+MxHYHiR3mkIRTa72TH527VKrlb/RjbelQWM118Z2QSnIuT2
XePLFOyMYQlH1SuuEGmCX7VBAeGL3esey6GKNMuj3eKRN2J5n0NI70jFA0t2eS6QNVQCbsCBwXiF
vlkvDoRTge3zjpb4RSXDU1MzpbCoEEUi84bzhelYDDZQihth73HgwNanEgEujLXN3eAQjmXcliW0
vcc8/KQE2dbVDV98OGgKRKAU/ePaPzhjK+f8+9Sa+TYG7GWcPUV6j2WB65iqlzwxdjFoRkxrhx1C
tYiefMROJ9CB2Cls0EskW72R8LTo9jbXZ+uo+Lyd6/hatc+x6PQ/j3Y9/wBqHphGc0qhjwoZMVTA
25UhgVzUhu6js8xUr42aHhAkZT8yawDwF5WhOKGK47hHDRit/T82AHHxykloqSzPpntBywfYB6Rf
detHHHfRO88OBAy+OETmo64nafWHGkzguPz+x23OrExiejOaiT0h5Kba895ZmwPnkFYoTIwORXAK
x+2HK3ij6WDjH+op689pqZdwH86Saf+V1MnJ4+UkNL7+klDd6NBNmxAnIKWB5k9rWFXfc8V6VlaW
0g5DJ39o9cwsrsHHWXeTGBy9cCzIh2I5NGFoUpqfrCbrsUp8oCV4arsbut1NNkOGPf6j5BlO2d5t
gRW/Ulpvh0rjLxmdRLhubQyicJj4hHcj2X8wc/JS0U3wHsg2PmAQ0t6KE7OiHnGSvJARHNAGajqX
GWb4XeBAQ/6ahFd/XgPJT/N+2dmzCm8/RwCIVkgEDSWLSrA+o4hkarnfoxsFOlgNCCQeptjRc8hG
2//up+DCkfMRWHK+UDf8oKiI7/WWbaTj+8fkp+CJ6TwQ6Sk3tbNK43RADqX7ABR+AtCvAE5+lqlI
OJ5PbDnNQcIt2MOi16TI19UgO0nBDXy3zHTgM5dkwnusep0oFZX59UMeRYrND4D2nYHfx2NdcB4G
Kql0ZwPXEBSzDfnvtKtw3twJvMDg1maIlEGGs4HGkSHGP6OYmWUGvH7LGkN1Yr+c5ozl2VvxwH1b
ZFvLT2DHfmloRCHI+/7H9AXAeijBLosWKoqkmoRM5jeQGe8AtLjn3MrGND6JimbE/iDlSkTHrSl0
24PLgQReWmq9sY66iI/Db9nxotD+T2mM+71ukRFVvkH3omnu2Lk5QUrh35OUIYAXpKDgdifiwF5/
tAGF2oAgJXnp0hHSLYIWJ9+P6A5sLcLPDkibmB3+VRo+UzOmVVfpdKOj9kQqLPUiDdKdqhKhd5bQ
MGOMMApwEmkMv1CAForGaAdglmRlA+YnVrno6ty98OTuZGrcGlPk822wDuenX31VAxZFQMs6mnxc
1xaWSAb/lXdU8uPdRGrMPzQhp95vtyHpczz80RFl2TWIThAXnWFFUIAEggdNTkFtYWq9L/SMy+yb
2pyOPaTTDeuI1bUcl1OwK/h/gCYHIGPJQf+slmWmnfKz7bHkgUPrIqSHdYGOByoBKM7Hr6lcK5RZ
bNN1aEyY2J800PgGYYDUnQaH2037mMC+DKT3u4E5JDO1RB0rO/hqmrIh6YLukSP1V52DIRqUb6FF
OWrWzlLpwR7tHio9YLiy9ZVwLlrQq0pep8cvTyEqt9VLlNrW6/YOCNgq8lrxRvw0cbefrhCpoRtR
+6zDeu8ee4PPw4+QLbW1Vp2n5xGpPsjniyfKVLCDiPZo7YGWquEgkEBD2w6yQUZVliwaeyJstmmp
tarfRsLh0NLZtnD3/SsBn29zOTxmQkJn9ENsGPYIXQRjsO6fiUwQM4dOjJo83xWS4CGJvjJoA+0+
F2KXPHF/L+LqCB5A5lxWnsLdWs+9M5WnPiVIK1Cm1mmDtNA6D7bi+3YQoSant6yhwjECsV4GGHsl
3Czsz7xkbwOmFvXXuCp3mQRCkCqPQRqDf+4nLOkeEoq0ZlUcX/+e0uprhQJhkALUiD2JsUnDqLMd
p5obIdXxEKN/Q0VKjwaHa07KuS0V4jM+srvpESJeviynTB+XNa5+6S4kGzedyXV7k0nPncjmzyh1
8VwMpFdf4DvtWrDyaA0VJvXeJh3zQ9dAEGe+HAxyJPxJTTlbNlrIR6tkce+EM4gKwf5ZAu7AJepi
XtCyuECjo/UfHc4OcAoc6fpSUCGpqQTkJKv7CILpzd1p7JP7870MzwzrMlZSAq/QzXtQFjy/GA8s
K0tNr+qZS0naVEqtpHrlVFX9gEYRPl1M5F4sMuK7+eJda71qYHraQDltflPjaPdG/T8x6DTBTSI/
zD7oMRckvZZqaTeo2+bItN+zQRgiHqKhxl6kZeQNkN2f471qT91UU77JiVJOrNgrL3VL405qQ+i9
PwMLUf8a2CLjiwy7Fo5ITlQT4VZY4+4OvlqESViopdlndO7f8eG6JOf/Znj1+cL4a/R2DwbsfGd9
PdBc/h2K++AHqo/TEwUJnxy0lAqLHamvIHc31FBGEFG/AGJnC3rEwwBzWj9gf8Yh97qBA6U+uIEU
K53cJbE9Bm6x8sEvEvpdtzIybmaoDL/wv9qwVV7ZRVc2llrdLZmoFeEFpwsdKNr0jFJdPtL3qJcL
RL499Vdbwip2HrWBTNS0uHJ1TiaVpKtxGIjtaarx81LoIKCGtokg1a6xTfXbO9dHx0mijfu9XEsp
CkKoepGxgHZnjYMD7Ak43nYv8KhD5hlmGWa451zWUi1cc8oRI/w0Dk857dH3i/lIl7mvvebNZF8M
6VpnWMoDoMSgIlsdk6AuFFeBNnWvjOSDMHtQpAztSKiIWxN/G0a8Vx7R3COTwNUUMZRtYb09HG4V
l3ATLjFKnqqWVY2X/V7zQ2j1fPrxnxWY1bT8SNoXBqrEjpHlawyCHt0F+nj1KyM3dH1WVO3ZoBDe
Sx7YzfEbO4vlKAAfkqAHa2iYZB1L5hqO2qgVlVN/FASi5Yj5KzMpWAJfQHHccXcIVylYDwbStMfW
QFCoX8ugyJEEQY0lbvIaEl74VjIpI/xspec2FTz5Nnl2AJc72eXoNhGv8vyfaTGUXTOZCbOLFtMU
ANFrb/QV0zEQLmvUel+s86kffV13H1J5+kDEtEtshROPXEFphk2q8pkPvvq4fgR2QJ9Tm/ZFbGzf
uqdzhaofDea2ZZTSCpPIRLoeKiH3zWOV6mHxmU6Uo168fXOPu05uTS9uNc5Oqtepds37nUK4vAPJ
cimfDf9TgJ+UHdMXv4TbmMvKrPBMDIT2uO3Zfzbq0Plvoy01PlOyqMqRGqsyylw4MlbaATohVK0k
bD5GuyevKNc8F2GyVuOKF+IyiFL4kbGlT8pOvk8i1IXBCuRhNCUdNkbH61ygiutrQaS5mPjpb1DV
3YmmvLyqW3Oehi2v0tYYmLtbLkE9vustpgavQBVjM/vcnyZwcu/BvYxMHYj1+iiVtYTPCcYVxPrV
n+1lmbLKX+KV0gNszRQzd7iReQiJ5a/r5MhuydzXqQlzOpVsfHeqVoZFOSJarA2L/HAo19rJyohO
bN4hogA2/0N26hYenDtGgFLdB+UTSmK0jIX4MgZpu3i24KvGyfBUX9zt1jNCp5bP5nz33LV36U4A
T4k+w2m1Djxp1WtQBsmki0u+vgxQASDNa1Wj59pjXCYlS+HDNkscEuh8ZIRybnorMTA5upCLOf/1
awUr+uWBW94ETHdW8uc0INYzwbkKM7LsT+ou4syrFOMBftusFh1LVGF3NXiF+GsThhB2pkG6EkPE
xtDTqGt7lxE+/X62bwHcsauO9tl0+4aBG3A+HgNchRNRTFq6rnMe8xVgmtk770jIm0ZdEyy5DeDc
+cdkpbOPY4FidEdKgoc0kk71OpwGEjiTQ+N13v+s8iSNUfrReEFbNb52Gur7YdrSgJElhfNKaX3s
ZkQK8f2wVbyjzQ9j6wlUtvBrmkSUBu72jHKhif5iA8on6KhD+wk5B2Y3bFRRqVTnYGA/smS5u/6K
E1HlScy+XOvKhY+Eume+CtWzMwl0Hf44th55o3R+G2egZJ/+vj7njrrT1zAqaUNXAApYfDr5IgGl
Nrdffxmg3CIC+P3LfwVedJzO5yTyXeLSmjkmVvrqbjAaRy0g2AASo76ETPN3rA0XV8U5lDe3VjdM
qE+EdHKm0MX4oGHoE9I37LjIWWF6bWMLgK1TOj+5B8+Z7U1FGdPb1+xQYe/uQHptjmRUKTfj8hfO
JXRhjC1C0+UKFrrrefM0XcLHxEyVG9Mh9gAYCprxHvw5e9+csNmI29MMu9AJNWa16RCdRFm9vbgb
3kPBl0Vgyv3gCaXc2HLn4m0a/Z3D3rm7A/T2IIf7t1l37hQDZUINzQuc1LPr5FeswKNAASst53n+
M5F9T/HuKF9JyZCNmjBobh/Ll6fihafqVMl/PejIKyN1VqKzcTTBEV3C1j7nLorIQrpKYk6X1LYc
/p8Eyyn0MNpxOvuhUvRKr+bCJQqr5t4GW4jEzS6nTh2GWLQ9viy+7+4s6DQoFdFgEVd6r2N+GjTn
8DGvnvgd01I4dzpaI14m+FErjadIs5zPpDNrHhBbH6ZAjOviVvwRwX2okow6lRE35ZB43cTpgc6f
gqr6HHKvhgrwuJc6zloTOuiFQVTn9Io5Xkn97s+rQfrK368rEIrs7SB2OXVXPbckTcP4VfENmEv/
ggeEMIZYaglLk7h9xhY7fAxDRRn4TiBt73ba6o5HZh6+9oMa4Dnixo3HzE4nXDJCmuTMnqybZmgQ
Fbk+dFX3xZs32l5mNxsX1Kt9h6wNpsv5XMZAut1YjjwoWCm+LuC9VGAEX97nax65kOnPULsfMZkF
ObxZex/UTyNT2Cj7x54zYPmBo2lX18f9x7wqkPIc9taZK2O3b2Var/ahcJ2/JO6YBj3TtlL8jqWw
HprXaPo4qNDRu/FiYoIfup/Gft5Owg9rq4s6nCWgGLouu5rq8gCLPhUxfJ7U0HTPztZ1d6g5z2/6
AEPyXaHnCSGsGezdOaIRHG1Pam7ciF56pzRw3VjpShYIsao0hbUvH3Ylglp7pEmDLuIm6SgCeZde
TZ7WF8qJw3vMejSrTaZBnb6JPpBJcz1TOL0kCvlZ+jdwojRcop5iioj4289NRg6TbrI+k8Q54hxz
Mdzg6cTM6SM+QkxrEGEu9hjQktmhiioaws8FZjsrDqg2TueYfa5h/SrF7ev6hIaKjrPfwhJc90eC
1yO6hPNRmKwToy6NiJn5DZ7UkxdQQ3MXOXYAMm2XDR0n163vDE+wGMofFE2RgvxKNgzbQJE8Hvcr
JttnTBUsboQiOxDLABWx+B0LcLjsJhkcEkMgLxPQz1Wasqol6/ReGvtMeJ3TiEmYp2NPtEL0fLRS
HlWg3JVxYSu3nN2YLWDLNJNG4SsmOh00vdRnEwGmLMd+cRqmpOPFfHyavDwxwljyRJPvpJauXEq8
7bxYhnGptiG/zp40YZS5Rkmsp91+NAA5gcincavkxX5hzn7A4Eb/LWw9YDFso8xVs1H4+SFSFAVX
rY4Ll5ga6fDs9lrK93j6wVkKIlVEKgZXGEcyhf+N8xo172sQHJJayZEEh6KckAntkCu1ElUte9rx
AJquYNp1Ag4heDRNALvJooGT4H2UBX6PxIhguTIIGjI5UT1BXitmY4eYOJh/ge5XZrE1CGS0JhUL
8eRma6t95IsTt+CcQB1gJzRR3lKq0+X1+lvxXpEGjdyqJiZg9NcEkIRIx5MROzadeVk7pWmiwLbY
y6eDMZLL2BtAcPitNShU/yawcSKY+crBkFkCsg6im9I92AbQWdENyVJZLLZyWWe+C2cjRD82TYL9
obcva0YJjQqBRRbMaQONf1p3RcafC/25ESzY/NyfzwCj0fn9WxOBl0d5i9UVHIm3qm/hbA1baDHp
3BWwE+9nnFnIJCAfLYjXJjEuQnTeJMZVgATrlo822YM6tv/6AfbR4XOy/Ev4NQTq90dne1uk9Y4a
T8Wgvy9ID0qeiy/3v5wThVBFBCGKP20Bc7zXoC9icffTq9M97eM0OeZKeTdd0lS+vCg5mKelcOia
Yp85OOh+DlcCqfoASJpNV5GVfyVcYFhI4HmjY/wUCV8Rdq3m/AJR00AuJeGhoyIHOvrTrgD5y2kg
WqaotPD7fpFqKsO63FBZb1v0GyO9/oa4q0lhtfsqMELhkto6ibg+klQSGO32fSRPgWQfqlVvMXXY
uy66oFsWjsDHmPJl0sCQfCK/sxhcg/5Tij64jxKPEX5lWT+hjNoFG4rS9vHjB/gWLlXHwzN5T8Yk
uIOYd5nNkWspWXYUNxEAYPMlWCjPgUHHnulTjc4O1IgFzWesG6Id0i++zcei7qOqZDT6+/2/CBsc
vcxh3wj8D7MiaKwusqUy6Icz196WuSguxDHf7mjTDFF7gjuiRF2iNHJVVZAiA8vlf7oBxDdoye3I
cWRqc5/6LZ4VyJYbWg2uIMjzS6kQfiar77aLSleYvOh/qWpz90DAVBqcK/cIXWmzgMMcQUPQjhvF
2IGuz4r/oEdrlMkcuQuoIJbGJGe5z0n5JK5Yc01mf4N8echOoWU0WzwqNBMCeC/9iLFgof9eT43r
InmMOxS7PFlwllmStE2B2Xz8gowvnQrNOBew/O8dnPTUi05ygxWTAZh3VEYUVEoZGtKsZHeLss3o
FN6vY8yAwramUtQJlW/egLmE9WNhHsqmsmOCGicgQbNuGmc4P1vwNmFV//2SQB9Nat8JmXHgJshI
uDQteklasRSiU1eN3whQ1gHA+p/SJgP0HUUwG8cR+1JBGDz+CBAT9YgW9gqx1pt6ia5vqDjOBRI6
QJjBFd+cOYG/j44yfKNfrdqtFudVNDgzJR20BgUZDhJxsxQ6X5BkEdopQQGTZNzTuSxlg1o7WqB3
IZQwyWT7+v733u3uxvA6d1IIPRG4gsFgUa6d2UZYMhm7FuLl0Fa4DhggczHDt0E5J518u3WsoawP
sU0kHSn9XXPy+LxFTn8pBUHTraEtjrK2wkSb8Tzel8tkgHQnDvYdIBcT0WWZPYuvVbBrve8epDSy
oZ8NmbxTex+uURWu7N8rzh5nqvA172iqt3ojkP5STWEw8wwaIpOVIaASPx2rQhZ9HRTECyQG6Nn1
me+DB9ww22PGfhk1yTLe9c/9rTbVd0O3icyIC5Uy/JKlOn7JfdENvACPdtwdoRw7mWVPMWDvdmB1
uhLM7IE4LxGhK95EryfcbXtWIzTVx6YrLC+9UW1xY5OOmaK2HmQPHvnuf11aLzMxYCOxABtsfyJD
mHfK7UIPsRsyd92OTIlgFEteAegYXR78E87qqlnZRvTKYAR15gJL0DS4o7z5D4guXsoEX8qHKAxE
7ohdQ4MRK2AjKu3fwIWDn5qqd6VeFsezbmSvlClVZ7660qRmktpwG2tH8VgcUiS62ESUkAfjh2BS
U4Q7E2WL2fKHRUh7D3M5cYHrn2mQdVutDldVNA0sWBvCdh5S4W0YHOl4ylrx5PgbGcA/AufKul6/
X7V/E+ht6iIOKD7Erb/jyTz/LWzgOYhSts9PkdvbgQX3Ff0rjoo90gTabl06SeN+ctMl3Noz9m6A
+2JWIqDQ6NMRQiwAphr4/bdQDuFuxUOmnMuVOJuP/bc8rrs0P+73hWA+UfezdxSi1Ebvl4qJ2LcB
X4Z6oDaOAY/QMioI+i3U3O/QJzW1e21JOKjjjCz889ZOj0BzKGdS4fNLKrkADkrCk324Wl2h3dN6
JbAHFg2Nba/eiE6Ak2T7lsc7jmT3RtT91pybHRJnpTHGX1sDh0JV+K1VpzSfft/ZdC0gOGt/qcBH
fIsjSezd3lJHds+XrSW7ZXcr5xrlNiNaqbIYTL+I1q9hgZT00h3z9klZBQmqCjDCR4atRWExzrDI
PRlMGMVTIj4IVEv6caqoPV2hk1U5Nez/aAUJgwvnFh9WT+yDnxSRCXrIvnH6O8KewOEVuzw1jTWY
sOoKyARgK6wTou5R/0XUoOubAo6654BnU2wrkAvHpzqKYpQofY0D87RJPoA+RVrfvUtm9QMorOSj
RJ53We0twHSlBBTmEgCJ7Ck94jzcEmjIv60aq2RxOZPZsjdq/zIjDkRuYfKPFbJ1Wol0YTd+kueN
n/3ohijbKFmXLuwna7OJzpJTn8/jXcgX7cBkA9Y6FZFLtb/qeRs3+A/Bny4EsmkC10oYAIQb+/9G
jVQJaR/y4TtVtdBiH2onTuZ10yN/hwDYuFV0m6per8Eg3rsU6h0k0rHybtPVym8M0h5SJviiCewF
z8pkZY44lqL4k3yUcl1cKyZlavjNCum5EAw7B55FQ26ghublz9jvG7kwlHsH2NbPSR2BiHNR7SDd
tRN9wxU4Dmxe0U9K8vx+kD3bCNOFa78yIZunAFzA9hvuTNXWerJe1StpRI39wlzWzlka8JKpOQQW
sNXb8fFKMz299LXAVGegU7QwtSWPwhkt7RQlvehFJ/cZEi+dMIICIFPjmFSaAV+voWqc7yPo5U9j
AoNKEvhYUnuuxcvuAIVGWR3HwvXuOSqOq60AsbILODZaGKevBYermyQVObQcLnXlqnFBPkcrZv9N
+rABpyQyIAtquFzhs/ctLhpPGD455H1OnZ8rRPJ7bUhPnTEHfosyVLqN+G23Z4/jJ0vt1JhkBYjP
yEPLJkSOg2kFLXqcYmfg2E1wGNAoKifULB+HAVF5e6S4XWCUU7cYqABPVU79EgDxwMaJOO1bR0ed
5LKVxUnTUH1y9dl/F859XiIsEU+SOciQT0aSM72n+e2Nee7eqWjmLM8M+8gzXWjiT86qiowK946s
f0fbUmnlqfsxVJTWj20haZFcs1ySaPh5OxQI9xkEqCzWwULIBbk9Y0Z7tQ5vsQf0bmPFaTpOtpjI
jwzvIl2gA6mKzM8kpUpmJrmPdaX2sO7lcvrnrtuvXpcACWS4HOE0NKaZXe3+wa0E5muTpx+nrkmv
aL48bVEdaNi6mwAK5TQabcv7dquTcvJQa5hfjonDnFXa265Fm89MaIzG9yx78sIBnW7I/D6KJwZO
RGeF1GDRM42QdRzhtLAosWp8WmKRQHB7Hwo0Dag8jPQvfVOzWaB86hpl2NOmtC6/mUqM9eyYQAss
8iMaf1omPPshc2tU4wWj3hGwmZBuHRP3m2eyCbJgrmA3M2LMcj8pbaFZghvTXvOEIzuLt7Psen14
cqu5M8XRWX2AtCv0idVMtqxxquIIQCVF3Zel7KCYMR4urczE3x9pQwpLsooEJdWHaKRJvl7oQfJz
igVbwEMNrJeqMId92t0+OiTKvrHMKeYbHPOIziStRBtur1e6IyaSv36suR8iWiu/zfSk8FLkFYAP
kelYmJznHBqodxz+MomtlSuCip2Sfm5W3KPCtIG+dbt2C8LPt15mkxiQuRNhBZljwKt5HdBUPna2
CiOa6yZcu4Yfdv03+t6IzHERp3z+G8Or40GQODCqzIhLh5APR4vUVqb495WJZdGjs11OidT703r3
29JT0vURlg63bZ2gWsvr63diMJE7Z3qp47x7wE8ed+8wzPOBZtlX2mLEs7PTSixs6nAwC+M0/lsO
JJqR6Swh7WHtcz5wq1m5X6osPyz80h9dMBtGmh2jE0WY3uPAHyTMlKos0MIs8/99nqSRzQhaI9ug
v7FjnyVdk21jjGQNnTadDZRWBSL4xZFKOGSkBBlddL3aqJ85hWIPbkhnM2RL+adkimNpFKHylQ+M
EON7nIHMuoJni/ca01svgc0upKrMo+YpxAt22yJiGH4QCmaSaAr168nNbdaCPEVuusdsmW2yCW4j
vGDJ5Muzc9tOvJVyLLQRNB3lJEKli+5lnXeIp10vWP6H3ihRx6dJlFf1Z/sKFdsBZcyw7RqAt2w7
6w1lbo2mSdHjBnJq5DQ0tvMbFw+7lxmRihVLbO0TwyNfUy3jAekCEs2X7sBahpq2+EgAjcD9FdW2
+uaVyngyllj7kmgIQZYhLXkn8a9/JvDozdN0YWSIHqIhnSSghd9NTuncyHFHoLyfRfl4IaC4su/P
MrVeNFb5WcNBQKLCyFahTVKn513J0r38O8SAySL9+5j6oJaY+qdL+Me3Rkuno8YLie9gt1evGwMh
AQx/ykedofE+2AC1JtroMouOBbpJTCRb8sa9/h18r/+z6MrQKY9316NRSsiLBSACkprBGMT1dINv
p1MXfy2n0bar5iCjF0SE/KIkVZFx6M/pm48GazyihYf+jHQpkl3yp3Gn35G01Ypia/+1jtOGja4y
2S8O92hrO6PcbfxDjWGGvEwM9q1HosLsmv6nMTV9M4JI7oMuaSer6qZp1Rn9j74ysRJhIWqs0B4v
Cmi9nTo9DST92e7IYlZ82tehgqVOqvOxyIFCov+xp1TBuKeHwjBMKzcjG/irLa191dNY4kNcXYcz
x1G7AQOhPq+YQRa3IC5buKKwcA4Usc52eUPEEsT4LFppj7pBTapv4AzcKfgfdU8VT6GFRwxR2VQW
nId5R428xsdgEUqmdU9qL+cNloVux95+wddcaHkp3L2e2TFoOiu5alpyn+Qqslj5hqVBWplLbVDH
96dpmbCUGjfPnnLTV2iNLd502xHpJeuVSRE2IRxFhvbdax4XXpb8JZeP0EmoFqByWJJGXUd7+wMv
J/nZVOCuITC60tZ2nk6VwksYitI4mV95Yqqi+pN1fBBxMvElbzqymgWtNarsgGIaZhuqA17FeQm7
1agM73aSZmM7SBlNolZWwb3QAApzj4Pd6o+sAdn7QjJYj/bhnzl0NN2cXNAAVcW8Dor6bikVMn7z
nVe6b1ab8G6Zr0/j28Wus0jV0ZTJnKMWG5SL8kuuftc1TONAPyY8ztg9qiTtzmfuKBTfyGJEi6r/
P3VKWZxos7OHRmFk9hOxBmx+K1HTSqXG0ykKPQj+GCMxp+wR+fcqFu9fGPgL/XJsq3vHUy50cmwf
nSbyi6e+2IILvND/WqS69GKmf/iAnjHGFK65VCdJpAGSEYgWBMpfqovnx0o0VA5ri7A5oeGUVI2Z
SzewTZrv69mevYel4jzInbHa/aAPhvqTs1CVXYM3P0wQBcwLMGx5K6f27JrOmI9q9gyXH/UkfwDX
3OIvPzUPzWPL0BwfRiioK/jKcPxQ5fkvWFXbhFUALbdsuerIfXQD/WvFIexCu1IL22vSK3wa+Oe+
MQPDh9Yw6hbM47GpYSdfU57dw2bk5MFsn7F3T84mma7SlfdtCGoqswtB5xKhPF/Rqp2AFQllepDu
/1aYqYvJHZlQITUWWHPZZd0jWQEYA6mmAAhl12+Wl0Zh/lAd9gH+1X9qyrn8JB7Ucl/+FvswQD+W
8IIwv8IpZnMZDiVBz0kxu60xqYP41Uj/9dT5GgVBX5Cex6rTemS6uiL6iBMhJNpCTN9BX9gYRH1U
Gz6jmle4YiE7wB2FYtQgCcYNdrpGHyAgcGXVYG/fo84GFu9FGO0/yfTiri7oL95B4blEFbxqvmqL
wK9IhHz64azOEeQT8jifzhrubvm2WVgmoq/XpRb+3NmtIMHGJi64Qgzxy5el0xamKevmyLtnQ/hM
HESoxpLgYGlbsXX8i7vx8oD/8p4C4anBp2E2uzLuDiRy7s1KgcHRHE22QR4oFlKA90ET6Nhzz9qR
+pMdX8I2fo0KDFDZS8xACb+FnfdvKD5GTvU5Hh0FsDtgvH85x5uydylXKBBtJCZEkeh9f2j+jxMa
hnpTnWi3ybO7N6OzVVwTCZ9aX6wcAltrXPzGghL8ZTiE2J6CPl6eUgLYb3T9x82qNMLeA/uWcjaf
sPcHsvybQLeje8QIeBbrQagKVaSgHAozxzDGoEQaQEe+w8g3Z+Bn75GjBWmCWKvLAEKjBGsagn6l
R+8l4DQbxPw4NQNz5Ci+cnM5dNmO/bGzK20a0uCEEDOEeKV3hXRDPHammzdpwd4GL7aMlpuohUuM
M6NvghZG8m0f46pSARYnfQeonCFyP9+d7euZ2kg+KXUDHX2CzQvqQh3qFLrh9oOVvANgUakBeK1h
cJlbM02oGfP9Zt2lTz3eaUxZWKNhpB1cq2W8kCyoGrUa2JRZiDdl3goPIgWCL4+o1rASdQeQw3h+
EcwXSCakGO8sK1DJIuA9PFOVq+8R6a00st5FnsLxWWv4EGIDZUObFYDTu0kOTNgaaUqufr3VJK6E
65IML78/ksI/bDmCJKI6+iFVumfEoMPJsqUmPr3XYBFeQybg1mOq8PWkbLpqyVH9eozHYgM+PU+x
k0oyjTC4OVnMqTL/R7PDAnEImPDBafZc2HWC0eLJMRyBuN+tdJAJABViJRXMjXai97XUle2qmB2U
7O0/u3+X/Yi/jpVKEG7MutMZ57yGv5QjxODw10uOlPN7QEFMKnUWCXRZCmexgUKNOzXJ53Xgjlo1
QyP1PZwXFxrPjxrNE3h5CP5sUCWncdTqGja7WYLWnJK10/kjJEcOTFiQBh6V3etZWb6s7lAoGuDK
sATRoLFes0BO/Vy6/xjhUgdYlHN6lBTVnzd6W1kAjmLRfxMEgdGNTgNwp1UT5oyPAbEVUdFmsHNG
Q4kOqwNO1qqtjouEIY6RXy+Fcjyf4QUb9PBMm3G+5GwlDuDHoO2VOkaM4Ia7Q0c6ziC9oowkif2M
D1pGdb3E0HyDZWt+PDcy1b0Pxizf8illv3lC64Ug2ON/Oa132uyu2lxB52rnx47RVy+naLgmQPRS
MAfntOMkoHUDEs1wwzMnhA30swb0sIDs+TLNQWFTjrqbAtGfQtmuQ9nzjJJki4M4nsWx/6xUdGUQ
bf9QmECSAGkqnokD4i6DIlIjIKHeuLALj0K0PopW9JQ2Xkq7LYye8O10NELP5xDv/Kb5i8TOhiri
jc+yUzlTTsVgRFgWL3iY9oICbetU39iRHslTEG6drhvmVet1PsERuNfY+sYdq5lNrdcrb+NjAi66
X9j9bToZGPACB9B8Tq/zd7bGc8ov7ONHfYnePzuf+pL8mkVwHstE0acUJMd6kVVCHLTifEDuFDzY
p2bFQ6iYdNdKbGKuR9gclfY3+eqavlLm427zvRg4LhC/eVv6ds3mW/IOCX5mXADLUvknK2lpP3hq
O4CRVtXjfc4IbzA7QxxNfcoisykpq46n3pejdqATl07XXzEafal27aUjjmusujaBDFA+U2/3s7nl
JdITd8zTywD7f6PC7QaqS7T6UyfRZmlNw9O2wQNpJeEOqtpWSgy87zEUUdLtEvk1dAnrt4aird6d
qsBsn4Ed4NmY6V4YDB+tDJOzvObJcfwpqDUSSc5GNw09yhEEBuAeq+CPjlNxoIQkxMupzWvvSh8h
5Z551mAuZ3E1Ze/QKQMGeP24wuthVRdvPU0aq9T1+NHl4tTx11MF9UM0EI3qR3wiVX8BYcyFwNQG
veawLGAj3f6gGyhMbxquSbho7wmvYNdw+SuO7o1ZThrZOJdur3rzpKwRJW/UfhE6I6X0hZhHVaSu
AC6Cvhj5J4NM5SZNLzu4CTC7pjrH7V+d79QtzgKiK+IP5TdYvqcYR4377CXjNxxTbx0X/Quo/qcU
x//hhkU4A6X50o6ZHwpWuG9SZgPtQDuMdy3YcZi3h9DLS1KtlAQ219cLTUqqmqvzIWz0DXYWhbR3
+TEHC6dRa2F5XkPKl5//jJaEQmOamQtPecfWH6gHW6EBk0ldAEzG+3jRjOdpgcjkerB2KqmFng7P
89kt7NwzX3S51w7R49KoZBxnFS2Kufq9k8DZmYcrTX4Yv6S0DswMtoM0e7/hDiKvn6fO/7/75+ny
OcrrE0lzGDfyFDDjmSYzIBcZiEblQh64C0ZTd393p02DB4TcP8iisQZwmbNziXGXU+gFp0OUA7XT
xLrB71aq3ofvpph7cmR0TnN8ukeWnKaeihU0VZxMoXsFrBhzC3yhkUq+LHLwLs/tq8DkddWwV6o3
x29+/90R1ADGjcbFc7SLHXcCBk5+8t87EBBitYda22PxqZ8SJlvVfb+gVkbFWKBBbf4nIGMDQxM4
KPgWwA0KHlkaot3Ymzoyf+v+Ou9NHOBxBnHIoj7ybPa77Z/4qgiuR2Yl5b81GMeza5hMDXLXLy83
gRj/88JtnoyMwZwtlnD72cgDb1HWffFByT448HpV6aEv1gcFdQpxWgjae2Cz87KP0vklRpFTWR//
4WTtSQftV5sBWaSzalBWB4s1uJPryeGTyjULqt9ZpNBuUGo3YCtZaRLweduiiUN8HuZqP+eQNMKf
N7FeHQspaJ7f9AUHMLmuyBvVWI7ZZ/iyezrLz+KAsp3QI4Vl4+6KBciHYZqM38aEeRkRJY0HY+OR
brCCOI83tqmQESEkuEt76nJmlYCXr2tlrTaXcNjoBEV6K4GTIQzN2nMlNFGfbe9DPoZzyX6JZlNQ
3PNcQMSR3IxkhpGO+DizBJvHT94IyAPdusZgTw5z7Pw6VVGYjzypM1ekp5EZrQdmF27lKlCL0w+o
giIbSqK6PaGSyEbavcq5aWw19D56wPCgksVCunFcJ9T8izLqwABrvHhg4XYbqJ9PyXVkMul0ubYB
C49xin145MUvODAIMbyxOJtYkJnzezDeQLhnQr7MSQlrGbk/OLjCA6hgktwxB6igyhXv3eMNcR1W
rMQ6Qh18YWg+4AVw3G5st9SG/8C9bfpU2mtAlUuKhb+EavTtHesCWEmemezS2W8C6TWvl07C8sg7
mVvkRE4HxWRLQEXrxMwpa2omVw0WJooBTFX/jfAlSzIsTLziMGlFS4YpoosxAIwxSxnTILzdgJdY
XSwKYrslOrOFu4bFPAvZ8/uA5VMRcgOozct89MoE9nmETk4ScilPZqrDO4KNsl8BHSa4d90V6QbW
wpVAVjkKzIsbNfTWs/XT1TkVyw6m5arfWUik91ML8oZr8sPdJv2xRP7D6eTkn1Kzi2hPdnWxVOLG
p98GFLvOg4XRdAb2okDmzioO1oBL59XCXR6+7sHp1otVZaUDDrnB3hOXpxU4O79vop7u1ulGT/Zi
GKbncJo9vwolJ02TPWEaNi67Nro0oUTvqcHyDHN+DkleEgDD/I0Wla/C/kIoW/yyyvcCgi5Rl/iN
glbvk4CoprzoneDpekZrTaM1ndxUqpHsCdiCGRWf96z49+hgi8TwOjudOXRsOgMjpqL/9mDx7mRg
vKwfS6PPRtp/uebvJ8OAGs8MQ3eEXJhESnAB97cxPyomjTTOS4C6koDRqXoEJ3mdgyPuOu2KNk94
XFS4pmeIFtWXjGMfH4U9TTc34iDvKe08Gqv9Rn0wxpk7VrGnOL96HKVK6yBppGyKmKK1+9cNAAbO
e/F/TJGvzf8a4k/XfTJ6ZNmQNfLcVLLaVnchJaEyYSy8n9XD77D98m1ZXux3CDxhIVues93vBjka
t65yfK6H/5vuoZtmhOq8Jb3gKEIdWl1xjbgKZjVs1S9XHCQ7vUgXdwQN0fhZrlEu54YE8n/LBwlo
7A9zXgxp7w0UdwO5JIkbXy5rDxP7WAG++lE0L7ZM/pv63gtvnEmHvC53UBnLxMHy6AwmXZgD2Jn/
QkXQ2/JLJeFzjg+e2i4w83DrKTqSbic97PQSmrNCe95WeA0tGgIeQdBrzlMAVaCKmmFUWKH4Ivzu
foVZzDrBXS5txt2raVGS9MJeKAJ1LeCRJTCmcalcfN2Mco+tLB/f5nxU9Ie3IC/sUA6hzu0VbzRH
qeMxJDPEY2A6EPpo5lpWrzaRRaFjbJ5cVAUWp+oUNtLTaVSgIo44vXSZ0IxbgEZFuM6ly/OJS45q
iz2G5msJgLTl0rcY/+P6ORFbY8VS+D5AT4USD4XP/8cqhzk4V2zGqAIR5dRXtp3hE5SLGsyRY6Fh
ccehrInSKk11Mz04AHo3XdIaqw7TA5Yif+GdF7qYXaM/Mg6gNyF8Ku4QNJSImyjcafWpskRcvfF/
HJYBQ9d396BjPiVF01rZBQ3bbTm8iaeke7iyi3A3dcqS8dVkMOZVsvWoV+WwYIOgXJ0YxsvSDnFx
BoTENvx/KwFH/JcGm2WsASikBOUuZxuFyuyfzwdY7uW1Na7ybQSZmJWK4bEI5G6XYNi9O8ydYSYq
0ygdt7EQ2X4QxZd78PkzJ5mMza8v2i53iS4aBj/jLPQxYyz6BANTCXBhJIhS9pyffJc4i5iJ1CKH
+HLG1AeoHlm/3i8sP0z+WBqrR/EDEhZ0wCuZ6l8h1iEOgHEBcBixAMHbmMLklGu0Mu0gVcPy6hZr
9g7QcO18Js6LKaOe/Vf2lzrCL90GfBE171cxqvwQYnUTTP+BZg6ydID7OuBPqoi0p9mLtnccWWGg
d5qsJBJ+IwGU2HkyNuTiNyUnueoTGWHEQ1JWGAz2VeZNhsRWZWin+Mi9iEVjA6B8OoqoS9zxXafL
ceMZk/IrtBSgPr9uSJRTrx6N0AhnD8Ls7dMaky0E2dWpUMCqAu7P6wfsB5Wb4zIk3Lo4tLDZRmEA
9Uo71NWdpq/3p6gPpjkPTOT4iR1TtRlo6XugxKOsZmA90cHUDm2pL981E/YlNsuTLxKVY46v+vsL
GabirO+sI/z3S6Xsu716kRCjifWgNWtr1iIccJY+VLd8AXJ672OcO1G0Drn0OpRnAlK1VXRqLd+o
3qJUMm+k5B97StvAoa6RL3x2v0938q6c9zlESQ8Pstd+f9/n39qZNwWwCbxZEOY7BYxJET4SXvMC
N9zx/ykWgVcudpQEXErKrK5ZGVpQQge41azi7Hf5kWT3x/gbjZxrYQPd8E396Ceyu81uSt8zTX7y
6E5rwli/Z37NzbNqXGW1ybpXcYLRoPNbmIB5ZDETQWrNNkwEPARlL21Vi7oBF7vtEOTXX7iT5sov
ZoAIOQSL8cjte6hNWf1KJ51BFlr4JumJJehQj2GqpHbf7vVj9QdmsoVJomfFyfNqcQegm2DzF6Xa
X5uIc7OMtc/9og8aq3Gf8fjRUB8bG3bOUdofxvoamoebckh+9gUxVKqMBgMX3kTOSQ0sCzBob+tY
9fbRlu99b1k3Cx7EV8D3rEmQUHsiDz3WwUYRyTq820g5544X0ynoi4FI97MoyNxkjzej3wqlMJ8Q
Gk/INc3r5rvnLycjR0kzbx1OmnoOFy+H3RJe2kg+1QR9PCMmtg8Ml06/c5q4XBFEgh+6HsaOZvFD
eACfh4+fA1bgx1h9DQ4nIJ2ys2lwl3cbvzaYwWIltpJo3N2B4eZBcrULlRwvRZgZBsrDTvX4plx2
2aGpz/rELpg6qKdbG3bU+IwIXxeE1GRlcMXpK/20MDbLqpxxxDb+yfV7mIlWVrvpZRqt8mPJlTkC
OzWbzGO62vf8LP9kB0z4wEW+r8k6e4QxDgyc6Ov8ILCwRJM2xj8joGPaCY4TWn3wKdKZMtkW9uMo
VqLmvi5MmTOvwMflWsXRMvlbPBzka/9E3BHZlrvIyUo1bljkiRxji7djjr+Ei3xqejhBqln907Bl
r4CTZ2kMhfaPdMBNahczn2LKTrxUxFaBnT3hytvk1oJnMCbqrGf3mERBuCdGm4TVefW4hjpyb7Cq
RDB8hZyQFPJ0Qtm3i3WuTiaVLA5YA0Nrf5mMn5PA42IIdr+P2Pft3e7loXOoADtuFU8cgaEy09Rm
qSQeE6LsB7Bbbk5eHml79v68gUUniQaGmVbT51w+ejN9DCOxPADMzCwIrcOt+j4YsD82ng1M2OFX
dTve4NYa81SGmfqjUMdFLuFR4h81lGh1xxfxGopoK0ZJsa6rsB8Wz4EyB78J2g2H5XGq0e8pDQd1
7+dtsK9tdZgQf/bOvtMTWcpYoVb8+/O+NgmWm8hAxA3s+SLEpGBl2vh6p4K9DmEWcVMVkCXsCHLm
40eIU/F3QfY7tcRysyXbRa/CF1ViONsyUxHdhMtHO0gyfgibtrtHpzSHRiXHVMq7On4qYya1AS2z
y0RygjxNTdoNK2NJRAi6m9o5dQvTTZyws6mXHYyZWh/fqH2bZhuWcbqVWE33fxpuN3cuBXPB8sgJ
DBCTKcEb/5YnrKu+w+h4tXJVLm4SKRyAsRP1q0Q1bRHVGriwblFiMXELIOGwDyoseS10umTyP+oe
DCQaPe+qaNXMyoyg7yx0aLP7iKLYAKYd2QK8PJJKY2VleHl5n+JvdHJid8xXePo2GnbHxogIFuIB
ppoN8XmxhusWf+fV1ZlcPGs3UV0az4mP/jHLu6rYRz1By78PoDAtsXRJ++N1FjknmeR2MNONGQ7Z
1rNxMRr7+vmSCG0BwFbQt8WgeRDiPzvOYPOpF1KiZi5ZG1ECqs1tVsR7yGK+6CM5QFTZRhuJNek3
RP70kurQwnZP9UU+NNFMnv9hxAQ08P0eJffCLd8eKf4Ud/lNaawkhgbAAG1fF1ROH6sJ1egyi6t6
dYnOwhH20Lb+uzFoFVUaoLRi7rNRpSYjUQBJBGzhHn7PtVj9GXyt+MFLUYBLqm2NgcljNk7nyT+V
C6wlAvO676PcEqlQLtzhGiV0ubz0K+NxtJadWIqa1/IzG8RjN48/fBf+6xozN2bRqQEuF4yU2rGH
mm1kNDvVc/dYOqhzZ7Mg2qzx5aPRPKTb125RadgzEw4IOGXLraeUYO4VXO13pZBL3Ted8AUAPnxn
trZvdF8VwbgRtGhEuo2LTMgbh/IfPMyOhl1Dzx6bVISGIxL99XL0DJe/PmNRGd9o9dAi0cpAYje8
RAMYXqA5UKGwaH4IkYIYCcdwtOiuP5Ov0Eczd2jDXIZ5MLnSL/vD7g0FZymeOJ04d3gmV2jmPpub
hzf2qDKKxFD1OYu/Z9hItMqvrXhOZ70yH8qwSsDYid6L4FJc/BYwD8rixjOr0CM4lHPJwvQo7RIF
oua5/NxzBmlRIwmHqeqCAbWIHgrHgDUh/M7gzdhpwffdevyUPBGisVB8aCUp9FyKH1oZ5Pc7UKuf
SqeoqklM3ZYwkGMhgEY+hb75S7boccgpGeUK4sYuQKKnnd11r3L3oCoAMLGoXe8foVlz1+ba6m0q
IAiO468+gXRTQ938lajmJ4WWbmC1vlImebocGr54JZAHNc1VSGCxuZdGrF83kyCVoFXQ+JgPXhkM
UIocQ9bkssfqbxKp1ZFsbjKnbnxzvzhlYC8tS+dF5SpdUOZcuQVkyuNeIZ6J9ZoFacwpZZ8rIQnK
vb4AAy8ubeV8SoDhv023I9awCqt1PuA7joFhiI0AoYfDozJe1WO94GQ5msTQ+VYFc/884P8ERry1
AQEb13xgorVijPThDn2yDueH+LdhoM0Rm9AgZlME93j7TAUmCqkQIWYNrOUBrA1AZOwH85Nun/ur
psyn0CMxJgfphvL8MVjsk6RgzhSXPB/dkPS1g3H4cdqQdOBufgZZZfUGfpaPUAEs8AazMO0d4Yqq
u3rJnGqhktNhPOJYlMLxTTzHnh5354rwmy42VWItEWoqo2Yrr4Wc/Gf6EuLb55SFLWHDCcPxCBPZ
akZWvHpMQOaYMy2x773XJ/mAoWUUx5K36Uaxr7NHoePDDpwvcz3v5GkuhEBZ5Z4EDOwTSqdZpRvP
7brfthjgZIZOd5IAId0gnpF0rwtdOfE6WgxFlW7s+SbhLg0gwrrgZy2Aas3fKejSu8ewqY1IGCWR
KnotIYzYrOws1XW1rdCBMDWHunH8hwV4qgUq86aarpDmpjNjYfrfwDLiBi06T3eJMiHzkRqScoCm
6Oh7/Hp1QODaSaE+4dZZWvvs9Aso2O+u/gd1BSUQDFQuvBxTAhW/0lbByDX0K9uVMWL9vHc9J1YC
EGshsb537uWf2DNZnajwa9CMN8eanY01EoR7as+oNOdZipkjaFvUHyOk08/sMFOw6jjCR9OrIgVZ
/yzciC8dJ63dYQrjvPtMK29tQobYpxtdCaGt9WbvSZPGZf52Zrgqxg1YVIXv8UHzVlC/7Pcso2UU
oEY2fb9DTYceIvyp0Wa1lhhkrO+o7izb43rphoxpOPuREFVzBKDp9ToTcLn/9Ui9xLXUsdmJXLwt
ixaQxDkO8Zf32G9x476JCkbzh14HqJvAvGK67GH0G4KOIAbIhusjdN9LxJLcfThZvxzKbXoorqfX
uINxtgYtchhM43+EixFdDIXW1SIaMoTve73v+hKWuYghHgpv+8aV1F82BmQNVkTyIyRcJw2Q0GxX
fe8OmwO6FpqFm2YJo/cxvAlZnD+bXL1AgMh+B0EHhV13RcFLXe3alTs0zeOq1udx4qjRwTjnJMyZ
Z7JUIPJ7FO6x/A8AHHBKPHZkV1wsdEAouNsizSvscExDtCT9CLMj40G4qLZTdzmEAWZkBh3afPYQ
CmV6ZGTb/T1qNzVKDhJQoEE9DUf7Z6xxthkPNnfwohXgy1tomklX7YqazMsHrClRdMEmBG6ZoO4Z
h3ZzlxgdOxuSO7vCaYYRugMemJ9Q9AR7oMpMFz80fhFop571uJ6Q2kmL8F8RIkrCOJ3CJjQAjMXU
GPzl7hcHy2mGu4XFU2nBnHSDuLUEgPxM/OyHeebNmiFy6nrHhnmxbGqgsTa4JQPDEPBTpXsTdM9V
Sq/pT3YkC+1LlFnSvOqjXMHQKkrQpT4AUlIlQoqLESbaz4zjCCsnkI227FYljSzr1vwcYCQc/32L
PsLkdLKV6R2lhuJQa1pT7Jy8EL5sj2BlrUG+fgaEjAAVQ4u4L6hqgvoahNtcwhskSLhHoGlKr5VG
9xpECetpVKxWvWqqOOsjk3cJ+qh0uUaOevoMOZVjSVZTVY5ygd9nEk1kdxSJ9Px8sMfYLoPMuxkQ
RuEuq4ahSlmGgcGdXjdrmKvTvKOlUDa7IZpmFhksL9O4+z0Ncr1o04cY68wWMUKpaJinS6efRpDv
c4un1Wqqm5BQ0rDwsvrAJCSNPX9ptRaOAJAAlcEA1BJ0Yju6KPm03MHvgflo84H9HiOdF3O6m5h+
6ikCdqyCCOjYnE8Gh4kUnwz1LpjL37cPCtbiErAjvO8HFCCnQ1b1QW8BOOirXR5m4sveZE1FfXVq
8QH08TJDsytHkJPk2tRjz0c0qIVUgwfaoS8NH5+esDS4e3xVjNyOWA3PxE9/Deassxgel6BunwwS
SME8VlWOgAnYXpONsggy9XbkzmiDBMRo0k4GYlFtn+poLVIlQ/9c+Y44Ggdh4W1TYXzXp58UUx5P
9aTyAX0N+tNwJG/oSUlmh4sWmySy+/fX25YZv6ht2pnq8FgdeeVD/QdXzrpTn9CK8tim1PlTFRYY
RcOSQ8HO60UIF8/+2qhRn67nT4hisLNHGo31g9uN1Gb/u6ASeSjNqKVziwA27LZD0LI7w+0sZmKJ
kEhct5E+i1TFrhBLwB7mD7HbHGFwxFqZ5AzbzH2fisNuvsCSj/bMRbfKhLpH3FoLDbMER9TJ6dkS
m6yAaBG4BACoEM6TY7Ah9NYGk2NiF/0S33h70KS/wDe3FTo2vz7uE9GPYeug2Wnb7wj8ny5MCl1n
rPftC9ek9qV0fxClCw7WbG13Fta6pFgyjMjkzJ8AdrR7+pAYhUNrQ/iBnjF6P/ZP3N4DFXAVabe4
1Z3Vdxz6cbDL0cvtbu7hM1hTJUrST71yl0IoOuiC6J6HDHyhYhtJHJiZoLXGNSasdoaXTSk/LZ2n
a9hZsbUh1DWbpGcwbAoDfDwEj5JBgnXVcxEbukJIHG97WoKEmiIdaHPYqVqkILQmlNQFxo/zOt4K
SgUCDsPOioq//csUwbBth885/U5E8N6Je1gF9n91PgenOvD9pCQ+oyEzsS2pcLpSFUj+0++Uw8Xu
AbONTbYAEfpl5uoSzT04qYCGVNiRry2HpEFGsxPStSSPVebEcEvdlty2ZO6H48fTaBs39LdQs4ur
zAt14jSA+bpJHymo4QG0ISgONLJLgJYcVDd8aYafGkqQjGMlP4ek5pcjxIUwXcSOwdZGOZcOGJr5
bfB+vmQTLlJ8k0aloq8Ez14j2PLEQc3w491+70zI4ESb+NZ43zIpwU4gcr8EXio/D5CBT83+e8c7
1QYTLSyywNVWWm5yFhTpSE163QGWUcU/17ZeueVNzVQDhX+ygwUwSgo7CLoHenlOo/6LsX9vpFwb
5huUcNBFYbJRTggAiDxJXL4BBR8WDQ6AldGGnPy8id0elpQbKrtEi66PeRVhpS/hu3I+onAQG3uS
Zy0htTlcBQuGFDEMdMmt4J9a7Xq9FSVfiOharsjA3qjHh1twtp6x1GHqEvMUq803A7rPlefdPXQP
lzriDXCX3hZvkgvAqMH+usXQ59U+c9h59rijW/C+qd7vPFYsUCdMB2KWLfCBp/Ftds9bWs+30V8d
sc1V9tFAZvSGKO28IC5rq6xJ1CwNereHy+VmUAR3zYX9hEk6p2WtUvK0ANgCMHSjy33jrcVmHPFc
dig+T5oGYM4DNYVwzZoUxLua8MYTA376na3d2TTNWjeG/wkhtiMhYqhiBOwpE9zsOoOrOFa52BKb
NRVQ7WRlpUfaL9yO3zKyfzuFiY3qeaKTC/D4xhZpj7bLqWb9lyT+O3fJ8pkohTsMBZSCtIgmewK1
BD7GqF5hSSW2M34xDyACLFqbs6uJxsiuuavzwhap2vYqBD41UDAS30oMVlSYNcMro8PD+BktvtlZ
8VvENvgbmsGNyV71ZADHqlRwHz+C413qBNAj5KOF37qTXtrNcFiOsBdgfOjqM3nRbY2Q1/EVvjDN
k9PKApEEejpzsXX+oc2xEHDxfpmT8K0Wn/FvD9ZsZFaYFjqkRxoQGqF8f6wDYOmlmcUICEuRX/7r
yiDtAqFnV3Rnm0aVfQ4QSlPBXNcMuPQi/qi4zRYkCHVBjv1Vn56bue9uoQUQn6X6M0mIcluyTZlr
uFpDXn5fmFpC0Gb5RPQUo9AOGKChPfSZtbB+Cqz/AGKZkBdJeNerKBDye/lP4mOyXCpsI3zn7Zjw
Xrbgd/0wGTa3rp7QHpmKyBbmjKtY43MNgy15tWkh6qRWddpOUASH8iyRaUfgN0nfqXlsPLqDdlJf
H4z/GFNBylRLTI7lnKLyzXNrTCKjaZfN1DqrdPCd2fbKGZnB2apSbGMpoJ+5h5StgcG615ljEbtx
Q4/H3J/qvQ+9I0YA4kcxU2waBzJZm1TdEJJYo5cfBWIoLgpjSOXlM33nU7ro5BwD99KNlsmwTNFi
JFBy/FV5fFmISKex4+yhZOclaXN8LkyaeyI98h3ksIDVKgbm+6CHCg+5EiADzFvqhLtheEu4JBzt
oFdiyPbcPixFPZLpEPNpAJiUlqfUtzpBGWMjpBA0weA4aXjsa8iwxWhsHjgwSQaVePVvIpRCmVhw
s3FEZQnLAyxWQ7wXUPI7SOjkgqIGHS8t307WwBxD6ds7UgAjMCyhcncH4ktCuqhQ8hnkWZUCMdDk
jIWObIVgonAq5u+aBf2zQedrJGNBZOI9/irYjybY3ggBQibrxwpoDnu5ScnQkFrykIUD0jY+AS64
1HAnjHFCepFHHwdsetuMSclEoqRtjo2QmV8yHBOiQKVP+ttq6OobiRfCXGg6zb0u0pRSPysm+RuU
lkycsjansok8iDsxwEiJahAERbMN+nLJcRJZk3Jo4Co+A6nORLvs+zYNnGRV3Aw058710jPwiZWt
UGg7iCbuE+XYIf1cz9nqD1LtIXhi7RnB8avq6Vq/1G8wWOtXQQDhVPZYnD1SavqBV/UKwU3rIHVb
pRN/jP3MPbZ24Fh4gHnBU2Ptp9FcUSoh3xDhEUUYjCClAH+BP3tGGUFAKyYbDEskdwktIpGtbN2r
pOWgJuDRMkmuMP0kPVTilqW38j3t78E1jSt7mArqrtSkIiAtgQ1AomjGXYqzU7IIvZsZ05WSEABg
GPkCRjb1LQaj0SLFxd51cHBBFlcSBozCGid7qdZMfvY/p5IshSyhtZaxaGPdvcB4fHbBioUkSI7/
Q8XWaJlGN0ZjQBvmvM/olKlpLEU/6ZjfoS3YKRDCNZbDRdlLmBDZXmO/JMcs94OXP1IgYJEWE8Xy
9dg4vIJ3eMXH5YLINuVUbBlX3Qu/9F6R2IjgFfKbGYMyvM4EKSy7fusEK3bP1Yyqf7MDdhs3m3R+
yjED0zKBcEiE70pnHqM72UAsghGvGQ381KjG4m6b5R2oNT9/YEv6gh3nIexZ8rpqFs/1FiAQzW6G
WhVj9FNJVitqhQbFl4wdm68Ex+vQSIld36rwaLV/jnjmqIteuvxzN7vW4e1FEL3ed41r8UURM+rB
hFeAytjHwvMuKP+dansP1atLCFwn03QuiMifaIqRzNg+ycIviNkZHGomiUZ3zjfb9QHrtCnL0Dbb
4VNqleUe3LQWezA1MkN5AefHOnjfGoY9a/+8BM+7nccYR+q0g6qosBYn+hqQibOblNKB+JN992k0
VMUgaxQUXNToWcpZiwM/cpOi/NJMwWCD9fUGJfzXJl3FzayrWRLPpciol5Ajm1+8hMupqJNYcOvN
TvSknAfG3lyHpkp153mVZl2WuB/4qFHH91iuC8zWBz1iq81JxlJaeSjMP42jIGGEt8ny3ftqLGBC
XvGDimEr99BKQtdH5jIgZjq9Bxw3QRcYvAJJ/TmjwzeH0L8SOvXw2U38towXdqaZSzERrL4smo5+
PlN8p9YRqKG+zfMUy7aiakw75iUJ1mfl9DyHQrLXH8dTNiMrZTOyR5OO7+GOQI8p5b8vZRTtgayw
uegkmmG3yQly1/uEBqcmMEg4u3ldz5QZLtysOJ030K+etzrQpVvghoWN3ImP1b/A9ULFf37KIRuC
K/+x5fOnDYVqN9B3JVfWeX+TcN7Nw8ZlInck0+l5c/mGNYhYWpNvC4qTrCMSxbpuK8ASvA1evkpt
9U7SLNU5z2PIPKk6yO7IfvacSsmuff2BJKEv01o7jWVy7SGAPk8iDJaYbZxJ7w9wvPqKySQisXIE
6zBY61B7wgE0+kO4FuvSMLEbiBc44Qu0KgFPJDS/irr+uWeawj8QOoSfyy1fk4QUHZKV5MG0Sa/r
pZWgBJncCHi9zMMr3tX6KtWYVPDlIRydiM84gbIylTnFrka1HNRbf3BFXEaELw0XEW5lKq6NtZTY
N+7z27oSiPaBhvVB3T8rSodI7BoTkwBM3ziyh5j2DL7KVaj2pWwwHQFy25QUOY4LGGCRyCBeUIb8
3AabY5n06SqE022X+AKSpuf3zDSzEA/dykGBCA52Hgs0vzcUZBXH2/IIJ4FSaD3oHCEZVUNRaviU
cUT/P7p/zHZaYWOwHTZQTms9fiQ2B7RI4Fzf0Ko+BZsKAwQxhELpB6dU8WrMhIu/tzjvpmIUHKfP
l2VOiu6tHVT3A1a89+Sl/H1swvGOUr4IEPznyodZ8P0WIhHuL4oQl+y+JzNf0E1HqzNTvYWbIBRM
/gc19eYdjAjryNIcokkQjyRQGbDcIJT5QOYfAmqzuzXrr/0RRQ3nzUU8EMiaq9d+fseVj7rl0RY0
FsveP7yH2VVtR2DPRCJmTcW4XFiork2FvHFTJqF4tfJnUbSIsYNJiU7uc5HDFF9XEgQuImdFHT1x
1saQ6DmvIdib4jerpdQu/Yw03viJdaG+nWCRaNcIkdkOIA0cSGNy/MGh6UeQJzOvTO6z8nff3++t
ZgDGlKKngOcqrhiaMTbyGe/3TlfjyYxAsmXUKk8UFERRvI9EMmEh1xJogxkmE+DpqySRbvH5gPZS
WpCn2d7J5aOriZjkvkTyrufoEgjlAWZwuc3x2NSsMepPdAbQnjPPIxMj1//L+jASc1V+Iv416B+Z
x8WDDuauvtQLKCkNUxe4Ior75FOOS+vCtWsJdxPGFAUaiWuYygK2+cUzjjAiNHbKr3PWY1r9/zBz
BQbRcVUQAKtIH12/JL1lDRFDHpTC4fJWzWBLOaob/lvVVLtM9f9ZZMMqq5yp4e7WyBZEvLmWmmiJ
sKc0RXhJjh0/e/ddI0lRvdwGZT6Gg5e871Oov00ALwVF++NsYzSLr4IXidEx8YqPM+tOl2MVfyFq
5bMkU7fPjePR9ACY4FnWHJtL68NmwLa+wnezvL7T0G30RHeMILLNhaFHOhjGHEN3zCV8RJvkqtmd
O5qBeUk+J49UIuyqXTcbltBIlSD7MolgwpXOXaMOjUc1uj3fi/KUBo7piKAS//EwOaQbksIM97Pg
uGHa+EE0/IAoS3ndJmaBTu9FY8X4TI3sx27lj6KHMxiZWqfW1mbDOiOaZabnS7r35Xpvlkvo+v8G
OB0l8POlE/HOdyABvCjfoFIAGYS8vEVO/ijOtWnI5NRLemv+9hw0Hge+wOzoHK+Iqr7q2MdTVJZ7
UP9bAybkyrcMw6FXHsxSMmwZw4hHbr/sNtOrWfn0maRqCg6c7BmRNgnypwsk3xk0hSIJGtl+L2VW
8hDJK2ArqDRP6APGKGObu8ZhH0rprfkMih6ICicQfseWCzAV7oqdy7q1rsL1rwFsIdVH8zqJ+Ufn
S932EjCJ2/65MNQ/hBJdokUDhuNibzDDMyGwbxFqU8H5l0xQSH7bOdM/PYJA3I9mnb0mghLgniyw
qCzrTJJeuSvWYMz4yHCOdR+//7qRnJfXcqejbx1FC1UWB7SNU48BYhF9ct5gZ4ovtQOgoUZhJZwr
ajknTsfpD4JgrCLXaVHUv6YWh3NMaa001isvw0+6U/384zpattbcZcKiFiYHdPXLVxEUxnb8ph+D
Bhj0Pt9TyWDEdONdTF6p1AKNkJiPTON7AXBl5WiGxtu1DKBaZiVq9xpsWBVMrUM48QbHA14nAEaJ
GXvDjXqX6ZE3Sb5m+N4YCWa2iMCa0jeN14yuYXIPH/Ses4id8TVFBgac+Kn0+Ps+lHmSA/w0tHi4
owp8xsZIHfvTq6fi2WY8hSDVJMfqfMNPEXOVkHrZEU6vd7vFlKawgaSESvTWUruxirHXy9b77t5b
slQP6Cs0Bxf8G2Bgh30QV58EGRyoX6ft/QjMdycZe3BgODsHND+nC1zuJRbQ0wA7fIA2Qqe8Z6r3
8qQ6EWmHrz+QxvnKGDdAU2Cd9BIZkYV/v9AQ3tm9h5pa2LMk9+IeGIRy2hoCmgX7y/Kixsxd9YNu
iNZHtHXAjHyXQjyfX6Ya27C4LBzB4tWDaJ6KzJ3VKDPQXxAhjXjsz3EgE/rxijd3bVyWyq53Le4f
qXyzOyDbaOLGFMTIP6WZT5KULvW2xJeIMIyzCND6cl0c18Xx5QtGp+rADLRaqfeYMVVALzptcqV0
dXvpJHB7Bl2lYFBjWZjsMGGhYnZjE37O1ZUyo37YSXXYUoazMJcLk2qBk1nufZq83UV8PyLMfAE5
MCbIFhHqXXBThqTHZ6uBDR554JUixSdVV3MHi7OIJQdXJ6xygrYaXiOutT81ceyvRskAQLxFicd7
5qvqqARWIdcKtg77vOsRoRp4nSidQB3bVx81PclIJGz72jOjrH5wbh6aQMWOd2C8xJI8QIGWvURz
H2isl/UrZ8Vnz13L5kZf902n5TGrWnQV8DzJ4tPidR39YGpgNeswcB/x+gIMuwMH73CottC5VOfW
Iu71o9hQqGBZWxwlkS86mGySkM4Pe7fbQKHKM3yfubeNVfbgbTjm4Mr6UsITrwwA+js3OhdEJPzf
CsvWVkos9FqbiReAXCW5omnom0bxiwr1E2yUVfc+HuaWmA5YebcyyQk0E76mJbtWU3nkm5SxiAiB
lntIcEyMJHAw4CTft4ASL+jc4Qdb++Sciz6WTUfDgWRg6/Bhg9bhRDX/XAm7O6QHVkhB/61rPt2C
ttaejUcmTKL75llDkwCoxBQOshb+6U/bAnO14Sb9doKJg3NbxsxXfppgkiRz5vZxnY44skVWnuLl
87FcMK635phA5It1WV0vHKFTE29Jhno3V+MQJoaRQTkRdqhZ6QgkTcZCrQ05O3pEz5dbAlfotkqD
BWYGfehjDRxm3OesVpI/SByWlEduZUMkhXRrZJV+SfvV0drn1J/nSKCNXnx/+u6dL2hT9IzI92Z9
Kfk5zAPZ5Cj3lF88nG3d4a68RTU0A0OBuWm30Iu+scTw+HfdO3fJdOXvfv5y0/sMjZcQTvq97tfT
AT9oQJHr+XIZEeu3G46VWUjtOdXyaziw7f6C88q719QcLdUq9rdIsvITwnh4Xbl7V7dMaXUnTOaZ
TsqDzDGowq+p7EihJb4buAjWj6DYI49xOnVTknqVYOB1lX4cv08YeeW8qpwqyBUfq6+ellIh2Q3x
tSQbNUuWxBH8gxu82IfDSywf85ZxKnvC0sbaUWMWe0pMlA1JFgFAiiGlGjGRTMVRDEI7VOPPgZG4
n6nfHj3aZzFz+pwQxbVn0KwvkgERSpIy65vZf7b0mvL1lak8YWMKiQv3SvObZVDSbDsXE/awzc7W
wKJobPEZHn7fBwso+7lhbrIwukstGQXNpBsCNVeJDKeTk5yDan/bocfqeeYUMY4VXnA9iOITo6yx
VQsqhLDSK+ACWZKJX1FGYaLDJ6GyAuBae7KxCxiKuSV+ZWh4kIjHONN6S/Pl4PX5Ncd4lAWTnrBu
N49sRS2BUp52RHxO+RcF3VWS86GFYlxWPJYTluInciReFZx+mYFV7fsWTTGHdo2vxuygQ2rwjWik
cgYisW892T6CYrOqrHucAFqH8BaV2usnCBL3t5G/QdxHAuPCAGxe/iMd9kC2YHZN03c3r61WdbFL
lcoukSbbyURQn3o0qWZpr0KCPwPXUV8UgcX7yVHTIs66gyK66/8jq4/16XVWbUbDwJNesHrN1LQU
eeyNKXkvoXafgK8IW5StC4MwidcyU73gI1DCl93LgYRUE3RQMiWzvW+tbs6udGtYN9I6zPr9jMmG
cqeofJxBsTyXNFRf7QfiBeS+h0FTjtN9Zt876Y5H6TLcinyM8UvixQSRRq9Coh+so2gkdLuWyvrM
/wO8EoLt8DFW75fGzRi/vSDOHU9pibF4d9s+xWaiL7ju5WfUuRzyd04GRwvseA0R7LNXEyzoWRIT
DTcXEgLBDITaYnTB81gA2HOoKbgFe0ly7k1WaoFNMjV1VZrCygi9/dk7tMulYpahGkf42IogFGS3
oWGLGOyrd+wDswp8pFRnUo3asQgtt1D0Wb3tCCvA1XB20VF8R6znSEY56lPqZv95yJbaRs5ZaB8x
cBYuv8CQJN2JTroQbVj2K9ble38mtQRsviImGh627WYNBoalAdEEQPbj4MWsZPWT8Sa8/4G+L/Qi
1ABUzrL1Z4tQlPnGMGyKmZ8sizt+RN0QXlbt+i5GFBLW5veUqs+FNaQ2b5wGaS2dVQVSSCm+Jxjy
pl10FzFGi7EELBAIJNNyeKZWrrPm/jXzOi4WLq8XmyFGVCj4x/omp+sX16xiFZll6taJBxG7xb09
dyeOWr4X2S0wmKrcqZDSaiqaMDaCH86uIwlmydKin7Ul6hK28DiUpLnhebgQ9A/RmSlXw5yDLS2+
Q1OdKhZoa6oHXL5pxXP/OrkceYlas0QjTELChsztdQJhNKwI3K4havC3rsMBz1K4AyYP9viIKnG1
K8iAOhT98Xth4EXEZkzJdArJRg66IVgd2SNjQdZw6DOuhFYwJddcXlstPrSJYvk4bQXnP9vxQ6Y+
dAoEiGytWjrKagBWrcSDWyCu1hnnPxRs1ASDgpW+fXFY0klaVcIrjjZnrXWoAsPc59N5tOtFW2s5
RmlFIOd9SUuALQ7oco4C4LFSY6QjLOI8NAb27xE0UKCp60eVTw20OBIAmBVXnOmHciopLhMcgvYi
8B4DO78r2S58ycSN2kxZ9WWJNpLg6uT+iPuDZNPV/YW7E7KV2Nq4RB+CdOUizZxPEJKkkbArn+we
VKN5Ih0Ru8HPwseyj4qPI/5aFRq57yOrBlgiVXeP6hiMXUYe2uh86pAsg0yP/oudqQm82kAFR0NX
kZxvL8/u/2czeov7hn9fk/g5M0VBPiTghQp/qzmuBU7hkNb8EesFqKSqcsJ5JfwQsftAolhQfVXI
Q1PREqqNeoU4SKsDum2SFZNRht7Hu7xcdt6Kr/e0bhnlsyBcgXlKrz/q1iFs6EsupLB3pzrDGuvN
YBAWI33HlGOyLXZW0DMr/2Uu4i+geuqjvMLnegIhME1QdBM/FF5rsb1aokFqN8r7abfXO20irIfI
ZN3jkOUgAWN/FWTIbqCv+g1M+1jQ33KwI43Rz16lqkHBN0E//1zo3/RtxEDzioAFisfAXPJCPY5/
jkXsEL4/nCVFXYHGQnzfQguIM6qiSG6ovBrR2FnAFoqpBaHsmCZLo5IYSOrmS+5ZeAyoDle/2Plr
Q180IPVffGE76Xl2ihJHQGMGQcga/qdIf09sE9saW4wfm/BYMLusCF4ewZ22fKJFNifEnkY7qHew
cKv7m2ho6EIQVS0hWNaHN5+2ZFTF+2vwWBQx1A0kHUXqmukN5ohL7vtko6DZ2jhcPy64nEcIUzT2
JV/zKESUHP9Y03tBsnuYxrxr6Oyd0fPDp2h9O8lxQvwrvRQfZQfM9Dv4o9SYhQAKGfyQoooZMEW9
TG235HA6g9WQtB+P8MLCqpLD8zKKhc2z+KZOJ6FVl/wIUI6Gix2aAe46s8M0XOu1a2VcNJYn13NQ
yMV+8+cOvBXBnCaXnucpjATvCJXVGi3Tw/ICjsvGKiNqV3DPQdKArRWqZ8YXzjkhgR6b/GKWMp4Q
jfjizH06OEaEL/KNvPd0x7ZrmZKmcfKPtIldJhRUNl3cftJ1OvQ5slrh64G3xgV+I/kfDhpqdiif
RnZoGXQJ2xL+NC7PHB9ZAaVWkmT8mwXSXDT8wQSXz3KYu3Q5L7/Ji8C7IcCQprjt8+7rtekBNb1U
L/JWcRbbrBbygcGhsAqmjeCZqUv1MsrHLsjIUx8gepMCYTtPrwze9LcwoLa6bwCvs9FHVRS0fx6s
49cnkOuv0R7Vo7a0wn8Ub+rMc0rI0PKvcg294BQRKjenrVpNKxn5iO7Aa7uoEHGF9AJmawE+bSQx
MdqhlG1P7C2uRINGdWzmdrORGmtwCX+QwKMOvA7ghj3MwTdyHk2lXzBWV76AkUx3mczpVf648q4B
I6Jy4ZjIqgE06nqplPDYrdbPIxygR6d2KfCs2YdN7VNne1GK398jjkrDwMRR6Sx0wjkri2K7RSvf
3AE6/a9q7SfG1Qj9P6FDbXClcVc1zFDxdQqSS3tM/YI3IGn0pJxqRSDcj/iPFlAGAAa2BaK+4eZM
OY9MfTjzOxmcw8lCESciavQwZ49YowNi4FCJdexWqcPOaOAEU7BoFfZDimXSFIGrJzJhn8AHIGHJ
Rc7te64oLaMKKLls2ss86e3kWXiu+uzsvr9XAU3lK9CzZmmYhHXKrpeJxdatKg+Gq6mgsecLY0/x
VRrlbFEy/96IuxdRVaY4K7V2h47D1/JaZySjhsxUUD9SxdglqSP7RNsjYiIoOcd7QHkrsY9Cu28K
F8uG6JXGAtvGjrqWvRzuL/9mosut9GnDFNhRVdlD5/0tu1Zqn6K3nWX4FYTlO/oI2oja0J3+ejMd
VgamYj/CgvV3Lj51Sap57Zc8hcazHWixBkUi0tBf5CIAQirRUm0lxNSh4jdxmObko8FqCZHOUokp
dxxkNhtvQEZp4VlTUG28UThkwpbETQkM6CRHa5//ITM+jcLF8fI2ivAxireL8YQB2SI9G7YFI3lO
Mld075XlkOyBa62gvxBxk6ZkoE1ojnJZMzrAq94AgmnaV7fYJCUYSXKTZ1gkKmEONDaqaIb1DOZI
i1EoNRggEKexM8nKS9ZODP3JAwQg8Ex2TFGTXKvGkYdVJoFBXYdnip44C4qpX+dOtYuKkYueYljQ
SY9ci0xFtEeiOMuWehRk6XW4KCSdBKLobGBEVxt8255OYci/kHpg5TE9Et17LhMAKRYWPTV3ijzb
ySGgATHBjW3uNrjhS+wEe0THCkoQMPCrnGMNpvukGHwCcpVUK84PnlEwqUY76ub99JNZaXsJ1CIq
FGUyBDFS/p8DU/u4WzGJV/Lgi91ZnvY+6ssqww/NMixS/nK3JtgjB2LZC9gOsO4FPrMEgQoGMMvn
aoLxlPjOSd0QYANPwHCrSBqbyu2YFRm6NgRjL2uIBp6DICucO/pZhwSMIqrHG8iAeZ66gozYbQSw
LutUwhe2+WVXHWMI/DCj7GRIfLZxUBcZF4aCGkQcRHKg5bJGNaPX4UUL/Uxjhp9ZrteTTVEzPoLg
ELnUmjYxxZijXtstZykztdX8HoFiHeAOhX0/850csHc066gP2GBiNE9Q/U8zPsx/5tN/mq11p7V9
VeIPLe0Db2Aviep5fsm2LvBoJGhltFNvWRH0ffjAiWc3R1CM/ezh1j01ILWH4Fw5VjSHc1uhCmAI
ANNotvd9zXb/ysl8o+hUPn4Ci27sn3qW+ZYDz7GHlcHBDqNkjOmdScqIejn5nlYFWnMHumYvVu8Q
IhplDhsY/ZWRS0zGf0CNbkm2d9oaEQdgdaGXrlI/+iotSf1BLadI8Po76fNL9T33mHnDvZlNloza
5p2Wby5kWq3zz9Q+y+R9BsILZrl7U3xirrfSU7Pb+CXTxjOGuaDVHdYUZOPbDaKplYVyqp5s+t1y
ubVtBMSk1MbvyOeaIZAV5Qp4W19kkjkI5OcudyYsf8n8AkE5B0y0S2/wtPIeNctV8gZ2i6+QrDTU
YJT/r9s+0iZavgg4ULN3/AXPcxzPpUlPu1E0oe6Jgxe7RnSaYioGkULMbCh25FWmcNRrdiCJNOAx
wk2vSaRYGDReukSTvq7Cpx2ZBhQntl7JKQksZ28Zskc3K9wRVQDm/Za2LN5d+hkziPaMEpSZC0gP
VnJ/d1U282cliB93t44DHlXVPYAU2A6+lbyX2YmQeyk75HU5kmF7F4HpaOKxCt+QDG3lVjwsPcjd
QU9EM6+p3HZWSFxU9Wub2WKsnmPFQ0s81UIghuxWU5Vs/ZpifsvUZQCzsy3LmqMpDafKQvdfto2R
net0kta7EpLc2ix+LbWwwc5saHDXe4fCVZw0OdDn3eMFBqOCBDw0C7wGESkIMODFjWg6jktawGae
ZimoTCGnTrD0TylHIXaSoioSJ5qDBJdTj2tFllcUmF/X+LZrX/ENuhLsMrkZQYyrDxZSmu11uk5d
oqWTaoZqBz85nYKVdiPnJr/oqfbNZg1B0qCHcZTcWYCXLMqiBAgMmVf0CuTbk4MeP9JJRyNBcqAt
P66Swr4xNgtA9gr0ccCQBdEFowf1Db9402SHylbP34ZsBEdI3vmSqESz/3/YH30mSe8lKqgStbbE
lO0fZUcxNCL7OTtLz0Mrr5v6mYS4mWTXgz3IsncrM/sRaCswvwv/U31/y/xPUr+Fyo6Ku4YiWg+f
pIW48Lzv9jdw3w3bDGe7m9aUCFDC5Gjzq68APuQSlCH+ctF9FyEM5oa3VOQa63wyI8daPQN8L4Ut
hCKf3qJ5cj1gJyLY5Egup6AfM2K7jdpUethNkGm3vMgCgqqb7pD5HJ58UVm7JC7BSPwvRlKplRSi
KcsLLrv3oB7BP9PlNvqY0Vkhdr3HgdbMWwP3RdLmbtfti2E57fZkeRezrHeZQVVjGSUnCMDOPj3z
4N4alaqaNuZf+4YUeSuLAdEJUDVKDvWa5IEbpYBG7JxkL1uFHmgmd3k1li2RIsiez8x8akgMcr4Y
aQAHDPcXEIjt3aa1lMKBvNNXLxa+Xx/WgNFUX+x5QZy9yt9Z5ZcC4qbKsZeH6SBvIgjUwhMMpxzN
RV7qFphjaPutp5T9FY2l2skmznAwBPA9IjhUkdOHv6pjjiYe6jZarbdh50C+zBD3l8XZn3ZBr55d
i939/dZI/Iqq3FQ1v1C1a21BTGhonoudR2zj0dhfvJ0aeDro+WUEeqlog/J/aPN6hGD9tFtIL2nE
MI/sYh3ca6gPj/Dl1EG/oSLmKIj+zGnDyBqzo+wifFJ9/zT7MTE6+04VZy+D5sUmn2/ySGOx78wl
BHkbuZb1MAS/7FXXt9puKApQL153ZAbwpJQ8p5a0NzC9KJrm+w+nWyu1bgV8pRx3UsdTDRXLGWUO
h11tWlGxbunxFmfApWm2Vhuza8SckcWYt6P5YYrgF9mM4qNL5UpzNOkrfCKpxL7KwmWz5CyUwT6u
JmiVzjnZnzwvyIo040J+J102JqLvTMMxjBNc5+yoPF203hP0rtsr77J9vbPR9HeOlkjSPrGFVVn+
/aqG9+GuK5XOnknUCauAzuYa41Hsgvx3MGZc8lLzmJZTjr/enCp++mA5juZ/wPIflJBzA2J/GfWx
jc91jpGQO+2I/R7m96D+lDeYfGaJRmdyses10rQ3EqlVDIaSmjFf/i+DS7oEvuV0VFgXKEQt3ACL
ODNN23GexLNLFwnG/PzMwUko9JAExnAM9+YBBM6o1C4X9g7UBmzEQDsue3QN88+N44mZg5ZkYUcd
bmpF7PDxCPuwwRD6D2pQM7A0ir8jS1k1d3VKG8imHOSBUY1LJ9hM5VusG4z9h665urMHbEbl3BC9
SU3FmcR/tty0cSb1But6jwV0FMnSl8cOVhiZUUnHTCpRGOMXDLbYZLY1hiCn6Sk4H9f+V17eqKwm
gg20Tiy/xCaZvvq1BjKMnY/9yVd/WMW6CixqVBCXyBVkcXMVi7UUTSlz4ZNwOYx+qW9/n+r8nnvI
Y87ZdefZ6pJcKz1oE0jWxAiGwrvT7aoNozzDsk59MQB6yn2u9mDs93kaXkd3qJuhbFgi+3j+j9sy
JmspHAarj3Z7nNWFLKE6PimS8JokjjiWwNH7Fo68u0VO65G5rFg7klDiEalD+WPPgXqtMM+9926u
89ysggjI5kXd0roP07Pp0SOm5MK8rO2HaWKZwEZ7+65rBiMuzXWriEba+Y4dHDYu3iJrkSy+PFwA
Hk87qnPJfQe0T7Vz/8WIdIfwiVEJBNUale6xTFQMRANuVEvHK+06N52LdgP2AMgcg3mVWfrZyyK2
QY1P/mVYA62vNA8fb/cqrM68b723yOhpb4FQv8g6z+1A5xNvbMwgKov9dByMsJMpceKyd6iNsbzk
e0fXZ1Gm+BnpDZZivu9b3uwDhGt+ckrBGFkhMzh/WF4ZO70ScbzHXJ3yC5hri55pvC09F0FENRlo
eF1Qlxm5/Crv5Zz8QCEizm0RorxScRWxd3bJbUlujWomDZVWHzdtcG2b0EOuUgSJ/DNiwt7FPikb
BAr7/MQrSwmy/eTl5P4x4pvULZvG0F9Q2fc26mn8V91S3dtPj0v1haIDIUck9o456synUAvHbH9u
LLHCAZ3kaMJN6V1d7Xk0s/tAs0EINTJm7leHZNNbCtGVBmpnbPYS85X5kjz9Hvq5/BsEtUjby/zh
vxB60gHthbvSy2ArtgFG6HXOv5/V+FXe+Ja/ZxdmO0bOKtRgt4sOj3h480MptVt2TfPnAKdDK66V
rVnBitNZ/f9G9i3mDDK4GejG3AlVXsYIU0ECa3v4Tz8RZA0WJp4fTB3AVxFBq39VYiaQwFUioFXx
1/ZQknb5c9gunGkCUgD08JysBJ+XS8poqi1I4HoOSPSFlFVfogE3oeHPqYwcq9Alsz0G+RpwSY44
ilf9eFudxYZIZLcYxkCATqYDOF4g5MSOPcfQutSnpawoIgP3u88S9uyopi5qv/TEeOASVdqfwHP6
/GpE7/qfuTcwW1b7G7MLYS19NddSE03j8xwcgkDa98r2WPl3AyfmlLEpA2rGWKnPWa3tC63NExZp
NZrkHG4a8w5SmkxWZ1YwuDnz7/z06+XsyPe1YavrdBhyZVpqeVR9QDm68taB2cANEmRTFQf0yuc/
Rkba8bWDETmau78xgHp7JgKXsVYtpc+KhjSmRcQO+uevbNOYdoJfDWV3f8noASx9dXFPPuNvvGsZ
vvGfziVfBSwG7ecAnSmOtg5koofMVbr9b2lN7g9uehNk6+FJOooJbpdCqzekz0ZatAgj1FJHmsoE
RlFxnJ0I60UGN4f+6UUP7olgc3VvBmCfr67l9aAjdpWmQr2Oe2/+3AQ9vWO088cRA2Fm3mE1D0sH
GUleetIO1Oo+ZVd01Fnka2EyG0LSrb0ZLMrHo4DyXivO+yWE9o445KHLr0cMh6dOqTeXfIgW97mb
5OBtFfpxoKgpLD2n10aE1rLT6vfxtO7UHm3ao1E/uraLCtjg21o18pC9ksszf+V/WkAInNXHMqba
d197bALKkUcxkr+AG4xSN48j5zK3cLhlf/+QuYFJ4A6UAbhJIA/X80GTc3YMWMF9tEDC3CFHCZ0a
6FJVeyYXs+ioh0n6zuhhm1hYGCKjKIngDV/l3UiYQ0BMRBz/cPTZW6jLcuUPxBd/SbmFqWJDHxQ+
kVAkDzrGr2OgYVRGuH5SseyDpXSmEX4StMiQFQmx3loVv4N/RNxbTQyDHBvVM1EQNix0erBPd6TA
2g00pWV6z9zXtgRND4buG8WqLcVn6GDu+Rm6ejLelIgDfvFvtfJEVE0n0uXFBTkp+d577s261N/K
HeE7frYjYVQWJV9i/UoJKWrSqOhWZVPK89Qd2hcJbgtNh8Wlo8IR+gz5ylX7nfcGN8vkANd30peQ
NHRrAXMu2Stk9Taj6oxJmBmBh6B0ir6hNgH0AukfX96VQeqwT8pULzu+pOtMxetcBC5Zhwv2xiAK
XEZl6tMytOcrVDSaW+m0zU5L02JeLvxH2dWQfOaByvpqfxm8OhcrwlMZ5yj3Nj8fsDXgig+Q3gNM
nxF1ZE9h1rXz6ai9VcmTIQSN3bfZjhpELZ2c2aJ05IIsgtQWViR5eg0Jle+fqSEEtQDUespTLHgh
lwID294OEduPPP4lS5AGS/XlbsCDxFWeN5sqNdX1Lk14Z3iXxZn69CJ09tUiPnybmNv5vNg7AZdI
WkS3LWObcHyWe2xxdiKM53QqN1+FbXPYT4reyBHFOYfh6sHVhs7Qim3F43YCGEckKmbhbN2WCoVu
gJsyoiN+IkmyzijEQG1C7IPN+2GDKkugo1SS/2PjBhkRJlmsRhpJ6ax6ONycC0xKwSyTKqkNAe+x
FFxuEq0dbP7Emo1xmmjngWbNML4THWar4t3h9Pm50X+9iQaD7Ic88yUUCyxmydNTnKp5HJE1RB44
9oo4weo5AAZHz2tKnflQvqbOzRtePGqVvfeUXhmhxsO88bEcsFVxiDQOG2ueqI6++Iv9N9hKd7XC
7rpA8UOcLhV75670GMarWhMjKiPX3CQAb8Zm1J8G18ErGQ3+wj/yxTj25t4o66hFeSRKC0KvMSyV
sVm4mErJ0hae7PnT0ctn8FLcCxEixup5fdsucmt5JNgHS9pNi4hv+ZOdGm8uZyDezg3XHpJ6pIxE
LHzQ8sh40AnhKuzIdGo8yH5xWJvUo83jZowyXjCAkoivCceIglyCrBRrRL1U2ubHrYD1mmnV+/7V
CY4nUvpEDCN8ABcY1E5wDOJ2M4XFSqvQyxhmT1JEpjCfCnMc/65j1FfLAm8wK3nXbhaNOXYZNgDK
IaGufR6HHhh7oSep26868Lrwk6YQcCOekVBI1mbmyrNJDLWGs1/AUnXxJ3EjW/GxEdOieqLtMO9i
js4BWkBHp4k8R73Q3hknX5v6R1G81YM1Jh4kVS5NzttLXUY77pUbCJaQ2ATT4qPk7X7iVLPM7up0
zZCQpk62i1fcSwtGZ37RDpaIrbTE0aQHvFYi6gm/5jICmo6Aeo0cwbGSOYN4D57LzdPPhysECB12
Urm0uDmJxB+xaxqclFPWawIAw8++o1EJfFE2Q3ttK7s8FlZM/yKeZrWwlUml5kWI2/QLyM40tQ5A
P2MXeTTJCJZdctQFQwKrjBCQ1liiJi24NkeKy94RtQpdQGnh2KPZR6vkaMfi5MTGd1fdLdeMx514
47nmss/jor9opNUwvm0tn86SDekvwIJ+kZwXdPz5fAaogYRmPWXmcLS5sehiUl/VUHwppwMAvzKl
NzV/iqsxeDHHTnfadu7g3BPwoEh9iXlLbcT+Urz6Mrh+F1VVa7OgcCi2EZVAO5RZAjqGk8GaRPg4
6waVulNYdiOVNtvwjyZUJdMIQA++hFnC8EPapn0092Fn7n8X/ELrWUBeO4j3yQCpwk68qc3judIN
El8zgC9K7h8TRK5m/oL9RZhikdC/XZ87g6AtEiMoHw7I8lhrBT+GoOSRSrcm8wGdpQ6R6LWTMOol
OGsrq4mvtkR/Vhc9IwWMpZAnuuoDEPRl/8SGJFgPGx1tff3OssL0pqmJkW5nhkPqojXUr3ndCmgw
nAWNTuAbHlLTEQUgXPcIAXLKANlEu8QaXe/UcYlxJ9vEEKnqk/mjDv1qmoAkY1d5d7nuLAJtMr9A
KQGaBZbU/I+cDh4orNn+7GMFkdRC8QYCYJiZj+9BU2HjgPCd86lVtkYSmQnl6Fokje/dCqET7KrK
wcQ2TSddfhx2/hySeYGRSJF7Uu7iQO9DjVVE266gzDTWPnVt0kE2Yhh5KqfSSwJOrqV7lKIMsW1I
xbKwFcvC392t5ZIag2liPfa4NhUJW92/aIa+kfl6yJjEX4WkmFM9Xewl2hoAxBIjeMy7kKk2sGX1
kLKr5iSt0Jb2oE8uRMEK9ZUtY8nN+/z9kC4MizByFgnpwKHYJuitJmITsmlFBpn0DfX1bQOMlQyf
J3O4AFJw1twza/rA6iKD2FlRVENK5RP4JV5AAAo80ky32/zpNxYCn4yoBqsg2e5M08WlMFet/zEM
0eVs4bwTTDEHT1aj4up8u1Kl38MiDRQXB80Bsw9EKJ3McyksokhMLDTkSgJZDTFoNrEjV8me9401
0NB1Yc1VhoEQAi3gJp9LCBIp9s5yhHD8L0HFFZLQ3rbzi7H783tft5yriy1Cap4rCI81yXWqYaHY
VK0Z9qYPdiDeaZC6YW4jyyQoAFPL+jWmXuhpg00F9LiR15/GDXShNHJE4sLnw70JNlfiVK3CrLhR
iOv1pJttjEbySoGIhCjWaq8tT1vI5Wv7IZOMXgMrZmtegGBSMjcffXl/4UXWKL9iiSMdxtrv9L1W
0480NolviRlxEwXw6uaxLs5XCVbH55XftBdylLd9bY0kTJmLd5M7z0zzjGscW9TYO8RLyul+XT/j
rUQyA9RviD7VI43JgreoJJgeoU+RYrAtYrMYu3sHvxSj9dmFY5e8FLFonY3E83jmj4S6na8hpGvz
11kNGsXStdT0MGQeMwl+W8RPJQUS2yI4Xkg90mJON2AYvDWsHHLbbGN6msggAwhF5+GOOcWWOtLL
w7yTc00ew0Y1NkQmELiSp2D6sW+NWGB3qx2wF5hWNS07HRCYh/iTpYZnZDeYpAGPoeUvUnqXgEGa
3hLPVzUKmtBKxJyZ2rdJv4bivac+f+c8qgR/f0Ld6buGZyVhIUbQ7jvEzgJypqC6JEHyeS3NZ4tT
1ZO9RcI/7gGq6SvorQbxcVo2aBCqigOlS+NyFQAETOapwMTMkf/VDdEMnFhGsY4i6JzzbyyPN0iO
xbnRCa1chuZdJOcXdopJdWaMFVHgTXdRd01+pOgY173di8r0rXCMp5N7vGWcRj4xy3Tf4ECQxOWS
eOcc32nsFge5/+QEqQFv43giawMcEx26zF4EsI1Tloi9U1cILPhyN5mKh+l2k3ddEiH3KUAoUR6V
Clm8v+cVQzUo28iVtDr7IRZoWO8KSjAy746SZZfedzCsUl83o5G8/SWNENKI2QNdIlNtCjTiMJh0
3XWd50FlEjd/54TPQQW7qu2x7jD8UB5kK90pux5MlWs8Ox1uNKsV675DWi0nGrr4w4G0s/siVmd0
tZK8AVZBtxrCKZlutqIi7KYrrikZZ2pVwnzOPcbBv5anjDTuNr7ulYGBoo9LjFhezOszAPg44lAE
cN2Zm0UvERir0PCi2Y9NxLPlUlYYvzEtZc3BHTIib5wnCPwAZs0PGqEJCTO3JTk1+SRdMCUSUZiM
PisqjPuLbP/kgb+PKJ+9HePFQc48wD0qQPwqn5TljUOarHjTvkuoHSThex6I3mijeqCRac7Fq8DA
Xbb27Yo27/8Fc5CNN5BUPr5yKIq8IV+uDEfd4DEC23xNQvH2hucmYO0W88Gmyp3O/lULGGdi0UuI
2uv9m8K6B4nYaA9fLPxjKvEXk0DGeHKF8Epgw0xF7Lny6pW8TTZvJ2dcgZDIR6r90L88v1Mwu9NM
0oJmAfCOsT3LHoOdf0hnvg5I00PYoup5TIOk5Yo/SkpSSI/XnC+Jm/uemV+j3xdQ4vbYQq5f09bc
U+FLkdXu3E2sUssG0RReCaLEiEx0OxjQr5AxeabtQ0qYhyBeJcLd/3sgARUtXeacpGXcAoSCsC4P
yFHMTEXPjNAQOv74H1f3F770y1lPWolZd52IhRTUU60MhFL2zcJMrq57GwJMOPWjIiwBsyxI1Wwt
g+0aeHdC+9DqVyorvlCqW3Nx63HGdPfKwqbSWFmORupO6FAnPKNJLESTYZ1UBP8AECXgkzA3GkPa
K3k2xc031vpUX5UYe8gXxSDd/HJwPv40ZuYPzxCh0ejRk9XXA7hZXmTCni5HacIS7JC3W3dBdZsJ
xa6fevmv72hESxiQmF3GbyjMJUbrE7N9kyFg8cihqTRmIVcsCjX2tDgETMZSqk4LEBodqWdyoyqV
BexFcFmV/SRjnmHAcAekwTHGWqFEKVMa0YZlQuLk6rqCAomfyIX5j++GCN92OEUyAoov9Bq1X7yT
x6KqRoTE+fVoZnrwbEv2indnkqFABm/CPYVUlbs7XjssvTqLzndfyWej+d0dEwdk+J7sEDO4zsjg
BqhGqBSbm+IWP2J/c1Bs2kyxGhZ74E3TXWnILwFpCreceXcOxX3I9vwru9s68QDFGpMofql77rn2
zmogB+ZGEoMRgTNzsy/35OjUlAAnYebOHrkCeULJDBihpYnC6LZDc5wnHeprDPaxS3QRRiLVwcLs
Ipp8T7sSM7brVtCBtswNq/4k8KV1lSccMmpqmufeUrr/foVPJXbXGnZ+U1n+zI5jcaAGtpJ7u55y
gJVptM01tJ5xt7VCsnlM2xpa54ptCuL0/yFGSLE+B8GGdUBdH/tEzsaV1Jcc85lNg7DJ0396XLcZ
dYv0e/s7i0YN2Bu31DOZGALZiz0bcovr0hA7kVv+SQgr0osPFtIiiJTXnRk9LeXhZpXfmnL5emIF
K5qo1JVf9kPfVYIF5WQIXCT5i+sJZ876vm7e7olqip1SR54T1wPvnUEUOtFDmqiyF9rV8vVPzBtU
aqn9a3h+AnySzKxBpfYUpV3ux9M1vP+ehS6uzb9lwlHQkwbqY+ASNw+eggJhiWsuyBZT0iDHwXUB
YibhEp4YlZVTg2JGuOzA9bMXPqKy2iegmxNzx9YZqxexEFmdhKyLJmbg0dEpxi3GkQfqqAe1Sv1R
31jFPVWiFVEjLvh2YNnZYC5IIZDuHzaD+/rm2jU+zDf4nxDAYty0tm0UE1kz67ziTAKKDORs2Tre
bndkm2ast+6/mrJwFr/SOFkuqYymbWVfp/BMnlzsTfceMtIanZ0CSQO9+n1AivxejxAozaoG2+N3
buPrZNc1V0XkMgoI122oLxxCR7jdPiGQ5eQQKGIOc1Avn8QSMY+iBWW5s9/eicaS4b6H+RDUybDf
u2X0x5zoU8XsV+DKL9Ur1aMHTqpHgLn0+EvQuc7DEn0olxDgxyImoFBu7edZhUh2yNjBcPwq6s+N
Cq5+4oL5kMIo1/r4ZXsntoT0wTd6Ybnjy9oCmHqnAEHwZFPDKPSR1xop2Svc3Mm0tGq/1xM9TYz3
rtsGdSHysQqvYQ2AxuOFvq2p8E4ZQANc+jGuxH6qt86/P0WmHEdZWf44+ByxL1mQO1r9XLF8YGBD
+qtJ7Z8iKb4XdFo1BsNXekki01oAWxZ14mYGGVnUdyp9suT+j8ViPLvumiMTyLpxBtH8x7gd+5HM
V9/dR6JaIGeRIniC/G83w6UiCLsUUWgeeChcLz5B4EdJMajMHAqAIlL+wosr3wP7OfHcYst0/Uie
X+TN1TjN0onQL672ji4sewee1x3lNaWF5MeVxsXjfR0Vdc2Xr2BhcItMwUYCKRg6AI3D4AYPngmz
fiNbgHsNoLVYIjqV9zHlVg3i9xzY/dtwGMzIvgUpQhWL/0eRyASPXLQAt+WijyXpUhHlu71V1jHE
2kFBtkJqwowzxUKzzhVxDdxzuVyixFinoArKxxanknjljhv/9/ooZfnkKSPV0LB46eDTLV40nNUS
duprtFH24AWm/IPH7QI3vcybwf06frJs8BsQUnqQYM9GTxPtoMTZ2EGOOLWo+zcsqEGgYG4N0ycm
ZeO2IM1y+/B+fXd6V7zC71XltmpUoq3vxEcIXlcrZ+WoEIFUUzic3d9BzFeEpYuu+X9pPKrOKiTh
1pbGlGwAFFIVWvj03wDSVMf1+CIgwiYzPuC/JMWX3RvEBDP2/FpL06bIEZPaTSMAXz/jc8o/ClfT
JPmBQQdKqm/DI9ANB4wVYYoGstQeUyY3rjLiYnb/v+QEyKS3/hn1/Pj1T8DN8fLcz+wdta9JJs7Y
3YJPAvhQ1OxSRxQKp2EVaMogq2PyDjADg9knXtuQ0PMEvC5ViS8AYa+EmlNz9QBF/L7t/pFwVzMG
G6AUlFqArglol6q6b+BrkJU5miHRErRpWRgWM8jmeH9CeA+wTl93O28pfn90bE0Jsw52AZC8Nfna
x7nDnb8DHZ/qy9od/iV3wE3wFJO3lOmuyNDCPaPAbGnU6/EHXVXUbNFkdhCHQf+pl4ZRyQP+QF3+
b55vVTEJbOtFzjg8S86qgERdvLJQRvloQGouN1SRwU4Rc38K9/o+dCI/1iXMA1/XqmGgDhgTSD5p
fJVwN1yG0GvEbyQhrdyMrxZ6lj2SKMDCttVWVpzxyG0HvTyEM/FKEYgiz4PLa/I8w5A03TNhp1EU
PEJxq7QI0J/RmgpuA/1u6+uOob9qw3ns2Aqhm0L+D8OgwxfjT24uZQgQ9kL2+t5WeJCGBYGP3S3M
CCQsaQJgqEqz5ZOGXcJsmjswE9yOt6ziUQFy+/hurN5vNkXcZs8FFaTqw9JjvoDMQqJsFCL7LLqC
yUkGL8ACxAbh8D3WPnfc5DLBnEZHuNaro1sc8wYK+yNutruNRI7uYxDxB5wKzfW9MxtozDJsPQNA
t7G/aXnkeSEf2jPacYfZ8i/F8p+Yri3DMO7y2GgOm6tDVT3r56pJsDxb/IJNMKx3HuFKo2xk/e+u
sFfl8zypD2/OHmzW4TOi3qDIijb6NtDNtNWldxR7jeHgH1CIgphx+YMYXZkZJa/bhNbnaloQxtVu
a4+6g4nvihLYeI/iqaKs7XHGcUzzxty0tuiDvV/QhSL0Witq+w2+nNZMdRho5H18163yor1J8V+G
SBVD99XBG02S4sP9Lp4aznjRMRYVi7lyGrPeCMlHYH6eMKBim4EzkgVvG1hYlk90G0VfW6UK3O+z
c/jMSEX3yfs2S6nn84t3r6gm3ibJ9g7gH6UroVVUAeCzKVjs1oF7lWv1FStUUwnVbnlDCM2/J+iB
i8bfq+cH/s6qrtV31yX9HXidYShyOW1Mi8Uu597P9iZBTJeVQ6LND2htM/nxqkCLCgiCb8BXRE/W
XNKeNEmjCTZC6D22tny/zwRkg1g9oTxxHUMxR7B6ZY347G3+ojxzCVkJ8m9rkq3LjLSuGEwA/LK9
gQUBCosP5N7FGvDqKtc5wBXyrksNK3hfAIXm2PSX3JFq7cXEYjCrGpHNPPE5utAkjNCYMywFdQao
Z4qZp3KwEaHoQ+CUiJQLSTPiuQC9PHRyHzNHcORUiaeIoqSK1HXNE3fEpyNnxbfO8jpz6zPmlHch
INYkHF1Y1D/QqbPH0ysJgYYLfyBE3MkeD3p3VCa2MvFqNswqUIiZUiScoFbSxyIHoDagUffCFYOy
SPEl7cx28YZZlleFmJdyPKDXNvl9z9U6tbxLFloOOwKkh2h1KzWW/x2xRDKy8VDfGp3pXjcIQd3T
gS0OtMjy4XK3qPrFK4pnF2Wh/DuDXRsXpL+lUuu89DDrHNbr1djbYgLW1PUMtuvQon3bDkC9/XFX
IOb/aMUCzssTb0PgxcyZnV1sBxYhj3bcoE02uziyhsgCvfCbqpxs+JZir0yI824uoYpvCeExNQgt
C9sDUjAJ7tw7KHqXUlzE8/bIT7y14pUY2o9j9dNg+bASqhkWGabZ6pATHkHciBDbucmPsDo+w9Yc
sRT8cFUqMG+M9k/Qv8uXxV55ouigz3zGyg/fE2qHn5fRiJmFjl5o2fKsB/k5k0gosi/cUMtiSl2b
SnjdPyT2vA3cICWKNtpdOcfE6sXlreZfdA4Hl4p6WwVZXCyZiG7QMlEteis0Uk7T4fNT85gj++Im
RAuJktGnQORcFfp2wrc+Y1n1uLgYhsOXke4mQmjgL76QJ6eO/9XcZnqN3Y2SZMRIrCpNPGyyQasb
9Jw3H+6ljY04J0hWjp6Ti28hYeYesEXFOR4vgllcpuwITogFrTDcLPAjZYfivLk+SrTrFgI6eLEO
yK8GS379L6PcpDxtDg9eQ7NbHXMM/nkIpFQFs5qfGeQe/VVwT1xj6TYMWl0iK2I2RSD8YRDEJ59Q
ztUKoLuBBYwRFO6pjSvsdyUBn37IyPOAn+kAbv/3TJYDAPOd0X0YY6d/BDe1/GnM1BN24YXC7XyU
oFlbwMKzhFsyyxAQwQm0e41i6/tgP1rif9BgT2UVJHr0ZsPkF1Ni4in6dSg9nOWmV52L1bQkzEdp
YcbqHWmcqYySr94zSQSfUEwb+/hBnyohYYXE1Rws8Y4mdDmsJiAwFUJJo4zyOgbdDomXNXAuXgfw
U9mI6ZQMFhEg7Qcj2uUtkI/Jdvfv0TMq4CGsaFxSMDxOxBsZXJKbnJIyFH8hICFKVmo1sWNtwygz
ovRiBXx7l0iimO25l2xvQX3ZyiQxB5NiHIIApioVT3RkoSODXKgORqRuNWncdrUFm5zsHqWp9L9v
fIkG3ScwwU2Z4oWgGJQ1uZF9/RYK1Se/MP+8B5u5mb8bI6FUZnQ0596MN0dzHbr3zdgdYFT9LVRx
Smglp8DxJW03sErNnPea7wtCAyGbSnw9eMAo1kg6ynIrzELz5CZ4u8v/b5ajf0o3nQCFWgQVF+Fp
j5H15mWxin0om3R45eA26iMEYoMJ5xW9E+z5B1300hnx9TdJJ6OaXXrvR0ZymnI3nH6y6GTrM+CV
eD3ocRj+wx+gbmMk+xcRCFQmNUEMu2zlApCq+TTWzGQgPtyc26gd/WpVFl1GP5ehAhMUl6rcPOON
ZR+t5gzBOQ5BBJnjRqe6syjehTHqPI+MipwImCEBLRJ//AtlyxdS2W7FH6tTOoVJdMkZYq7uSXuk
wzKaoMwwSaJuZxvNBi23kMIWEwdcQu+72sq5PSd5t/yRr8goQZKRebgYkdweZFpJoUuVWrKYQCjx
1PBeeunp1EzFAIrA8qK2Kp/S7qQ+vjftbQaduZi/LBmWibO4VQb3J7zt5y6iDDiBccXHZDFiEx/V
+f0wl3oJFl2HIhPCbDeBlhu8F9udTmrgpL2jq15i98KDf9oL5UeDFJSrZ5H0j4HWk4n1NEKo1ZDn
Pvwz6WUsNJRCBxvkSGgNzq6PKSZCwqe13Lki8a0vLZic1LHx6m3ufu04y789Eb24QD+b+E6tya1w
U443R30ZOlcF8M7z2ibg7qVxTZB8M7r7FBLR/TedOzE9EmsjhOrFEFVspX6lcDMZmBpdW3/BYu+d
EVQB98BfK4cb2cV/oST0jNEzp8Q69gwLrQRbNXRLdSAocRXj31pXDsr7HvnMLAvKQWJ3eq753TcV
meRbn3yBBsnrtqoK8AKS/xwvAl0j8Tz7Sa2F54RO27myDLi6d+Ltqihg0SCbZgy/wuiSCe4DUtKt
mhOXCrCd3/fV3/XRviSUppLKpT4hb7zODssgx/ytEQIWuSpGQMG+X6hCNY7rs1c0taHw03tMB9+o
umOOnNO2DE2SNCQFtWDvHMVWk+8mG/0Td5m0VzEFLGwKNiLgxT7V5/lSualmmgQSUTdTaSBWacTf
NqeJTRUzbQ5FdHPc7FBZXxtv+Izp2Gn6b7FBXf1ZaWgXAO+DiOGErruD0m7sMzLtqHwNgQI3dZgK
+HdyX2b4up7I2A6iOmW0GlcL8khSXm2FMipd0IyymAHLu4PJ+hNxlwymC1yHFS4UZAajFEWrFNtp
ErNJdOv9qhWqwRtCEk7q2BVMmvHvBJ6gqS8tKEOadoMbNtw6YUVqycUjj9uHkPIc8QJJspEfgz4u
Glxe6TgnFYhyWck6g0mw1bZ6jiDo9bIDhcjqi+W02C4xvvGbWkA5KOje/VcVH0tyQ6dkM2EQ6FAH
+t2NGZGj4bsmoeIgba3PvfKjnWn3Kwhoj8kG8IFOiO/yJrdnqhb9qEIWJfEefZzomXKFatAfunZu
wuObW5opibamspXDEtuLwQQmCl2fSWVvPrV3fPKfP1f7rv+TKrzAUj0bNSD1gN4akC2nLe386z5E
irMwxccIDIufiEI3xUoP4hbHxGiCbp3H2xFsXCVhAQ7D8Sht1H1NubofvRI7I6VLBS19FdNk+Qaw
7CT/IgliA7aAEgvFvT2KEfDPGF50g2kNcBAMCrG9kU8u5KKjMaCMlmMNZdEutHGdX0IWMbpuuzwV
/NlZ5Q3wGq4FLOl/MKoaEfMa0AehiAbKEwSc7qix+YrVfwRzroiQiYztDqh2e2xRiHwkbSBgJPdV
YbAEuoT3IGeeLrMcZaJnKcDPyMTmISUwemrifoGuxW7hCbSRFIsxZLM6TUgbQJ2ctNH0Fg9kmGLs
en1eXi+XcmjghACaN7v/Xs9VduxYt/6etdayBSC1Z56RfGg8l58BEidBRov4Gigf6jpBfwxSD2MK
g3kWGcrOJbU59qmyjk9sEcShdSYNjzMcRatLNV06DggwyD0jzY8DEkPjlDXeQA/nXKN6zZc3LQQo
SfYRkgsZM/whz5INDG05VKavkODFJbc3zLjtxIv8Tj9eDGPu9cDgC8W+0T0jy+TjxHgvgKpobjRK
RD/l11V9kwgr+FCN9+XkIFJTDtgXx9sbXHbVY2tSEZSpju/ANm206lx4P7xR1MMPUjAA5l/R+BEe
3OAEID9C89dgXH6m8CnukAYZ0qH9PRCnL/S9tji632nLdbJkBrJxuiAw1HJ5uuQ0T5lUfEJsAj64
HYnnyXbGsMpC0YbYyQcToacS5LupA/iARlQqZWWkz8yywaOcOcUxhbQgPlJFzpqli6odv7Oh7nGO
cQYPYc5QkEjsDOTF+iYVs4YyJVU/5l7rpF76Hi3dGpAqbtLzU5EG6JbHO9Pa/zAlU4EU7tIDMvyL
jPoVBNmxjmUrMn1PEac4y3WEhIQWvcz5aYFeWtrvV5QdTamThk2Or1BD5vC7jOvc5Z1vrbPzFNaj
HRjbYjz/qt8Myz2VlRQYPXMZXZyJLP5dZ7M8fbj6tPYjWA/Uqrf8pH6UB9nbTsOhiBD9IPnq/xux
jMHbr5rF3GwP/Lsc9GeYOmzOJHZ6MDDKhjoA51HGjGUoHCcfU7HqupOytyFA/olI/BeZJpKFLp4b
dC4FePXlhffdXUGcVTDI54slvfuTUIF6bpilfz9666w9SV2tjQXx5kfIZneNT2Vz3jW7TvSpUAAX
ssH8sMXH+ZYB0pvQc2inPALju7w9o32dqAo7F/pU0z6PbxVFW5bj2s+9SjrHaEtG5OuFHd1fow3a
Kkr85H8OHHK5eKpvTPQWoQb1v8apT5kd2ZIFUrqC9FAbVzh/ZUZT1cpopF+Fq+9+4XQL2uIz4pAf
KYuJ4skeceIwyiDONrPsd3O9A65g2xcCcWiZR2GTm9NvvQ0VhMNqX8M1YyyGrREOBvBiM+OYJqBY
rwIvJ8O/2+rFTCHba+gGWkjcivoU0+aXcuJJdzp1AcOu5xQMi6ir8NRjKXEWHK/ADDYd2gYpUHYP
I25Z0n9hwpHvXMP2u5zzMLpKprq4SoNwRCdiTLM1DKI8AX5PdqpxRXx3FF+yvCtHhn6Ut8w1WXsB
cQuDbcMhNJGRmDyXmBBTGtVNXJ1wM7HHWvkp+3q7K7VC8s9Jd3/PnCjt6EEvhEaijFliTIDKgFq1
Z1XgrDlPVWzo97aR36TsEtl/zDvUwqZmbOZyox00a4uEYKlQPmKaI/3UvJxSGc1pjTLn/rYaEdsm
YYGuUqN970IkGGdsA4q5T2wq2fTukVGlJUk0WmIDUDD+7ogJmPY70cs8HofOqP4Y81RX/c3fzPXB
MhO+nPnHZBT8FP1tFFXYgFvIvOzJVRvjuLjB0q20ftVr/qaOOjlPclhFTcvPpj6NR9TvQ1/7IOG9
ZvM1SMmfgPQaYPpkEe2Us+VI8bn+df6ulvEnJheQFUDGWXuNQUY2FiNbF9JZ0kPl9i7Ef2YzCFQo
Uo5hlmMfVsqFNiXZtwXKys6+nItALZ7sXds681FlTeIOPzqQX2nSA/zTOKKKdYrW+147l2NnTDi9
/vyKCORmGBRoND5J0vRQSodo4U9HovMPUMFrrrkeMvLOl0HubnruvVoR6xEBjTjgWOB55/vryepV
V2eTYw+Btv/k3VFhtlqzMYQ63zsTEmI17HPRbV7sH8TVydEytgs6n7uoOZuTP144s5CJwmp1LVOM
Vg4f+Pt4CYVx5zCgZkXJK5+8EnIxySLKJYrdnxbEPLu73SFQrvy0oZzR0nWh2sT7gCsxqO0LEr9n
rjBSbYKVcQhnIB8ZOAtfqUx8a0o/H7YxIdX4T44jxyYZZ1OPLOemhxWZHLKJtLabIyjnwfZpnZ6S
aKAj7zuoAmQCK4r4eJY39FeYGaSDMm9tB4c+zogwhuXxBL8d/S60vkqr6YABUESHBqW+W7v2s2AY
sbY+BLxcY9KXYiIvT5/4aIagDQXEEmQ0RzzXPka/JOyv5PpzgkNTVjR76pDpDPR6OJzER5zkblK8
rk5Lir1VXCAr2PFNM1YrJpUl7YiqS9J7sTyfH0vjbD2hZRDKeyLkzGA7OCEc6uyjhSW4mxQOSyS9
LQunKT6QRzA8PUKbDQWbR8KX8GrzrEkheBvjRg9Yohc5q6LEle7QeadUUE1PzAoZbjNXZtJ3C7Cq
viXbOfmcC6i18guiOSJEht2S2VpUFe3pXzAaohPDA8jdJcqmQlx+d5zM3a11iytEihsA+dquqych
GkwU6NN9M7DZ3scKcwhtqwsYLNQGmMkynw4owbNe2hYYZBHc6FzrHUHx4anV3Bmefb15coxsgUuC
1pHXrQfrY3CncS+bzxeZ3pTQMSgoPTeiJhDMJxniGf3IVy8nCwIfWjRrekE315Vld/TfEtENuFe6
CXVHB94HtbczC4ITWWclEanIzHeJ8cH0NChhi43xgZzqXaYP7ZSbulIF/I1+1d85Sjjn4josBSZb
B+AlWluZx6AK9G8QfeV60IkPmt5Ymrrrr3e48YHY6AVK1OlOtrMjPRGkDd3LQePWGrQGfBjjibxh
1iw3Dk3onaSjIAVFy+jvo8h5gcHW3WxOfWvM1T3NPDHnyZxY/KbrZNEHEWfAouiWcNVvBJsL2ZE4
/aNjP5f3uSKA1CzspAOZ6WoC8oclegib/kX3tEK65rOurgI1BWxGUomCFW/xTiaQFchHvgRWpVLk
CzMiME+nE/EAzfF98JOU62nXDkUPrt4bBhG/uC8rv3FPnkU5XaclMHF/fTQYbNU9diYho02hOKSv
slTskhIk9haa8Te+klTbcTnf4KhX1ggEDAxRakOXpC8nYfeUz5amauW+lLqqNfuuZW3ihuyzK84H
+Em+QHqrHFOGOsd9fHybt+f/JMCpq5LoeS8rPgyJH7oUsznwCnxKgTvNHFJMttmPfVHf+8DQXaLC
yUSgeuxDi/bZ9+O/Pztb6gJyI5c4nORKFjcQnT1ZBI9X4pVXVeFIfA/j6LSwZW5SJlv49BI3s5Rn
xGkLUCC7aEWRCO77HhKXRxa/DZ5ihlfhZk4yRAddJTLbYSqcd04Yvq8+LxA8iIprBHt5EFiqh1kU
5yNApPdUF55qgSTFOM2RMkLWikpkRke5+U7/EM+Y4eMLRCN+VAgu31omCJH2SpPUsrTwSpwqoreV
NEWp1zEvasc6EQEkjeD5SZ4qULhBSb7n2DjJ5fAGzyIZh9NQ035mfpQFm8KT3g3/OWJmuLWeJWbq
rwaS57YnbhuthwpUGaj3QCUtcDiybzdWSFucy3TBKHGwMAyaiLPr340WbfSRW1ke8auz1MhyfODY
5Vlhix8FN0fdzUF01OF3/YIocf5gKDAOo93TPn3vbdmkSkXdyUf5y5zz/3EXfv9fxSmrnxkvyCnM
jZUieZZXA2uJ7AmxH7MpEqZ7GjuHzNouGrCwp0aAqG+F0FxvMkM/Tbwe1a35QqXtnnfczVghg26o
Wo7L6Od3f24OfsFOFTW5Id+bbhqzSMxa0+DA+zyeGjLWk3Ht6HxuFTuXDdvo3VZlCiyiPlQ4GG6w
USik7bHYKAKhmhZG1nr+V0UangGVtfSim0SfvTuh7ain+7CygNGjgMZ+yBVF+baeTsAVls5c25x+
rOQX+sbZGupo8pY6rvpFotiHfLsEkmJUKoK5UaMfQQW+7Z8LydEXt9jfRp69k/BdZLy+3qVGbapv
GUOY4G5QweKRCpJjFwaEENhODtiG5djEPkDJ/vEQDio0hpwMPkSkGoiROX/qGsYRxC+mXBlcq72D
x8hJySdxsK7P02RSNuXupJQlx7le3JQIAGxv9tUdB5UbnqF1KXVaJn87xd8hXU7Ig89q6pACzkjX
BQUq/eENF+Q8VI2sVLgVQLK6HNsxey1VoCa05q3tWp7ftpg+9FcXhli3t4s6DmQpix8i76l/ch7K
rJVW10aEVW7cwjUpixRKi0vXaqq9/Wy0A3Cujfh6saoiaj6ZYUphC3pGwKCYuBkE47Vc9LoJfd6N
DjnskBShoTKxdVq03XyxqBJcyhuTBGBQjOiOgnJ+umNCtJBRYkUj8tO/n3hZmaJO13l19+xH0G8Q
Gox46bQfdabLZpbgQgRm1a/AarCC9Xs+Hp4SYKrvSbprhq18xQnd03deQhVdTKwBUV6bqMSKbqTQ
cV9lrVjKzy1iQPbm4hRJOjBSroW8aereCrcgnhiS2IynJ8AP+pGxQ6Ke3059T3GtWE3dvwp0hFTg
gni9mvLPtYAZZxQe9Zte70D6ZqyBVunMnplsh81EnMorJKqDT1zhxTSV2IEEvcz6ejWdFnJsEtLx
31qm/1RhdsgTzIzf/A5rraBbzr6BC8vVsV6/oHD0ys99tPBN9mj2B7GU9/1QqJiFKDcqLJpKv5z6
R0jGM2/qBtfp2Ky99ivG+c66ojzPYthn9xJDrqSimuanYnqEgBchag9TKhRJEZwq+4uKvEdyEEPh
xzDt6w7CS8EurPG7DvZrtr8rMXecDYIJFbQStZuKrbsJ4MMjNHIImMxWrTihO9NhFhSalMK+yNfv
qEKRzVQiS5g5KOavtIIPXIb5lxyao08E4hwJl6ZeMSQQbPz4BYOGqX3T/u9Hd10R9cy10+zadZvv
xxGnPhcu0Ok7lH8zYsiY4RlVSMvYejj+BC2PTlyofBS3T6Na5XT03JzYIwmTcxAOXXdGld7Hf55I
gqy69PpnBdkctnhxTppruj6HEcryr/0gpoLTgPxET6RJXU2ekq5u2JYv+mny0H9bYtyqdC8zKSTU
sLVXe9UdPmiMaPTHOZDqPTcw6T3ntp0IT6mzIY3HHNLY0Av/Ya3/pWYgwVsKi6tHuDo3UkVBFahp
RlE55ibNFlOtVB5vYzXktBasFhz7G3Qea7qV5N8khIF9QAES4tTdRJ8OlQvYuEipEQQtdN1v+iOt
3eFg+YfGwUqsjHkvuS+6HHAqIjPUE4rv4LagC2KZOqqP37nlGBLFBTHs5ALQnPv0AQF1bIZInXS5
BROteC3FByAVLomk50zm9bQm2PefTmc4eQ45Zni84SojRcEsczCBvUsCstWMl+a9aED6r8LLJjD0
HUJVERE5Hkzavz43REBqmu7bgGsAhgY/nzL2qb59MKgNC2Hfcmo1Wg421tqkhYsXIKb4XAcVyaCh
euTzh4hQ3AQ3F8w8E3k5nWYUPiekTw2j5+6RuLQMLtcV9o+HYvyF1y/FL5PXPo2mPfwyXzmCb8nu
wu+QGOQWOCKQqf0t0Qn2MolYwrVPlceeSI19HAVm3OhisYairCJV7yCDXr21e1pabZLM5jFIVi0z
lMbqSy4xdwTA5+KmPhQzO1YtKKz4BhNS8VZqFhn5U4BsFT20kWrkVjfrbDXaIFNfcIiEBxNV4wue
aoWSuOBKNLiUB+bnEDWEUyvAPLyMbRP0/s3Uchypf1HXON4fRvNYEtTiamHbj3F+xWxqKziRzj52
IwNjLQWgs5GzFdxbaWNYQTLdv4gap80W1YYC3hTQlWDgBoy3ayHykmdj5BUKzlU/klH27TjcG4HF
ZJqBTxDPHF/qJ0tDACSEhln+BHOwncZpweVR+NL5THUjWkGdyfwEyn/Nlu04+iQ47Vu2vqjTQM5l
ad7Bj8DfKj/SHlnwpFpR7wdMzP5nm+qyEDzvDG6JT5pEcaGdLdmP7tTfOBz5EFrv8yCQTf3LdMtD
TxkZeYd3qc8csFd+ymRK4vExEbnuCwG85p9pi+P8Wx+sUabGTBWxELyQglV7qwTs5oFIkliH8uto
GYETtU7Wq6Rf6HLAzboTZm0z40T50vrFngQFCIyrhOGHSeE3DK8Mj8qeYXG+q7G4XWX84D73O1th
Jvxxs9lMDyihHLreqbZiZOtQHwiuVdPf1EE8005pG7ByLRqOcen9/fIzvGBR2q59Rxu5KicDiKZ5
YroszBdqfcuPf0W3DCFc4dvA+2b8z1jYTMHrD+dcLDLkat5jbia6JBkSMK97bS+KsYugzkcs5b4p
gIwJ4OAd6JiIODfXUiNAfjX0vNcVI9ILbGxl8NmvawPWU00+t9yHrRfvqf7zWOCJ+41FkEOJ2ITR
HxlfWf4kC5o4VdOavKWbX0g/pA1qBSdpo51C68+pNGef9TlbW2LqPv0p1tTZLyKC36bdRmN7lXNL
HOYhL+HnWh2AIGg/HsQNayAVachDNDZHTkv+AcgnIAn6UnruqMtcbouabshioQGDUsq5hR9YVXST
ht4DZriEInYfoOTs6W4bF0FM05N3b5l1VSUa3QEmSIgfUO81CJU1s+M76YTWhR5q4Zf/LLBDp0qF
IH22qh13cDYksxSGR5QgcLrGi1AgE882REIowakyafsD2AyFAZUIKxNyFuavkQJdu/B67iW6uSJH
O8nmvBKPK5v9FRifydw5B0F4RosuCrzqBdgIIMuQ0hSbCs+MyxPpGZIgNILqENqOsoPvUKGmYTlF
HXZnEbRHBX8A762Ngf2UOzMYocaaI4nl2UyBYVlCWVA6/ag077jBG3EG+dr3jjzYPu0wdUoYKMZs
CzEKKnT9/kCmetUyGyuRMq9fCrrX+BsM/JqdTqSjuB+nKgsCRcC3bckFNtIfO9awG9XqGyPvqisG
o5SID7qP3AfC8bkt8feJKR08bVXFwpMJa6keZd5oMCbH6ZfvOmSYUbRxcNNKelEkv8LSwa2QYXZp
eaooKfNBXo+aCSUjlNHgqD57ej3kphzVy1LQUHHkrGzW9gjgVC01D7hMyul5TF5Y5YsjNt/o7NKx
7Od9q0Z2bkPiWFBnA1X5YUiMYmsWCRN7RX//jk6fhOFFH07nG2ca9VRUmCRly12sUrx5DJtLoQnt
Ag3345ssKw7X7n2O6XFwBDrVcEuf2ObY+z+mZoaGIyX2xhGKrkUqPM1dDsnt/MbjoG3a4IKqXW5/
+2o3zhfnUO9wFKV51w/9B0C644BrlnjByDFPq7k/wEwhAfs+l3Y22UFB9AVGZlboIpjhRTrsnGij
oFWQh4EFFXWxWjvLpm64Q2t/FtCaYQKAIlg/tP6cYZAwTTB/7NtIHEYZ3tNsuWjcmTKmnkLnqX/K
cYdM09s70zQuNEQwG3Zw8PUXAjCjVwuZBOoQNAFYzGdAv/+lRGw5HyBApIFLVPXSjNS+svaWyTAW
GDQKJGagKxjYl3tXyi5seXFhLWoAeW99fRMxmHrfWjzC+8z8cBy78RUnTj3NI5ZjObf1StRHrIlG
BYNe2mZG4pd/68lojendguUZs9HyY+liQZUG7KOY52co2vJv0aJYMdicAIA+AWTzbiKtWlZ5wkHe
2xxnQMBRqYW4VvMhoZQic6lKkPozjCSuSyucXmU+LFwi/TwJ0dIfGW/XxKuXjMPggK+b613pCfCB
IhpeLnIToalQcFKVWmKZpsifOOjpdA1TEsISEUqKco9NVxTBYY149Bo7KaBicW/PYyQVHaOFDsaw
KrBGnYwHAupxY/OJphzv4RXIeZDW/ly4oOKkaScUsJ9V1QDzG4QWI1CXJe7V9sgzcKc45mYhVXuZ
sxfJycdX9a2tpJ9C7b88MQq+WsdtZOFT9VjqP7GudqE4agiiF0cqpMHfbTBoQLCN3sv18ISLbzsC
B0zISBiZzYPYin8wnjuGPrxafdyM7g76v7XiH0y9MQh9GWmG4xJoUwS5Fk3oG2J8ohM080hjC+q3
lPOvCOWvbxXxs15CgkUdcwq0oDHfTguzO3a+8xkDb2AvW/V9RS1+heo/OlUvTseI1MKICOKm3Y/8
mziSk2dhKls5nTtoWSlHswvgTk3gwrD0HZ5UHH3d8rZMLvg67KC49RGYspi3MzIG94CC3QqAwqyQ
NFG4o6NFNhJDkXxmyj+ssS31BxJi9g4zngOF1IqWbflvigFiJbAkjszCFCdrljm3a9LKGMuhW8jX
P+BmIbuzEmHUjpvv72zIYtKnPBgpTS/qpLljfQQLoHml4FvtcqvDdSA+IQ3mIw/thUzwDSC4CmuR
ZLI0NdHGVtbjDpQSac4ZkUsiB7J1YPFk1UjlROmjbJQSBBdpb66cnISxtOP1bkKP4uObGIsF8e7H
h3Qt+YLq3N5lQcke5ppSOGvTIAbEVv0oT1nc6ojsvWAnLwpnlHXZZXPRpmKPwqhSq3G7hphtmDMG
mVKPiAVgDvLRjv/pNZ16Q9klkClb2buuQgIsQC12GSn/hyTQdkIPUbchPwWOQheL7xSiiBsAQXyN
wODsrJny9HY+29HeW6sEuiwjmG/FqR5HT9ox3kmcfMl5CPpZ5JSmk3sqr3FO/yHsvabinMzQO+/h
sDd2LQpM2y4N8UpRd6Twx8NV3EM/Kv6Ca7J+cv7QkxxumUKKCeuNC5GP/qESKEJfrPClcPTV7ZX0
RS2tdKuYFA1Y/YQE9usn8IXFkoSzMagWtmlH3PFPpo2sWHb6yle8fz1cEW4bDjUJwrMsTTyl4by3
t0Z6ouxkMm898j1Keg4pxIIk9GoVd5bpaa8YhYSjQPAoo7OlwbvP1bp5wFmzq7qUF/fJMANPindm
37AUjKP45VTZrzuJVW8AKNPABbl3ZCTwvIUd6yLhGGNn1sak4a3xvC2uo459iQPALnmXjcdGRqXJ
AqSx0jFtTv54WMxXQfKsBb2+PkKwG96Di3CONIz29i8Hnp/UE7m0JK0Y2fQvJKHd/PnVmryeuSZB
x1r6BK24epfToSTuTaEweLY+omeMFwGatyCeeuVoBDNskQ+6CFiBoHI1NTsQkoxwdMO6CrgzAQw1
AXW1L9v9AUF39cBxuQnP9rK5GGqJaJn+38Zd/vJ2+PvEaAK5qxeMkh9L8l06xxGwCmQgkWE8eOm8
eCeXw3kjcni9ztLMfDh8thN6ui8df/kw+h7gkk7Ge2i2fKIg/nG60yFzx1REF7cUDvQPPDQFPNxb
aOl3POehBIAbqSdUPdsvG8BZEDkilqRohFZoEXGCma+xk71kS/Bjpr+1hvGPFDyMrxuk6dZdjxw3
VJLkXNbRTZvi2DGRtk/1tJtJIaJR5140JQ+xUhbD6a8l/cttyMBRQAiNBEpTkawIcid1y32e30tz
AkGbyJm45AhZpQznMmquuXkgjTpNSsrqxDC3SkYWmnlZx8YpCqjWO5ExV+H7h357q66wsDXoa6W1
d0GLTciyTmffvkaRSFgE0gRHiXtFjajrhAyo/o/bpCMd/o97ynUN7tpL4i4NDYtvVWjR2Cqi/Sww
ddmc6H4egkv8Rppz/ARgzl1gcRhlBLoVQ2TI0ebvhs5A8JZJ1u7esShNu/tn4UrKAsPbYIoMtuCb
4y5wDq0kY4qmmXtDu5AL5SlUXwiVG6ohSPiCLDkRh4CZpBQ7twnaLB6bhY+UPA9FDuhPey868Ryr
exKs8cKsDEsfNVkaQbIF8a1Ca5zXT5KslFoUM/PRbIuPvT9qtaF/qeqaVeBaO8U0wj602ngRni4m
rq6Sk3S2pWo3We00DdCY5e7qF4GZbPXLz1e1nTPKhgV8+B4Ve2sanijO362s3pnGRbMkyG+NpZqG
yJKMQ7Xtf0w5EK2Kk0GZKdqOkPlI/FaWZnXz3IQJSrmUH0Qm04Zr3XOe7SxsNcfpFjSEP3nmn3T/
4Y5krbFTFeWiL9EXdlCAQGwahdW+BtdLsE7BlRvpncSMS+r+IXHOmAJqhermk1lXbZgisAinqJ+1
gb1mdTD0XIXFKOdzBwn7XCEW6eh0qmdQL2W5pwQYpPo/FxImsRBWsrW2hBDHbXl6bRJUjyEdLqPz
pP8KfklRxlYM6/SJSdHq71TM3uEgvFGd13VBAG9kCzfqlM4mnlnL5wg5c8nbI8O2jx7/ez7kuaYO
dAQSfwzM993l9wV1tt8cuobQczWwiXfUrhrr79s5pRcSXFhBM2DRlXzK/vbSH09xHL+MjIKKriat
m5J6I6a5pBF4zAUXMy/2cvWxxc6fjnCAnCu2awZJs9afbfGSq5NtqJZpES4hQrYZDFqxvDDx8bHa
otVyv52W+V86+BYqKrkpg8hcgjeb4U3XgVkz7u83uJTMM6+O2NA/XwvNRqfGGdItdMLloBVLvl+x
tYW+zgCDslDIgbxfZbpVXY+n+RPoy4qS5n5HtzbydqIGVFwVkNNvLmIaXVmZ18kQRAPlTJkcSax9
5oPmnAZ+tfxgfspKzXCFsX2tz6W+DH71yoqLjR7sb83ELAa2yawHF6brsFDJDonAesiuIPfbZYBF
FpjyjUp6t47nWPUHa0pxkNvGppYasUdIXhI6v+Vfp8/m8Jfw14lA6nsbUm65yBb5s4i9AsmGFQEv
vhA9ffLWlPd88MRBOhS5jgU845zMNEH4d71J+fytc36ja5cNJYnNl7+cjW/lvtAy+edrLBOZluLQ
cXkEMaynLwZeTCMH75lCNyal7O7N/MCpvhz/EaYi+PUB+0NXevXyJF/n44RwZLHUy63Vq5uvLBw8
qAA5PXA0Sx8R2Z/laBPEhpuvb1FDbDqRnyDKj0he2ZmCenCI9TzjYyqVL6N/9ZOgM5c0P3ajjzRV
dXDcgJcAaScWflYYVFscmhIQYzYYjgo8bgBv08oXtmRSvG7ozWVQqbzETymc/ihnwwvQ8DWktx+e
nHK8yO/POJRURTOblklI8ldHrs8pp9T3wooFR1LWRWe5KxEx77cumU15dudQgJpTJxuVJ9adoc3l
tn+ANDiiihZuf3M8NGItoY4Mx38kn3Y1Rskv/XLaOYiyVidnXa7fSxrOAE4iyeCTay4F3xOosku3
fxN4kTF+c0j4eotOpHUjwL+L7c4LbvEf90qjj39/cTummIevVUA3Su4FpP+l4blDCi+uQ96Q533S
4hb7v3h2nmg/ecvbYy6TreJM6iavuWseC2HfnXKkrhxvRv9KZlUMKRhlHPB2Tcy6s1lN4oCR5qK+
GnXbIhaxx4e4MQzGFfVpF74VS04nGQjVNhutg+29pBwA4318LPG8VZrRQ8jECFCgLUhc5azPvlV6
Du8ExGaDDUaqXtIWItzEqv9k+P2zt63daQ9Sn4zpNeuGNP/JMvY6Pa/yPHofra/ylwRm+XK/DQZE
iOkEgT/0lGNvEG/sO2CUA94sHQP1KL6aPL4+yLrI6gnD1beJWyDov4vGP0+/HIqKMRuss+CrAPYi
0GCfzRYhMT8LbLSnCjfJzsjtfe+DAd7HvCzOzh2fosOp/bQcrI1v/ti5yAw5pAqEx5Spa8nbc2Fk
MMHHpa+/xSGMlR25cXIdD2YkgskyAR3k9yeEDKDQBRRij5W/QO/OphTyZIVWrOgLPb10lwm0Izhp
W4UmcV18NwBR/PWZKsbPcy7txBcGrFva99NlqFFVI30eTknT+CIDPSxupG+epS2PFAPJ1rFVssSD
7VoEEJKF6WLVvl77T2IjXFSEBNsoPgIDaQidUBofNUhMCXy3fQTeiudHpQQ6RQHa4jjHSrvaU0SR
/tAq2l/woSrCHk3dszb8OYy/ve3vL4PD4jP/fCKDeIL/zoQQ8iaMKlxVS13A1qSSFyknVdMXbSgG
5FGesg/fkkA2P3fjkEJYgv4kc3iFgsNjzhvPo2BPUu7sYu7EaaEgeU8FVjakLotWlfTmIHyaHKx8
4BLJR3jZowp6kdRPVWRL4vOkrhqiFBeSbQg6OtiXk1BFFUnPZZlzbNqyAOBFuXWr7J5JK7dJA1qo
Air73Y1+ZAl5mxzCbErtLaW2UmZUAfbdgp6bDkqi2fWTTcRTijqd74f3zJ4a7VAK1MU+6cs99zZE
zJBVFx0xEiH93G/t9Yr1A/kDhMfM79tlC8XrwHFTZJ/JjQyYDw3FYz5AcwN/P7ypxmpgd71JySx4
3a3RqUK6IIbqmS2tljZGd9+RHYaXxR+u6Q+q1/1u3wGKPxV8d3WOXWx4rKUMjJ73UcDjhuLe6F7u
3i4nTsoHSTyDMSUfca1EU8GyT0kCBwkE91STAUwl1XlgKFmKZ/yGjZwHgVdu2HyNkyOHaPD+FBxx
ogvgwnaNS4itMZdqBOXGU+KgM3HVK86sN7ddB/1Xxy6l2ofTCZp2icXqry7PQ+EKfe9eK685zv30
F+rPn9b8njq00fqSYRJg8pOtM4mSf5UG5u2XY4CmvnYgwUA4ZovK5u55A42BBJw1mJ2uy39Az6/S
9FXVqAZB+T4ckHqNyk4Br5WC8FZPsYji3LZ83D40BZQkP7TNjyhj7yU+0KRhbVgdKO86s98VuSRR
NPnix+q2e8e6jCmC/k+VUmbD5qlQHx1Y7nGowysnisjpdfsGFAMJHtT9dSrag4uhOaO/khXdY+Jj
0Nb4H6opv5adShwBhcgeAaE6q0PKD3qqd3PvItnUztXs7sTRcmyoKVsgQqlQ3lIF9UOgDDay1std
RKFoE7YKO4iiCf5TN55aVXGMo5/BGOugUs3/V8jHZz0p8qdE9uodsG4IyOqCvXt1n96Jiwcpdrif
UPjeasjW4c1a05nXSLEwBQBbIg7AXEaNHAh6LaGkwSEABpqIdShEKw0Jo/bnq6J/PGnvQgpRQu7Y
HBgva+aqo12zCqPcuwE3uLevM7bjGJwoJ56crMXIDUkd5iW7q9t0CxmISngb5JYoCbmIBE/SGDWr
eM6D6M/iWyINYiPw+zaySffDMPkA8DEpEvTie1d7tGmgve+nBZ49MZjfrkIQ9tfZ9jLRp0hLHwGc
xkmTO3o/bd0bM9R0ezjlHrZhOrinoUT3ZUqeu18MG9c8q+twb8B2mAMje5XeqR6O1GgZwK552ZT7
wRfHlRQLoAva6lI8DQ8HRjTYJhRbtuDAAUU914B8Gerp8gk11jWWWsrPU1FZY9cPFF5UQqoGrOJV
fmw37qGdTxLb9WFK1AhW2qqsEAIafwl5Hn277fLD5I5KP5nfukMvjNzT7eHAICudqaqi2H/r4LAj
JjQ0expzIpHMhi+c0fmy+97gD+r2a7VrG40PFDztgGvuE0DO5uENmbI0sz95Klcg0NZqgs4Y8pR1
IscYaaDn7Iq1c7S0VyvuL6kqsGKcJkcz6vCaOGQztCv+uJeaOn9USPKkv88jPcytYw5EN2AbswhY
vzk4xOihNN6IbRU+tBtgSfr22t+B5FZDUEAYB+dSW/y0TAuHu2JRZ8zEELDcjvy9Ze2TgqpnotKX
XWa+MwZ5fECLsbTJ7rE6q7z6ZEokjpAA14aob6Ls2fldOyiI9+UkS1vIySbXIeUbW3afqoOzRQ82
M9s0jsGfLGzoo6TjF0TWO7tnpfIGBtfToxBHXL/Psk4FQEwb8vBuLblaYk+HzGx/PGImQJpchX6F
DHH3iy7PWuXUiwgXRy52r5VBcjfMS8kyYmhU/SxbBECW3xdr3FHfyyUTR8xwfAAkjxo+kS+RWoPI
7v+JJwCmyxrs06yLJGki0ql40AteT+7lRKcFpKVtZKSp6WMYqpsKipzOw0Fh3gku7b2OdCRornNS
1P8ZZLBNRmvKdV6yzDyl6SfQeCMKVFgRDcPKSxLWZcgAkQXe1ovxxWveVkjcXfHyhi2yTrEb69FK
v6DN9MpQR2HxJkIBoceEPd+0iUkc+WT8e/qyN6LICXIdAPMStWvKz3h+1HCvTNAI4jD972au3TPp
QJHNesTvS4eLEVluKGuT5tES2GJ2DFtk7DitJ4tFzsjoIOQhsRA4nHTDfPhDpUTflZGWMeAFabI1
84EI9gfBHfBps5Vs+lnK07A6pVAlLF3hSbcuB2nkII/ykfmBHt7HSrRYIzAoGipJr12E3/bbsyPI
cgWc4mI7H2eyCXh6WWDi0Gpwb2+y9+OJr9ULPSD2jnzRgWtcCd66O6v1bA0cHhCqOeqwLgZW3atl
L75eJlsM5iO2oG9UPHo1gn2SF5ZH1+7tFJC+YzGduDnvL2ArvNuNRgFjYGZeoPmTO70dEH8Q9KfF
tStQNvjtRcl9/LFlP6jouiu3bVELWJc4PDaXfEoNh1R42+HvOJDN1jWFB0dFYscGsM9hM7N7515R
WtAtwXwSYPVKmmSv7A1Up0IpZ2FK4E06eBTwAXyX0uP2NhpO8QXW5qS9Kv4IclcDbSGP7sbR7EyP
74gph9H3alU0ww/T8gj4wYdamT+obaHzcXGL6vQN8nwNEEHsF1Ml4lSEL7KhhSB+Cy7neRTn/9JT
euBwYTnlw9dQlYYf3zffWHkTzcQzaAZ6QFAhlsNMbmpPhIE63GXrvZIWY9mS6l/1FIFz1LJ8z7dL
umCUT63Si42yzKIrw2Wha6SFsqjJRG+Y6y0hDj7eQw4GhztWGn7q8B9UHeoaKiONxU3uTJgJ8cLo
4ShkVfHo6en3xGSlcBj6+z/9lLdJTMLkHMJ6dyfgMbLwosoDgR6UMVmBxrcF6Pv1buJebwCYBNTv
phpqxUxNloQQ+Ju64gzwyNxdUh3zAt1Pk38ZhV4t9eBFIpFmxaGJNZtsiJp2cb9mZoHGHvVkT0Dy
3Hg/Cz/t+TAr3F9GjOWBAfhad3nfZVv5mTn/D+dYt/YT7BC90/DWjnRO5s9lOFdJNtN6hO2Hm3RM
ICo8UDuCit6fMxuyP8cV1V/4bOOL61tV79knXTMkDo0NBRSJ5JKNldY8fvTdtHkgNJQnv3p72Bpr
ECGUC6Ubcw98uul1dSDN13YQe+orOH6hjV0Rjg/ql07aGOw+jAA46NbkBHVrxDQL5Hxa1eZiZ1s3
eTxLojUiW6daVglwg793l3Bvz0i4eQEVIBkZBYdIuypxZ7MNepzRgSUnToxQwJEMq/k20GuiP00i
l8xGzGdZrehGK0RZQkZIYgNYqMdzhdaz93Fs/rd6/ZWk0pf7Hdo9vXGE9lcvENo+rtdmt3upPwm8
ZG+n1A4ILqFM9F8SbpvC2q7MX1fymr0wOXZYVMPcvlJtJ5VJDjk8KGYbXddfF3u0ZUUnU4WKHshe
lQCk3tL71znLoti7bgly79J3oaO5tobbpAGym9P3inzON/BojFJQhSQaGGJGWwPHV+YvjjhNp8jT
LSbCTrIOwDlruT1pwBvHCdqezbE635/n4wZaYL9GgxbrxtuKIS89bFYTETCft/j+YcatiSTPvipL
m/wuq5AHBX+cfgLYMRIgBiSf6FuQSl34+xUlddj768j8CIF1ZW13PnVAO6nDqQWu5D37JdcjQGDr
Vxy8TZhz6jo8x3R4CB0yyopoJCeVKkX3EUncbtepUBNdYJAUw1qAOgsDK2E1IoRdI1ICh8g76kmS
/5njLtMJ3XnIZKzKeJX4pWUgE35lqER9VR4qz1A+7KsVxLwau+dNb1N1kgpgwpXTuBeR8s2IXgsg
IndirgK4MJmnkWBPAYQ8BKKTjWDZ6mk7ouYzy7t2CFC0Ee52XgM7dzrMHWFsMMwp9GunoOoPa7PF
SaW7hLqROZN9K19f08em37F7nFpfEVVJd5/fGTLjhx7dZq1JpGjDPPR+okeuGfyf6ggo09emUvWm
cBhAxsii6LKPTeNp3TJM5P/KOdVNiH2DmHMPr8L/Rtrd2WC68FLswPV+blilDEUIMsgj2Fg7QxIW
EsGPSAi2JwlgA2Fg45YgRgNNaQjW0Z8/HQxngcnaqfDZ0WpoVo+KHHet/3wyglt0bhHP3NDA/1FV
c5aA+KVg3WcgW4kUTDqTRWt6lU9KH6Dw1JUx9eYc2gYmmnQRG371pUpVpBFcJoDr8hWyw/FeGmjS
UUcV4bwoQssHtnHFSvjIcE/kMhJ4kihX+k/s2nYFYu6iLntnEGXBfCUxnwnUPbto9qUtjdmV3s4I
j7zDUBXNoj8Z6ifgN25qpzVk8R7m9shVtJALt3RWvM2WxnSTpqlboq60mC1xZXlkCx5u9NkZ4b/Q
CAydRkGs3AeN2Vg/fto76LYrbQa9m0+bumd9N4aa4FfZ3YF+EPnhGIhyEM2HDEOr6gNE3ORiUMTo
S1kXGPbjHl47ySm2OIGb92edaBmWw3YVI6aWDNpVHOR3Q2PA9Otmfp2f1mOz+H61u5PQcvRmJVAS
ner9RHQJwF6iFbNssVE0Zx+3FDnD/aJXlt89MUV1CoUCa+rJRhP5P4+MBhceF9KSgCRGaIqBY+go
D4C+xWvyGAo1+pnYDxgZEF2tkmiTde2cyg/vU430Uqs7hCsrOU6lJ+SfyjmT2ZRhwARQw5rF0GYc
Cr0HYHkpHnoljclgwd9GJruGDnyPsDTl1rmEe4/PlDFSCdU2xXwg7H3HudR9jAhwEiAjZu+cx7WT
JSigVjZqYaBxezcZz9ZbVvWl77IJ5SCazVABbzIh+hQVyZ60AUNJ57vFwI0UXf91TZxYeoKflN+N
LdgMWBH4BTRizqS/Y3BfhNrNuxBJI89InxxHoafzqK7xUGfI2F0RBhV384l6hVqQWzNGvSvHBze0
xjOexFkiSmW9K94Y1Sth7AXEL3AEUqxJYZlqRB8GuQRsFJH8hmh57RtTklUYdwHiMqn4xMctCQ2X
ebl8Dcmw8p/LHQO0zIuaEdnGItH9E6x00fHY9bWq/3PyZsy7SPfyPskqMvLaAT7RpSj5cb7b7f4t
vLRVtImna8hgMg5niI5rlmNnsJDa4z2xVCICTbkhNFznrsBLZtBylLiSTygQmb9cumhi6wcsy2YQ
8APAXnZLM7ggMS5mEggX2GMnS1PNXG87mSYG6VqhujQBWa2XpdWG7QwwAAE+7k/KWSx5i+s5UI7Q
TwSWGrKf610vuLmNvRvSm/+E5TspH9GA9K0i0GxBVhpKrwJKBMViTTQd634sCVEOpqrxfrtzGhtm
mPgrayZ3Bb/5+R3B36ba2dKVnmEXJaXIOWWB6Ub3gLbTQJUAv9sQqLc7tgVmsg8YwGtF33peuRgo
+j/fDjlHXfTCg0rEzII6lEszHucWJ5aJ1U2UE0hdx/6wwQ1/BIik+5ePfdxjGgCByUnYb1G+M4v3
60X3wr/+XUaSpqGx6eXPu7vyBmAfn9NBRevFWiBe7FHqFMay5VTPJ4BwTLKcV1okC67nfrQ9NiVx
vpwfh0AXbLbq2a92W18o6ZDADryIlLO2WfaFT7/BH77LzZe4FLfHYgCwxNmLY1RcEg6+raFIcV4v
4ycqj5bm6rnYMi4SX+CiILOhEhABAQ49isZ84oiT/3c1/Jl6pE0w1/zwgen/3ppKeaahtawArdmB
pEfty3Xxytm87G2OigXlrVQZEwKs2rgL6dnsTY0XUCWkY0bxt4X2yy5iVy+xl7ZJ3wNHa0RB00EE
m53Ydj5h4Dp/ytHbHIPukoEllwxz5Iu8v4JAebALheqlHRIieQw3C+B+dw81qZhzLJcM9ZGJpsMw
S62/naKAu5bCupW/8qW4/LqqextDT+CsmD+MJxDR8P4TYJetW2xRI6nZRNAJgI+Aq9pMl0qRPV5O
81oQEGJzp+WlqdtEbNB+IFpOJGs4qVF2KNIEUs2mXKg4kvjUvSLGfFvSHKqw5gH+/ZdjcCpNdTbf
0SfqJMbM2FDRIwyc9jx5Aj0PogGs8IKkkSBE1JrO/If6XG6abVF6Z4jFPjYvW4L05KADKUfeOO8+
clznIW9Is/eqhzfKvDoozeZV2Oa+Wdx4z3uTEWuYCDVQND7NEy2sTbaBrYA4HOTAWb/7h+FQNUC7
ufJAGRn11H77J4tpeJCCoB1XHtHKpu5oUa4eRcQc69NcKQtvEOUg49CyniZO8yTwkMSMNjYzWawg
dL7kjTS0jlEOyRz1h/CpgSABzVZtNvZDjbu2fEZO0fulFZ3rhLCRStxsJ2gJ80sXRDToUKUlsXWp
488MH8ZroVIvsRSD+M/0OhxwKbCrD1KvausynjjHc4Xzs+ADo9LqY69lMoZPqszsg0irugXSSVGP
C6ZVMgfbFz/AKqamlw4DUiJBLMUZqTQUVKNQbrJN/FcGJrSidLUxkTX+LneORDc6Z+aaSHPmcCvO
WUL9oG55kj4Djn+irnsVwvWARTerMEBqJSa9g/jo63yDKgh+/JBMqjsfJlmlwN3QYaL8PhafNdfh
WqiJz2oSNjn9RTFOXgaCII0SoYZEgJ0Dh8c5Xnruf4NdPhTCsdVo8B6RGinCHMwdfleMzBYuCYc9
MceBsdv437whvCX9vKS3q/oKQOo2o0iL0NSD0Gfhsv+GZaLMSK7NmSV58lmCw8XDktRp9znyaDRn
Z5zjW23NYgOqoGG9jdqZj1zFubrcTeMYNM4R0fbfLk1Lsun9DlE++VGaHkuIiOgeulyElUc6Zis6
hp13oBDbtSKv7H+p2TvFS1VPiVx9HjRT7/Zuk6LcPzyUfaNvpjBPFHK1kty6c0XWAYVPJ6QqEWVF
/2uP6dU55g04YEoUnLtims07clyJUOv/IHcf0xXTIyyJSUT5P8OPRkT1QWhT9bSX17wX3ZaQ35X/
XueP9kBRE9UPwOwOFipEOq5UL87vET1wVmPMGGN0eKRh6+M4Vfzc8Bf3DPxLJhZrTy0swhDry/JS
dHoi8k4ios2R8C/ja554tQOjYc9TCycbiyjWCz6UxjkE4ePAmDF7vXHjJLVX2L5p9AbzylWD6Pl7
O+EiII/1A2Nx47RIKm/NpPEsQit7gQe19hdC6D898DOk00lx80HVnOiR4ju3Cy+TbgIpvuMv3h5U
Nq9/C2MB10s64NIjqyz1ekdW0JQ2tnBwORaDOxZ4yAFW6/QAbu5aezWUGoCOm4opFIvOkT7vbYpq
EOUp8NSeijJbzC8I7fbVM8h6dwnqYO8AiKQmu+mZKLAPatNB9ywpJR+vAMaxzdMbmFL8EFqpt8Bv
6/pYx80RNGPuuZcEeRjbNan2LJKxTtGQdxD0UU01JwNaoNuxkSewfJwwe57y0ByA6ZM3LZyaEj30
FSUDAaGKD+H+7mTT1KnVQaz5Ba/fcvjuTMqGKFCaq7KXriVl3KmcKFSP4E7vXPmCCqmvCvIQCRDk
vcLVS4Adrelw8efcCDQmrn+huXlHc/ER2cDzxb31R2WFjCykg6SwmsqyEUNRxWmdn82zMmFoCwal
8lVUvgkvpk4Soue5mryBbZsMP2vV0R1YlfUFq9WVK+0rzu3kyTamns5JB9va9eFjXtg6a1uewtLz
1FXFlCVNnIJrrakxuRvMVLauGvb6prqdT/okXDYnQP877MDPJFCeim2UlvsYdZEvy2LhTUaoM5DW
Atk4DVLyUhtLhGtuHAsp2ZBrsDgkt4UhUQugiEzfbvVI5v+u+uuuupir/dincgOthbMhkfshLoAI
7RadE9F+/BZlj9HHULTutrsVpAqxUTK2O/Sow6NQPfVtshT7++ZXO37APVmseL6WiassIG0rNPmN
HCqqT0c+LJpy9T3DI6iPjmYhauSFcuzmTkNN6KeTxG/XepLQgBy/82QFFp6Lv7fzoMnrwxVSMRWN
6iP7sxfMQ9XiNB8iLuL2h61KYZp76xey6+D53RoFcudRQRpCNf+CCgS9yDRJv7NbWTqVDtU9GgmZ
lHen3mr3Lw38AxQwKzb56J42yj1WJHdA1Pwe/ybslZu9AzkWDnrnXvOK4E+8xs89bBPR78BOR5hE
vtCXk7x9Jo/sb2vowLssJpK/Oe2VH6bsnQWMZ9DWPG3e49Am9C3mYIGRjB9eu7CuKCnWi+CE6jJ+
uV3BxjpJkqbljTtpYgggZRFUhyo4M3TxTSxJjo3pOYHoTTQPRMV0BfVECs1JeKxi4Z7rX6Auqbxw
Xo6qnmEkklzdETxQyB+00tIdnDgNDWVXn571rWvPI2/Joy5YGr7GqNi9lnwz+Fw4HvdQz/ketwKJ
cpe/oHPPouh7mCbrKrQBqWnYKKcgAF0s4RhfOy7xEG5Yg20o8T560pL6gVBrGZCY6gSBrZiRlrLb
PnwkJrlUsLGyHY3OX5T3ax//5hqQlVKv+FhSfC4L3gZDA1cO2Z4TZ9Ha2m30ulzQcnrWVNXKBLQP
sRZjAs+/wBaZjPqVyGbmYlo9QJa8hdzHoR/aByxiPw2+dFZAxCl5r5Qlmf1QhVSZhEtrjjvdw2fR
63Y/kfRN2TTz1uRS+f8diN9etzLxLt8lJVDRsJj+obnh2gZWXnKZAczODRx5pFgUpFCONMgWedcQ
CKt4dKiAzKmYE5DRAzk60kUVTAU+/vu1FyEHu2VgEMsWkz8KOSNYpk+d/atEYOMQedVbRtbX+6ih
16EH0jXwQWOO5pGWEh5dAoPiHFaXjD4iGdFjPBQm/uHoMTrkR5s8FCO8xlWAedxVp7m9e0C3vgZs
LJzc3dkSC25x1XCMC9m/qtNn/COacx92yTT9J/12K9Av83E3SchMFJrd7vYiwFIUko6wv/wKL4qw
EAlLFNKV43bbBuEDZLpzh/RWv3Pdka3dgDWhrnX7qaaH9f9vG6+EzknwL9v0rFs/qqXGNWmHWuUq
NDw+jWUrx89DEWjkgjxmy+o7siUgMXcv65RvGPyjzcTg9IdDPHOF0aO7OjySFpmPO7TsL8ZyqVge
zum6ybyKjzqCpArTvoRLGxN44sSrlq25CYn9wkb646k+QegyfB2II5cN0qmPfH910KpLPQp1H5NP
dbRDfRm6Iij9jhTaDtjdRD3JA7P699ayJarOTDgD2+F/Y5ZkRiT2tZRMBmUzZ4C6hTm0yldzeYeZ
8z+Uav+lOL8SUA7Bmz79DRl1SYvD4PhTj8V6I1iLYsEVjds7tTacHdx46Uv4qEWVsFTbLnPVnQVm
b2zYOLEBM3Op5rBa850MYi8mECwCo7O9IZWYalr9uC3ECvrDOVjnPOT8vkUW5jzQ7Bw6Uy7gEqQF
DSmiryI+zPEkSsoWDAOs21thrj1dEoqMjqwGsz+sjzK6EOjK9rbILqwDyov0JqvxdkrPRtxco9zo
fmsTQzq1eCW1GWJsqpFEshbN7r6fkoV3JW4nZmqzzYumYheGgpLnTavYbne8/pOcXLJ7KsMADOF5
bOFgTNAo0VnGAtg0Pv9ql1s8EHhj9UY8yeCUWIsCWMhENmt0YHiDVtmX+rn6bxe+9wRdHDsE0pYE
3a+27vg7AFaqrKb04/7ZsFG5RXBfjIw87vl/UvhSihrMkTcyWP5nJ5YyB2Zs63+3Yw2HppVFTXQ5
OaNpx8lW/k0GiAdn/ynzO/jZrq3+ssG14vqptu4oDZcSPYWUHCNowzDEi3QiH38VprbXpa0TpbZu
Mpdkh2HXYMGzYskhqVua48y+//AIjTQ4Ab65CBKQPjpYDZ7PPpuXUQlfSdhQ9zn+Q0djo0ZdrBdk
9ai3bTWu/XdSABDaHgJ9ZPoZ+qLUMpFpO/PG0/GvWGXNj4zX4EB1cpzo5JWHVPIKL3T17djSB+My
+rx3r/GsdR8J3H6EhWdMhBsspMfNANWc0LAo/kOcvlEcOqihsjf7/7LUetRHP+NDfNmK4I/YtI+x
oQCdoJS2vhmVUSK8ssiaVyfyrDBWxUdRzmM0KZWkWFH+sWHq/Lb4FOYJKdpLLXtc/bmqkHJffGj0
dxQ+QxKXx0wTeuy4avymWCR+Vhlm/GPSVv0+Cqbixx75v3p990E5N+P8gsvBgK3VaH8hYnS4hGFb
cbj705slE6VeUuHa33Ic2rYtF0HsJ3+h4Zv9PVK0bB8AZ2Vyw1hikV0+m5QNhJOVhCzuQKKCZFK/
sf2bCHlD8L5vUmh3d3btsO3I7CDaFSnBSo2G57FNOBTNgpUSJI7JhEeP56/dEscEpSF+1wnm291H
+ooIXSJqrPo+lUoUMSo53atqtPm8vpe/0APaSwLH4OzaQYAKVyyw8x8J0lT33rqxgAPsi4qWExEq
0ekuBPY833YnE4fnbH1ZeoY3O/JNSenEVzQnmYOsJPDUZNrDaXysUhpB+H0FFK0xWr+zz5ACU7/c
1pqlg0H33rxl0xE1QYZE9A9jgz1H5e9j2w4bNBEBcKepCL8ueFEw8Fbe7XNLF/8edH5bOvtwo5mw
ZdLuUtkjF0AnrtALD8ioXv0IuL9b9WGx5Ep9SnnvnMs7+cSWCOFLI0N71lcLFWQQVNvzf6vTNzoj
ab2S6zGJanEdj3mRbpjkXOUu4unlwfj4aXs/J4DSW57HKuAhjmFSEScwMDOAQo38vApeaq5vWLVH
XdHaBLrT6OHirckFP5/EHQJmzXO5h79qzZz3MJxzGa0GaE8i1XdQ6+MOLiXbzilQ6DWElytwRIfs
GeDNEBcTEQTI13ryR+gybWphwMJ9NeKcxTsSl8LlOdj3tEIhR/2KAQHZ4jI6ZgZ1oPYttdvWro1n
47KBJMMAXJJ046RoFPmR2lQXOLk/I1xsuopa5nmVQ6QOTiMEETxHjQxwC7RELoFYIVjqOZRzFB7K
kY7enD2wrysGgCIaWHJz94luNdPNLxb96aJSY9n+BOoR1VyeXX6b8ZIwsP2RtfgHYZltS6gCCm8v
vcMSjEkIi5jORhIkpvImSP2sARRvmn5oJXhOUGwRmsJSg8vNulak7KVq7Ga1OUah+KCaZZoS/CSs
7VYFBHfIUAVoFH8Znlv+K2muguVPOl2hh/C29KJIFw3dg1e6/JePpuHrFzQ/jRHcWzvWUuawWePw
ifQEXq+ouoOv8O5yqg15BZ8PvfHokQhsnHzCG2xYfzP7pJRbAP+Ig7fALuLEEsauNMBUtxvA2mBN
sw8SKCtYOuM/5JdDwuVBLJwGOLMzIOPGLdH7uzcKCbY3+Sx3LGY7iod1uNITeg5of6MCHFCID4+d
5kThY31wVQmKxsT6wmZRaaGE6C5zpuEkts+Q+vaQrOVoWqEAw/FwtRr/SLU1XYmJdHkG+xqwJodF
zGmqU6Sf9fgatHkKctoWNxyEaTXPMVDBMTTpPrZPnvxPXvlCgWkBKAcsZzmRJ6vshkHiOvkBIAAI
EvkUHGA5LhNiKWHml0IZaEQQ4K0UVeK2WQEd0x8N1seX1Dh2CHNLhghV0UzYweQzDA2YFQeA/yXo
eXRGWY43F6PbAxpYI7E4p8y5o3Kn0R0eJhs3rDJQ2mYgPb0AZLlp+5rNNl12qJeS+nidqnglYrhT
CJdoy4prLDepdZf9rfzWLp1jaVYSB8yEWLf8866pgh5tWZ9UNYb/63b/PkKczJN9iftOYLbFnIis
0sfb7LR76OHDHDnXTJCwDXy/hI4S03yP/mi1qOGyE+XqK7N/L9QDyq7Bn4t2oxAago33UkyHBWVd
0zF7dK+QbAhWTbQOtQsVKy5bIfQMN2UCIpV+RQP3E4MFnpmOXkZipHby2MBHslJzUtzZYdeHZt7U
Os9c3Y4B78IOh/2BSeLujJoM07+lLhO3wTAOlS+nIoy+ABZ08Cyx5UuQgeglLFD7xgNCaEcsiPxN
e+ii0A6VmhRXp+eFSlzdFApfqV6HrsbcOPYb1nLSJXihhQqetaRME02DFmet5XldHXTEotJz+fws
k/qAbhOcPCv70Y0JmO8Q8F9ja3PeUhHGUOGeVxRGyrBqC89fwZQZ2l4igqzSXeixAzRfk85TRtWl
46blndX5Gi0DvIdSgRfOHj7VzapGt82xXRvyr+n8aFl6QrYKM6N/+jL7H6nonzhbhWB/yPx1drBp
EeqK1qBX1G24vyx0rPnLZiIkJYpDjY9wts1FGXHOfUWlicuhQHrr6cNiVIq+z7Z/pnIrabwq8U/0
WMv6Ng7D0cNNwoRr3cTNNNFLssRpFK+rWq3j/Jp+2Cnm4b1unkVIRh0FFO6VAV7IUMNTy8oA6gwK
azkwpZX5e7Rh1otw83JgxnvnH7QpyXal3jdwdAvxdykauBoNSny+UCVeV0zPfJR19vqmNlnPB1i+
vVxrBCXKlPzPiNNLhvAB4BmD0RikjLuxcDeL8dHeGr2hZufACFQJSRutVikNt9es0Hzk2RuIf8pJ
/ZAYQ4WaafP148Zy9ns34cnPFXEuFYXBUN+VYBwyVNbBNjLZDQDDk5i1DdMTexQtxMeFdh3i3mZE
WMPlU7Go/YOC9HLRQqG9DQLax42ayzCXf2C4wcquVtC0CWpld1SCDOmHUESG3E3rPru9FQIO5JDc
RcnptHdPLs9dKNBaQg3VbV6013Hq5AZ6N2yvxZFoYZStAUInlKf0MTb3PmkFQrL6hJYpoloAXrIP
PEyKw6P0buNVy+7oxp6sHafAKEaTfgdLtWmh9ErpKQqvGAuWdmvqAnWQKTKq8aj7jx5TyWdpmt2N
Hp9hw86ev0d70aNQR1KKiOWcGYfSRPlQQnr++520wpkw7VDZeEimAgf4mHfuQHME9DQ8KJrYRZoM
1krMekxPdX30fUmt5sICrIG9G+wa8MNIdTMSj3DcGpp4FVHAYfIZxBxOYT48odm6fjwIjdU/VC9B
ZPbXmDGrYcrTBVO8Nv6FXvzWvMM7e+jTzY687i28daAgZpRG764yb2T/88vbVUEApYkebEov2oLk
S5I/NPeu/lnXpdgArqrBqq+EZF0Y3WFmaU5YjKTUWFVC1zxCRSkskjeqDV717UexMvbskI1OwIvZ
6EKeGRfQrl/hKmOjYv2h9ItUxbPXhb3YH9QfD9h4dvy4NQjttSazmYp9AFEgcMpYmBTEipqnjesC
5Fls+639CXvVwNlslIbEGjhLTbpLHl4hEG4n4CYNqDVeRZyCViBP5GDGiZev0AEEF1FgPy8oMsjH
FjAU4YqGduvXVx58vzCtQiToy3CZuY6J4W1zYnY9Wv8TNvwF2JvlWzz9hLHO3CS2d/crATn4kxjc
CfKQij3gXrq6W0LhPagT3+IqQxgHJ+OI03qBiinUA9na1/pwTyyvSxCy7Q76Y58DMH/eqbPNXcAT
yBLO3l19EeQilVq6CWb3Fx5BnCeFMCIW1iuXbmW7dFBzQMy5nvLwvBeVfDyk++iyBugbgRIlxYrZ
Ss7ms8QVlR8uESJyl/8yv1YtrrUrkfr7H3xV+tGs7ndp/IXpZrONbYaRcLQ9uEkVVz8znKSTa/a6
rFmN1kRvuhQEanLNj0em42whUbhssD7WBycddcpuwo/kIwVgjuyA5NXd4qXs2+I/oRHYPc39UCMd
r33QJxzR6Z9sB0HeYL10zNDXm6Y3fWiK5C8WloHVqbUFtVr9RVUZwKGXELjv5e5E2jWP6cdKXeF1
HOw0wBQ29iGl03F8fNzYcoLJihGKl+4/p8mwpRwkjeAtWsZ7kVsq6m00xB7u6E67i6rg+Pocepfn
wj2Y21JdX5VR2dp6I8m9PwWrQhhggRunqvKVr3m0iliGdpkSSmMgYOkdXgj/iGUNC7w5eNlzuly3
L6m+VfgKRy/iJjQDDDjfAhNqyZG9jo4GDBtAUcHsODcD/gDd2A16dSNQjvYDFzIUZSxKCJWeaacd
f8I27bI/5avxNQ+6T++qxrJHmCVI55yRgJtn7ROEH0fmVWPThcrDpT72eVbA4GHXb8E8dOMPmwy5
sn4mZMoCVhDySruGv4pP5e5IkMykmDbPbgAMrUammdTW0L0tM2KG+cd1r5HnoRh29x77V6gTbopT
xdhJn8/8ln7AAI+xwCFsXwARR3L7+V23WnayGk5Vj8ldi3pq3n4QAyb7XYxrj/2i0bEawDlkQC7R
Zz3FRtJhrP3Dedj0Uy7Ryl3rLU+Wp/TnmNtZW65Odl7HIk3iaFA0sUYiJgf/Om3RUFk0gUfWEsDF
YbOyntQBTQBzXhQEo6ApDNz3pgK9Lx03tiup/h2NpZPrDnmIFN8GH+Lj5X+0JZPh2+oawShVM6wO
cr0Gm41yV7a1ItyxnQTE31nL3yyHFMOpoTP87QqUoi3KszbWjrLnyCVhgg/4b5fyrSNKHQOmcM2q
TdulAXcCv64L4GQWDIXsdY+VBMLdLpOFlDUa/FEsZOFsSAVstBdJj9FNOIod/HqCKXy9bLhDv/jJ
sLvkE+JxuNPcP0qeH/dcYE35zjOEi9RJPycFiWBdF0Z4AjzW4j9EWEKVrjvhCipfX1ucfuVjcmaM
fSHhkjqA/5MuImXf+1hk9xoPPyEU19QeiMWW69D3uaS1YWm2ng/ud7v0ViuXcHX6nDGDQK6218aY
dhh6AhDsX5g9nS9iLhBKokfnAbrVCixArqgjb4n9IaOkrW/uioReMv8Bwq+zfzFxacqWHF+uyYim
a1FA9OHC8V3RS8Fbt6VDUGTdNtqfl51BdFm3jgFNw+8ryq1cDACLe8RpolxnscgKy0gStrpnTkV9
pcMXgdET908QCczNovfeRkimDbsa5swnE08URrOjAs3Yn+ywBTV2J0r9R8G9jVzt/H4TySgJAvon
831esT+449JaAW7xBZ7SlW+kYVuWaciLeh3DxgbBJshP4GfbqpBse0vd79Y144uh/c95xjryIwDs
mdzqGjvEuJBK3E3onmrHWPUBgHPZq/49MYKHHpZrFiwCMPs2EAnTgj4EFd0dbUlgDzQuk8WkjZfg
UsLZA0pSyURvJzGORTGvgxvdsaIIJTU+52qWgZpe1Tv17/+S06+4ZtTg5wrvrjX9+37BBznMjYMv
0bqD5OF6zQEX7HO3rpo2w54K6pKxiz8h+/uxFrg5QpR6NCwdSRiixz0JX7s1k3qXcgxdLGg6hOhx
0sBHC02V0aWGFIT0VjORCjQu/pw/x7UUsagPq9o2CardQ+Y5oX3ZQNcmyqMFakPjjUZxI2uE8lr4
Wtd8YIMdysqHBL9rUTr0Ai6SoYcgp5kb4Qmm8gG9hbCS04Y1gENXjaeb5GfmWhpdDcroBLnTVnQp
ygxEh7yZfhTj6HIEuGdF3EqbjUeGzIKF81QCN3KNgfl3MGc+MSMghGCKfW1cmNaQPQgDV7GOELhL
GyOcBu1AvivdhhBDicGOE8suNu4TFO7o7Zn8QtHhTmvbPLuSzsxIbaYYPwyRla0A29QSeawL5tFy
joQ1rFG/eLjr1wDeukMDWn2uJMfkXLZ/Zm4W2Z+va/gDk6/XxRGRYSpP6B9vEd4Ec9eQ5tuLJOba
656bLddWjZOvSuEP5UxLPodEIQozDWMKBUPzi8siVg4BvPEKnsExzh96YbuO/gQ4+MUX86/OFG1c
E0PFxLBy/baFi0dw2pPuz/lw75O+GSJ5BfZ4/u+xzphSVXxQSkJdze9Uy/yE5Q5j5MOTPgwMmCfE
W43/ND4ysQfhKCIvcsN9hOLc3mmn8ucqgR3hVt0Hpq8GwH/AK+xXFf4rppfamNKR8+Mo2mihNqwl
hO0J0LnxvjymxNYVtZQUC6xum0QgBPM9VoesfU2eyWmoJLKv91KEr5yIB9oc03o+NyGlsh1iOkmn
k2QQOwpGamHppb0frp7hV0XmwrpHuOOpA7fjonKk/givDHKKuMGbmw9wmM+n+NDVlfOGsezyeQ+0
IXzZAgfVxhrLQSE1lrfDoxkP/dgsbTHa73QkoFdNchobq90rwmothj9TIEyfsWA6GVQMCfPIBQWh
+/P5mEr+IogRnh0j/1rw6jE+jm0I33U9UQRCQve4oVhtJi7fMv+yMnA9vA8P0/L6R0pDTbAtCzrc
DSfS29f/S5HkuftXl8uplAAHFHdgq66+kbbF2VmQ6JQu/Uv0s/2aFaMZdBoMtQ5PFQqTjp9Xz84S
mULwD2jJeUauShavwRWjc79uZcSXG+UwjW48Qc9P1VUoyApsAfsfEWWYjt0CB+1/9ObEPzgKhlWm
pL/C6HqWXh2kbtv2Gp0OJvKSw00FjoG3dlRxQG5oSx3m8humxdGKL7azjkBI2nMeKYlh2goqJwRg
1KJmcoDkj+mWnnAvFo6AucBwVEEGzn/QaZxwRHEnU2bwNiJwV6tm2ZO2Hm2j82/uaBInMvhfllda
/0uug9sXOWJ4jUCXjmAOP+bXm0ShVm+4UpIw9OaA4I9sThZhWQtnxCokeI7QfKq3Fy2WDtVOxayD
qVEXpYmACsbqBJkkUJRpwfUlQz19JW53Oz2nnh1bYJ0yTqexhHp2skgvfQ9VUShe8wPFOWz8mwks
AGumCNEH2okB0Cno9M7A37rIemhs85P1fFshLqRhYtIuYVkmwVmOg54aIOWyjS7HEBFxwF69RHco
2okwV2SRss23+m9KK2f6/jijLTn2Qf65RidN7u7v4P/5ZEnCSfXLxnFjIqPN1vPL3SGnpydczoJL
iPVi86JJn2vmE+hwjR2fSddJ+w5Nd+69yzLOoSTmWW5iEVf3UjDS8Z4fnqEYHIslvqgN25ZQUiNj
VdNnsFtQ/bjo5ABIlfAwetxVxNeO7qTO6o1/fN2fRk1Zx9bSGWlnLTK5rE/phvDu9WvpGhL0c8pK
lozwQqHY2UsiSWpE+JRUd3BzKz7hNnfW8pnfvjx5ec/4P43uaTki7TgimkpKsXqpALq+2SvD9Olz
OXz8WkkSlv3l42wpGmakm5Ji6GjE02vEr7OdLN9sMEldQtJGCaB7hzbXNdiMe39y/AePiGNl6VsA
uljRdAI1W2MLENiWeqdHfkNdhEytH0QGBdcAOQ0gcMEOAf+Ivw8VclhamFRNYnaZHV6O4/R73J4F
zzyFyD3S113WH7rZoJDsMUoPQjJyvaPc1mvAlffuy2BPQkTETGSVS+JI9ZfYeOH757SfSQTSprgG
/p23NSIohHDxYJBRnYkza09RujzExYhLVNMJji5ZsbWr14RdBmaYDXnPqTbmwmw1sa0j7SXY2gbO
htwyHDCX8YZHpt68D391GWaJfOzXYz6fREhSVIMW2B6uWS5pMFcJBumOBbSaRO8bWKIM46gCU3Xm
oijlO2HR+ih+sXUep8R6T5qDoMgpEZGlToFjvoUD/q0RH+Gf5iuywbT9q1AGaysFymL70ATC69t1
Yjt2wYnEBmjaT41jVm8853KizALZW3c88QRkIlt5wRJByst8GsF6ZDQUrtcxO5YnKTVabyeaVr1f
0fuRWJJ1LGjaOrqsx7wtdKc8ey5KhrJalB41+AWDz7xCVgtc97rq2GAVbza6c1eRNJHq24pIr0Bh
5aNikpSTqMUCwVeGuGaJv0PO8FrVZIrNGm+vh8xM8pPeRsO8npPXpnH0551hxr5UY0BYbf1pBMbB
/wQ3FAkIFxN8C+Disd2fTr7eZRjMyQ7FMcMnEQ9ddiDqiHFzb3gbcWJJPnsibjQjCi3H24iotpIc
DDn3Wt5WN8qV5pZEtxUf9LKq6ygZHVhU82MufIhy8/BU9HpyWonFTnj7SmBMR5qCJCobRPR2H2Yr
L9Jg3ji56TPR2lFNGITwjtQzEjvZOXArTfusSipHnzWlX+uS41DqjTWur7tJi/idcVhNE4f9ysEO
k93+rPG0UzsIgbJpmM1RcMTjybyOapOTGuNdSAo1X6wMNvDxCOMQeVBUF+fs7qsxHxHfZ3iqnc1Q
I4SwY6LlmO9Tqpgv5MZv8DbLJsgbLz2SH9WLCoZgH2c40OrCKQ+oSWAUapbxuM+nFMrtp4gPgeAJ
NbimxMQtZNldKypp7JNdRwEXQpIykbQ4Glrati1M0jGDXl0mit+OGHcWsicffmKqmXRbU4/yC4V3
/KRhnLAs9lDkCKhMisGOUEuhILBLwl7n3Kjx8aiU1SFYiHhECFiGZfIC+554nG6E7Q5LYt9BZ/zE
DzfcWInzxW1XLEAdDjAq/T5CgYkueopRlqIMgxBe3OG/oMf7DBe+kK0Zo1TiUe5b8hRFk00ARzXs
NaaChiR3ZfGPOSEYp/ew1fRjHS3KIbzvf+uaYtwPQKEWeDip6lbUY+qRPC1E0+DTsioypPM4xeJ0
XwSqLqkBS02fZUcJVT3Ls4CotGAudP3NRW3ZEdqcsi5VmXyO8YNsIpQRtpPhxf0z95LN/abAQTDV
f9LLw//wtmrLdGKWVpZp2GbObhqEEshBv4BLK7VHZoGAUp/4ejcEltUgr9ypfgvjFkJGE6FROKKm
8YJx49j5Tcg9iZ5ndq+dW8222U90mmU1aZJnq0JAFJmIHk+AxfeFbVhHgp/thNePBw6BPQZN6VPG
9P/BsYbURX8AyFoQ+uiPYSpcaqOFI8nlxHQIpEcmxueCGfzyHiadV6I3yF6cBJK0yh9MaFuaKVq5
Fw9/9xcwsURGDFWkQt8nDvMHu5qAk53Y/S7Z7QTq8uLBD9Z/NNVqMld7Yw765ZdZFuztTX+o7hPu
i9f5/FBJ+s0Rs5n166yYS5gzVIfev2TB/qp9KU3l8j4AoYiAreFvT3AXNlat7fd4FnRpdM8rRrUb
58n4kg4w9SAie2j2AzE5IE00Uy15vIcplxJa7a57wcGmbCbfnXdYLXjaIMj/7LyxyhZDacxgymjM
jpexdG7SzRu2vcewMWOI6iw5DcslK0tcPDX1aVI/O11V2nV/AQqGGihMbD/+uDTRPikXM4yNyg4X
FhUnL3CQhVcnrcpc1qBVHnqEhKw5DKVNtBC+IYxqM8AOOdYFQOJ6x7h/O3SqUJ1cYJrrumTLUflN
4wlnT6Nf2fefNrFHG3leISNOW7Ilsj/1rbjqzLyr8A0AbqVX2p29x6Ssjx2kaf876pfzehcnJiK6
DEV7j/01jPdb6l6pyG40AbEFUx5Ajw7ZFZT7kXTokkFHZAff/E+7K1AG631976RWYr+Dh9nZk83R
wR/f25eXjhtz5JYlrSEqq5tbod+rPfjBpA36+jdQbbszRv8lGB9qFx/1LwfbWor6SJsyZbbzGKIA
HI2cCbUtM666q+DtmtpCSLwxjYiUqvG6JbtiA+VS0BmNom4i6CX45wShnCpbvu2cE6nmUTWbOboe
wqcNusY10golvlOYjNiDbCCxTrIYBYq9GcxcKBP5AmBQAsspXmNsh3ohSHkpD1BkJYn8XwQ4kDTM
p4QADvSrqNTf436LtSFiXqaGmwU55R3pcxLLlyfCe6eLPUPjVExq+ZB+KQNllq6T89mP01Q8cD3k
8DxNdUlnC/tCHDT3uNHMWeS5mknR/bK/srL/kMxrnTtT3N7vpNXVT89X+ExGT1VIv1765x3PMvek
IKaOutY4WWiH3zDUkf0MiwV2NJWizIB2oe50vd+qnTPo5Q1yOyVVpw7VrSdEWL1rw03hibNHBXKs
BfNX9P5WZwNvA5buSQ1eJkDGg29PN2KgsMpmB8dK0mXfSnc/BgDXNpUA+bDazlk+MJgL8rby8lLp
Zh74V2EeW/P4P8sLJYB81kQH9kY4zOMGS5FlRYfjJfACy+L1MZyb4O3ktn36d+/TskSYlE8brwH+
CrM98puNzS3xEDh+p3L3YEHoHE7TnT64Kl64T5UHr46VZyQ6gakmkVBw/ynoZ2I+sPWB7WgUnW7K
h30l7JjXks8Q4DdFSKYx8QviOIIzfX0f/rTKZXbehnpt6veerHwnMG8R+lRyltmY7hISeyVu18Z+
j6OpQmAUBlatHSEKX6xCFu6OuTXxWT1A6LKPZ8M8uWoVLEne3ajL0kokSf5DXiEgoIou9s9+tD6J
DGRgZ2bVjKfHaHbE2pgQoChdcwmgguDAvIM6VqscS6rd1uzvspiPg+92VIQE5ULc2toAwsPbKYtz
SEwx+5r/7qRiUhf+Y/FekhJbyH86Z2G4V9QCYzCWzFkX8m1xiWdWddf0Cq+B8h83wgwOGhsPp54G
h5JRWajXHVRsCb6IDqhqbq3s8U3x5sPY/DjW0ckl9uBTycHBqKgIHlMpctUTGaQrkrdEhVS7Il/2
zlwEa0lCSJ/vNBP8qtKe8hm5wZ2WV3/SgPR9dI7In4/XOfDZhRfXQEYEx6dxLN/WeB6WHs+mkH+t
C8aaImCPu6RNd9RhQZ87l5lgUHuJLi/Li7iD/uocxnJcqp8ort864x5cqmHNxZ3K/DaUGyej788e
4H0rsZCZ6TxOQNC7LOPhx+6ddVbrIh0t+H1GFlWCnj+FyBogRkF/DvbyreCgq9A7EKC5cTRn81GV
1YfypzMIIAncywMmDayMRHd6wcysUmK5QDvsvn9Zj4vIvYsQg2AIbM2LgSIhvyM2oJ3gW0qaTpa8
dvFZF5Mp5GkUFFwBFFWNSAbh04XpftPj2FuzeH2zfVCx3ECLZquLoOI0xnN6Fb2+MFWHY9AUaZ5E
sFID89E3SsOd6EzNXDVJ3VR70IO3rnAFSDYP8y0bsJ4lcU2+BFtla4ELaIX24josBlwAA2BNcnng
1abPPu39a0nQUozDncJZw+pNcZ8eh6gRWwTtox6TxQifMW92gxKEoI7U0+5v8xszda8bgeObjoft
6dYWQ/2C6i3NKGP4D8S6KXOy0YJ5ozVTD5HGCLSE+12Diu2wRBXDdGSmU9tP8rANnhp4l7pLjNYn
KWVUhcSTiLheH2mc7TOj7A9LsTfzb/JRrqxdszoLROnGKmOswYqnEJ53z2GsvZmx1gq4u9adCo32
tEyzVyT8/ANC3zq9pj+kO5QAzuJMRuyEtyG+xwBu2JZOHNYra+QM2BwetAQN9RP76Pn9dAxSszFG
oENY0yYKT8ZIaW2KQWMG3ZoKLBV1JtD6bJQFB+vkWct9iJtzlSy4BHcvwc2PXRSqWSHCCjIjxfUZ
nUkZPOXCDHTrNUw5jqhVZgbj5JFT3GLPBiuepki/76uwElDwH6aP0EZcBvVZQ5FCTRZ5UhYOJ8b1
Jti9jpLHgvQnkSuGQZy8nD0FImzhc/rPhkI8AoIsb1E9t5WgMzWPBzuThRrKiycSzJ32lf80ruwW
DV5YZNDtAAyxBQ/mxTn8bwbHKclGVshrtYHp1qf/qsZqkq/wBF2R5u5r8+Cb8BB0Wo3r2uwbkoPn
ieJoKTAYxSauZEw8njyORb4PLzf0dBKk77whVQLEn0EUt6L6iVTgEBy8DK12peia75LJickZMW/R
iLKhdSn+IaAoAzABLF7q8bJF/tHCOt345gJTRFzl8dkTRpqfMI2/2nj6P08RmPfeGaiFwyswNh9D
8Q/6rzwSJTcLnW/CwhGBe7SbjpEIQYn4ha/f9VoMVD3dawm7dUiyY9xLst4odPT8mRnJbL7VKieY
1gsudhPJBRPgulHwHG5+esFy2yi//jE9mdHXh4e6OePORyzzQjU1pUSp8197FaDkd3ml3XI3J29E
gDrcV9eQ94+4UenZ/+dbFIUKCcF7/vkn21O6v6MfXRsc0Rk6VeE232rkk7X9YwMOgaGGNhlEENVF
fu/4nju396vHuMnBylZGjHW8To1/ivt2kkI8aqjkiqWpmX754AXz4ct5//uFMfGzWqr0YRdtE1s0
2+6HCRK9DYKRDBvjyD5tJI3GliMrWgp5F0adbmEJqauCprD+oAE3RbfSDjEROuJY9CXJFMVR8EOH
cKvJH0dPzN46SfHszplUwW3VIfyDbu5g0+UTtO56pdAN5aqT576dK/RlKnyhZpEjRUehqAjI2vr5
s14yQBFH0rlFkq/2H54qhkVZZo7e1xfTtM0IzS0ODCKZoo9756S9tMxtTpBqHF/f9CBHTVGu10+u
n9j6Q8p1o6DXbSwpBaYYpmQKt3FNufZuWt9RlIGnyaRh0KlfrrupK3X2p+szYvjrWAOSU2C8dZ6N
UGYZMGEpzzMsEV5D2yfaLFII/uGDh3mWZognbh8Wby242lYEBCJK+PiCF4t02Dg0drTC2Hokxe2y
NKJJG0vS5fm1+JELxlAZVyKYr3hU4xvpYED3bOnmBBWREoaPXHlGHx/Wr7owkqEazjdWauxDxbNK
7h/0lLNxGtcFAZ5it2j7uo7kcKTVKmYt4/Ni/bhnRgTxG5lBL7RxSc5JzSk9Z6aC+c4Euiwy15/5
tfBlhXIW/CYGZly0wvXt8Qvc/T3hAEn+bdGk4ekVHgCeABrwl+SwDfIBCv6ps2bpWjA6ZpAS9HQK
xIjQrIABIKleCociRleRMA6PT7c9qMFOYQVsCL3KivxSLr0Ke1qf1ue6iZqg2NeVQEIb0FRE/NLr
RpyaOVe+j/f0KyIbJ8qRikz4xSCt6O37wAQ3B46y6NayDkMRUfn2mswGoT6SZJZ+T8f/QLIfTx18
aYfs9zx67DN16pcccoFDWUqVhCceyn61ShmZwta2+VF/1mgxwcHHjcr8/9nnkHj+RTM5SNDWMvOK
OVKpVsYsdxpNmsbluPFqI+k0qaQCDI5HTzNM+zpzjXwfbqFZqzAm0a1cES0O5miVSSMPLzKzQlgH
pAWHI4617Dz02tNcdEj+qfkSN8LP7Azh94WEG4+dkgJss2YfOcm/RFqYTMrjGy5E8wbQfCVuhnbq
Rho5elRyFZg+04ovhDSPc2/TrAAmdePYa8VCMu5/jbPra50oQIYXapvHHAR/23LP35DS9ly8Lp0d
9B63cTM5mlDxFUBgViKaR0M5wQM5GlCZwMpwUqC9n4416sLgnhsgdZQ6m+PgM/24kkDrrKe66brj
MZoyFid33aUWJt+yxZonUcXixvwvtitmLxy9RmPpt0VJXz6fGJ0HkRdWUGDKow8Xadzedbc+/xqw
MTLhXmAxZOvAECwvVUuQh8ECIT7nETnD0c7IfEkQZeZtVr2dPl/gJkwqaL3Pfwoiu9n++KiRPkDe
3dI8TAmHxlgXn4hfNLf4dStAHzxl15M7oMqesL9MjFUkfWIBDizHa5ZBpGGTZov4wMQxv8/R0jAe
Jie6g+MnPLijVfyBLMUiLi3YpH4KaR93oe+Oz13ACadjrJPa7idoFAaDYkEldpoX5R/pQ/OCg2Z5
NBoWHcQzd2XwhjfkRxJ7eT8Aj9IYVmUullKgRQy5eSgqRWsxtl05UifChateDRInFUxCyT/n23N+
cr6osQbTwcp1L8kE/m6/8mTHaiC0gXkd//3lV2vRQorEJpKOmnF/OPL4ypHMCvRQgAK7EKP01w6i
2iqh4lTUM+OzznuecNE81LhOGNoUFGrrRZckDya34yToUEK8fvml3rJtyzNvdUyODO2eYhGy/QRv
iNUr3s63DyMHJdQIcjFhzgYDUpWpC3Do0Uo2mH42DpPsQEWeq9g60r4yNMazYTJvr71D4LiqWtQm
BbviFA/o3XlwzA+RMvKOkZrJiC/1F2W/J2gRLjX0iw0cAOypWiCZeId2451n4TYzLRhvE+fMRAM8
qN88T7DwsTW232iOTaVTv9Fk7MMu1YRZtTZRszHIqKeKLhRYVDCDmVLvJ+FpfNY5gjvvMhH0UhmR
+o4uBRNORrsXuLkiWwltRL4/08OuRP6S++79yJ29ehMfPHdwPOVaVsdVlP8aRD5wfQV9RKDZyxRR
MN3ePiLQpUxCwU5GcGBIsJjWCuosNbfp+7arszT8ZZSBP+ru/27SiKv4sootdJKfT9WovZwgfXff
rzy+4VVa+ZEBG/aCK35inHPboQS/zO9XlXzkh8vCClNkUWPEYfaufb9kc3PHomZtmkY716KkX6m5
Hohe6hb8stfojqBeOE/Fp67DOXxNFhj44iwiSPK2Irl2xKElZow/Bkg9LGvDuDszeN6+nE4EuxjM
7gKLdoV+xtAyI2jdVtkgET6X+LX50/r+TFBB588QW+xT2E9JuCD/7SL2LcShx+93cOwS3rxMS6UZ
+ZkREfmswaHN7EeD34Nm6BGQncV6cJ31Hk12zlI71LVdB1nklbtZR6aRU8SW3xc7wE9b0mIatwwL
oA854WMx+Czn0o1KMu+S9zqf1/pr/IpyF+u96+cBwh55tNArDhP1gzdULY8H2UFYYOHwlT5pxXcE
NflFLgpkd3YBcjKFHpyxijF7YFTKJgsDHg6z/SAhu1820kmlCNb/x+0KAnecItFKTHEPyhS4miQj
SI28fpeI+D2fZUd3XeyTNv+uS/45HCAuYrtRKRxkVWMUu4CTvYkEdFL0foIYfhuMubInNsJencqc
nBp6dVS0k7Uu9Wn2lI/g2saRheO1WCr/8wWPDUiQihezcNzVn45+pldtzozt9swm2B71MjJfgQDN
kuzMnRXPBjattkS+ipehDvl6LOReL0yye+67qIknJoy8oQaxfZiQYaBJEzT0Uzp5wv2VMTT2Q/kJ
nV3Haqe9cP/hLTIS30aRXU67KiStTul6luGdzhUDmu9/i6hogPrHkr68i5vXAqhhel1M9UAfhV/p
WLr4EAWYjYwDjCja7kWLnKZnIYfGABw3dTgJq6YypYvU/ofk80dGAmV1FbLaor/gp9kQyezwC7Yh
rXgHG6QqEk9NPfx1T7eiMHVPFb2y0QcZrU3D2wxFZd9CdtZp1mhf4hbpoofsuHNmC7GGFSFkCwQN
VSkK5BXSeYS2ipndPoacVkdNgLfdMX2cWccZFd6tL+9VLJOotlyRK4Xc/PIjarnD30LbmxGa4qBf
dzJ//fMvFKRtqPhWZO9m7qvFDLqbgayw3qQoDD8jUHpge0+RbFvSnIlZ5UoO8v0XyPaqK7vaqJkB
WtquQeyiQgRMaAg9dDFg8R6Z+bEeXOYLTvYIhi5ajJsdT28yMibve8gPXXDCJ0RkVatieMVtV0Sa
MZfiScPW8tyPEI3KYU3wNZrbMzNMise9GoTd/xYtX4bn5Mfj+9gU6A90RXTQ9EBSBToZEigFq1Jv
trCx2ONopS+dyC+WNIhQ/EsC29u8UFGQqJPRS1rZS2d5+9W97mNuV0wZWep3SUL7oW4gkj0jFuoQ
7nlz6Qc9Lx7P2BLihI/B20f0x3INRpewz2bcunW2q/nJJKM9d6WFovpoM4YTmP9+20j4TjaLJWr1
UEEOy6MOv+9WzJ1uV66Xq9zRNr5L/tgps7JAANyy+mLczd3YWJBIOcxKW2Kw5jWneVWv7t/8bgeh
UumGC6an4ncmg3BUQkEzv7wESb4lURQ8tgFAae1wCwU2ZQcHX+sp0YQhRtzgxwcPN49E8WkjVqsH
YCLyNoD1b1iK8JXoGJdwzHLS8B9IzxNjkOr/BSsBSMCZRBQyyKT65KKNB7n/yUMBo6CW7zBhzMLq
7HLD9//Ne3lbpuLdZQSIPwIvkE+e5Ve5xf1I8fEj4Jl65iIqu4oNv1qTriCqmCZOZMBuUs+OIlpJ
5UPPvd8MARaa2oMBhC4fNGuFGqjHMTT9lUCmBF/6anLoRFb3AEj0BzOGs7WtS1plaifK5mr6o6CS
vq6HZZKI31/fsV+izoPVZTUJx9zexJINTTyCsffj8r4E/KDBb9DqyiKYGihvKaBxQYaNgO383wM/
xnL2G+wkkeg93dEq0wt6cifgB//sinXbDyTYIdC/GMz0rTUwDE6Ihpq1Wx3Jr2Pv/reLD/K0iTUn
uw9vv01gcxiakjYPasXyS3g5AFxTRKU1otwajPjxAQfXB1yYY41QT6me3zk9rguYfxTNMLSB6UOo
1kgt+BV4Q40YUGPeJszydMwI70SbPWlOSl11TDLpYSaYX8YQbpzMpFD8p3LZF8XewzRN5Vv2tSvM
TBJmRZwaexkUfOX1fiAubEkXdHmU93Ev5h13lqi8ua1CtRwB50eyxBcAxQw/ZhIqtJ+bZO7JM8xT
6SkRZ9uStAjbxVUzjRZj1SI0GMJa0O4aUO+oJXxjcRhIz5VvY/QJGHDyjAAiyV3lqd+n5Ko0KnBn
oYBN+BOnEt1PXczvhI50gcq2lK/JpKeUTA8O/Auvi/4u90hKye8pyseUxGuyzSh/iYxAmwapQ0gh
PkDXwi6t+EnBgx+oGwWQoTea9c70SWr5bRe9R0Qes0XAox9jSzCmMazMcRJaCbfRDjxTP0okhlvE
maRTcGFir9gWhq17L1BTjTSbQSdDs53A1BHcP95UaEwbgUejLVTv+kw4emCyzfWpVqEvw4amF6YX
bRr5oYRIxPxb9+WkLyd6NQxjmP4rc8mQdiSQKCeUP4dIyfMOczxZyzn52Pw2j/SDGzCO8TGHMGwU
aUqV77So+i4D2id2QLiSNKU18wle5Atz+atxr4q4jjHGsNNR+GRi3vHNSZ/rdXNevkx1HDlGo4u2
9qtmBU3roJk3aWeGBrpKATWmcz1Y1U1dMJv5Tmnzc8dVjt9x6RyAzTW7I0kSM3qa0THCnf0At+Z3
Ec0y/nPX9J61k9C7PSIqGgiljWLilF7eq/qh9aI1auDwGLfory9hjWvc4r34pbypDfQ9xexR23ow
eag2wdfp853epm4AltwRur6ArlLmP4ncdrcvyQvO5A1EPCCqBkzh6MIlLC38zbUpdjG9d42c65MF
CFUB0nHh+UuYe0WMCzdSEfBM/LBg6UOf1oxMABLh7UYQE0KL4dliQCnqjwSolK29TI3l4pmEKsRL
nrYtYx19bKKRkFyjVieBXxAVetzw4vjE274sz9GvJVDy/EyjQOSSqGLRsnBwnkqnfR/ffQFLwPic
2KyFtNgdWJ2Fr6SHalIkQXOM8tU2yepYOr6omOuxyAHeJ11QkbD+qobCY3keuKOe9tpAGR+qaAxS
TzJML17ZkXzqXf1yaIZIK/NsCTAtThT5KikNfBdGaRrGc8augxM4JcXOSCS1MfwEeoLt/+5UNF8Y
NIOnXBicuzCWMeV07kb0ykKyJf6RvRGp5SoyODbD/2TFDcaYU29bsH3Teu0rNEmOvvm7QTvilekN
c6O4JFZlttxpittrBEhuOYKR5PXdy9faErYShQtuQCk3537pvGg1MbTmLs7BvaWN8Yf/Yr9HVeAN
Axl/cXEmA/wvlWFhpoOaLzfl5vmmtF7i7RffWEHZXQv6nagphA0RrReGsLP0ZYOFpa2S4Iz4LtnD
ENNPDskiu5fCSoe+4jEtaJbc7CvbqIFY+x4e3+1/fMBNf4TlAW4HsH2KWRJheBvEQVT89qOzcDf0
Im6+iX8qLAajRh5I5kfYaOAgINhTNE4as1wm8WXFgiozo1z1dTsrji7Dt8A4QKlusm5LRoqy9Gal
hnVYeoCn3+i3px0DA85qbsjo8oyEbZYcbhdX3K92pPxTdOyYeV7mE9rHRBAqoPol3JxOOWYOKw7B
Qfa6fke2ZxkR0GPFwYV+DKA6DFNpJ9gURQfawsCFB2HtRVIHX0WygTiMwSQT6DJiA3Y6BsnlZne4
8++M1kOCE+FP7fsxENIPT0U3xxAyo+PQZATlWxvXwgERouZVDpwhyuVSdmnbJ2QTfTg1pI8m9YU/
NkfDpuLzDz+MP3/vBwmLfbHZOn9qRN16nnkhRXl+Zt1BSm2PQCQXQDBI08l/9eOPafP1Wc5JgJcD
b4uOAxNaLmH5P0ClyaCa8jZsnLCC18PZHVhipgzOy+uDLUh+tLBrY6ASonAE/Til8QD0TKYd4JnV
zCGW/iz21xFkFj5BymAxcxt1XX53TT7PAY9j8+QTUsMEZdUVMOgNXRLSMWoIEJK7oYmqZpBmD5YQ
+IuHDLB8UO4UCHs0wzD90veCwTr+bThiZ6pT2PagpNBH0Jj2t86rUtYKcfR7I9I+UbC979CYeZTE
u7cd6ZJu8Y7dv0te64yZQjvt9e/bKTVKxQUqcUknNemD4v6qeBRwVnA8l6yezM8cKfRaCaTRurHV
1nhGsJttfDSd5D5F/9sGlpNRjn4wgs1+3jEsqPMWoMmyjv2IAmL9oNbzkNNlOZfn5rOcRialg8yO
FQSL+jN3Yu4ZuL4MQqgwdc1aTpjyJYQk8rFhcn119tcaLk+E4SU8LlkkjkLkDfhTUZbRSx92E7RG
h7pMp14BryKyZ5o/VwqAd3tCVWuDvrBjnrqKCzuK5KHDpAP1iF9vFYbE+We4SoGxAnONKAg7q/ga
4ZtPfUJkzmyfgDZrriGnnwhmaPQwMWSDlShzSBipNEgGOIBcDGijkEIvtCMQlOQcudZs2esQKAt9
Lhck9ewb5KsoHorrYqhta8v+d58ClhcTrM0Mki309cvhCUarGXPpJWanDODG8PkzPMzw+HQfXCG8
e2PzJKCgyhOJOURUdrnPxZAmHJ7IzBMqoptLY2sJdFF9n1L5Dt8WbXLyfKNscmoh1WbsTnS/RN7T
YuI9bg9N4aYbDZq61wCtoRZ2L9QRg+yJ332TIJPOi5+5XEHG+aYBzaJpfBBdNFKf5J3vSudqzBct
0ygaBHSazLkOxMlXygCKjKsGekX2ogh+plh3XrzLTW4dVdFnQ6XLCWnCopdDe9iLHukIhU2D9iI9
8xdpjjseVOvQ2u56Fw6VoRgRmqnif8b5mYCCqDVC3rbVkGuLyuaVw2BfJAQRHGIcxYQIA3A3RjJe
q44qPnAuPo4LbHf0eV/JcVfFKR2jq41ONjlTtGqjeZgpCB+CLoMztsQGDQagaqZ810ACtP8vFjmv
kXLYqV4UOGxhxmzHUCX+lzBnwJZ8Jzv4AJLTZt35Jpj0iIYBVRJIF6i4bbBTpt0MjEHBzen9bJUb
CHu+um1CoGLNyUkPxmS+VLJVGzSalCjQvTqKxAOMHVbWFMXyXN4aVSYVToBjAki/sSjzQz3WnmTo
N1Fy5AoS63/uQBJVvRY7bGDT4eVZn4MLBZnREn7WSCWBSt9a3KUaVMcRgAm5UPcvh+rrOULzrR02
ssWHizoxQDaLpThJzyk4AEnLr84RcP6tX7oSIjKeNvMgbr/X5Eer8i5b2P9LURNkhtGjzoUCwRK6
dhPtFBatE1Wj0MSlMyk0BOOf/b3a9AtnA81ffBz5kJclHQO/zB1jnsd48rqmO7qNMr3qbJT0Qj+u
8SD6QqT9NEV38mUA5soagHIwCujBvdcNUN8RpetZdxXRDTfuUDceYqV4bQP75bpwz2VK7cwkw8iA
G9+cVfODkoFamZGP1DSBYuWu0OEAAUwv+DRKQ629POtowbJZEMJc77hzLlv/k2Lt2wETDWW5P6yB
rWhsvP+ljGI8kk0TyOoAZ3kLFOJdWaRNkO2yAGaW4u0AkSo8vSk5Cd6+b/AdPmrpiibHqSe06CkT
g9hV1/fvkRvbPYQvK1zr3CWVAeAyvyLcq1lzW27r8WHoEI5VYKpa395oahpkyJmK3q6g8AGopzNF
e+Ccqu4iz+d0YR4ehEanQRt63Y5uVfsasclNj4cGVV9sdp/PGZQGQH/OmIqWxhXubCLPKiHOl5Je
ctV3iGPDye7vE4sEKmHmWj0jOxa0GGjEc5JeepSG47aj+Y7ah2ADVOerZn8ehGcoaDSL1CGMc0ES
SpKWElS3NV3d2aBK4UIzuUNYe6tVPNBAZn8AVP+QCW9BrRT4pw8y+QlOcDv3gVFmpVp5rrp095bo
JfUcte5b84tsNsVDHJpofum0kJlMvSQIar5yLTzxPo1FCoa2rWsUXvdQ2GMuwE98vvPfKjLOL64r
e06xryjfMixzPEGSFtXyYZfIh6eo8eDSTVe/rh1WesVAvd4BPWjCXNT0sCLAzJM1Vu4V0EoFiDf8
Mza0iGJVhRdguzh51k8cpUvpVKwDmx35p7+vWZX8vrLvRvF2TReKtUVHlqj3GScM0EEq8BWTHk6T
UbZ++HbPuLgHXkCmS99yg2q9Ua7aak/N9/Uu92bnxeyAUbO3IupbupqsV4KEw584+DDxZGlCoXhL
2JLRybPrfYG6xY1B8CKdNhxoyRtXje6iJV1KGRu27Qj4hUxqI1xjZ+vI5btwnxQTDt7htaYtb1X6
xuLvLIkCplCKn4eEZkwXbHQ46ZhArRUFapHyx2LSYEMYKw/qTC6XTirsv4jSMTKkFUUKcCBI4K58
cQ15DXC3uXB6LyFetx2G/tVpuUA6+v7X9iz0+agRtj7JUJiywFbTTGsrSeFsNiqo54IRyMif/j6+
P9dqu2M4B0yWTPxSkWH3pYbPMK9Z1xtT3vZUkgW67KKe5bp9KrUgeNSn7ZNCYHP/U9E070BKsSX7
TqULJQ0dWzwAi3WgAiiCvLHRUwIP3/04vDYuupEmRX79VX15QjgYe36FBtAUTIHBWVpd+fS6n47B
w+bcl6yUtpuzkNfzsTS7UiCjd7eoaxQZmrJKdzVQ7v84yNl9Zj9z1yHS6Kkxq0Bc/2pw/ZdT3xU1
8s45gumkSshWcGxo4xnptxImx6wB7Vp8LC8uqnNKOXQUeBvNb4tnVy3NilTsB38Dh8L80+VBj6oS
YcpC2yjjaXHMbjIHL1UUYsye4Iht33HyG0QS0j1nKhSXYl71Jxg8rWiNHDa3fpjnLjOKV83b7tND
/bZTTryVWiKdH5Bio/e9S4dXvgFAf8UCIHle6efFQ/roew4KMrDeoU9FaFRPg1K+sdjB6NtePWkU
jj7FQXPLrz7vq9tcEXS8VoqDPnCShfRW/oBs+Cn7o4AjMeShcDaFAoP3hElaCA5fXdJG/khC7tFQ
816+5xB3DUuQN/fwNGWoWzJn9V5hSefrJ3dOwS57ayoE7fG4470lg8UX2h/wbtAGzqTC+b9COmpy
YT8VXiCofHCs7SW1gMaofm8CmSyzt3YkLcNkuVwXluFqnCUSgWaBqEWhc9dKLCuZYnkhgZuMaVgr
O2xUagaIiq39R7WPdwMQZjI23iqfImZYnTJkMbK9amV5LCltObiktmI1Jp09wk0HM2R6BNdXqWG8
KGBHHxZER5AdhS771QsfhbDtrxubv4jW1WX+IwH84WO4k96j1+GvfK+T2Gi2lQEl518/cZV9IZWl
2W3e4/qfOOvy/HDYDPEMTeMScSAKRi2XbZqehilka6ftfoXsbyJt43HhEJrVGs4Hhife3ltwdvmR
0rBgzOuP4JN3y4k7o6DLiPaM6RWxiJPLbvbyBIGkbtjLLGR7VdNqIig7XvvsV4kNjQjBWEdbOJA2
upKxCjAA+JKrQh1hEugsx+7C/9xq5xYprn5ZG+0yJw2ryLOWHYyqdHqPpkUSYAqu8OUFUb05Mda0
Vsyy/IyMzxkGb7G0gN3bs3RnGJvEoGiojqQEUxxhK/ymkE7jTGTct4p8Jgr9olQNdOslLfkTmB8V
E1TfoRSovSb56HR6nT/KUnS129IFoH6QkHb5wNDBBmuzqtOWued4f0gJsTvozvl+JCcGZWgkUneO
bBOzXhxdch+JXxkrEmus/uceUzksvbCvpNUiGxYtYbJMIF+Ym/0yfaIgXZujkJ5B/aZf1g4Tt9DM
roAeRW8TFy/O75LIjZg7v0GsDspegq5tmEVZJd2zv/B6BMnR+lB6ZFhOahyb21AFjIAwDwz55D+R
eUMGyGSANvMazwdtWSR/4/5yikF2X26o5uSKO/2dvVa+jIdXsqetGh7kG0fOL2BNwzt4mn1MOc7V
bK0vZg2EKbNQALomXF3qlYY9/bj7zio74Ns6vFGPRfE/p/x3Nh5JUKPqWDHPJ+JeG3rCcuqKywmC
rul865bVxVVlDknkWGtCKbAFt60AXC5OoayXBsUh+9zfcExDesVpI2Jryh8mNjIB1oLLO01YHuH4
Vo5xQzsuf+Kf8hu9uFfspf85QG1sqBdaWUtYfRggrqKwHqHRz33U/EoxkMqL4A4fuoncIARDboWy
uSIKYSKb1AgSOyICBiKFG5vrqn+Caie8pvBrhkz3G9fsdFoJXqmmIJ7IV6QQue5gtWkrCBkaAQ1e
/xvDyMg0AqLhdmODAH/3E2T4AVbdUqSW4LGsOrDxC4bQICeKkY+3M+lPF5wKZplefLjVNpX8LDgb
+AuT5CVu9E3XDmbkzP77t+g7LlfsRUQWNQl5SA1EnFOECQdFjd4YzvKH8qw439h0moXZLiduZPuq
ZFsIBo1/et+wU9moeUenl5DDkmaNWkSGmaWldLNXsF1o8qNSQldq2+ukxUaoOjlSJrSxEvls/tkW
QZWtHNQKdzrLqvmLRPAK/nfc8EZR/oGP7kuNz7JuYmQwTG9bqChAaSslme1D5vYvUTg0Cu9C8/Mp
02plTzZOSA0GO45kWltWiqrojJCxFb2gIS7FxATb7y28XbMIVwhdsQP/elvqUVNk8fH5zLuFo1Tx
0ZJSADauyhRZweiBgDOl1S2idvCJgSc+4qR2/a3+rioTszVqaPna7vygnFMd02Lt9MXqFjF290l1
XoAIwl8zDFwx6rvbSQSuC4DIRjh7rUmZj613zc5pZNQAsFbS8eOxQvlYU+NfjzbD4mfdVhGPi6Ld
hHd9DmU8bdr80ngy4/Cr90o3ZsA4qLblVSv/0hRKLE9XD98iSEQ22BEg+RWX/cTmppuWFrA5+Wds
7UdBrwOQyyxFNmzOMEncwdRNFGyW4niylh4wBOt2nKNm/8R4bk3Jky9YHCQs/pwI+wlJSBok7jpV
VQq4rI/bvA/AKz6jnZxDF3ZW9K+wVvPOZ7/q7sYKcpV/5LXRtduSLuIK8zsUOJyaH9eKcDjTa2+i
GowpvJ5ggQMdC7BirIYsH4qASFJi23WRU6Iz94utMpJWLbDHnpS03Nmd6zinSwIxWYLbpS44soIb
2kmzp2ycbjYiKe/6qdQ+qAG+PQo8WzKWhp8TjWq7p05l65kKuNEHqG7Avo4h8kh9DUI3rqcr7WG8
V3OBbQ6y59LqRQHzFcsQK3DpFYQs0Un6DW8RUBOUZlqTemuu+sNy1pHrEIpXst805A2VqbeIaHie
6B6HlqvZ9OYSrqH3bY+VckyYH0FQhbFYErflRLhcRB0G1baR1ppXTb2tsHQ+ptUargOy7VuJfTS0
lzaEDEJ38Iyqo2DqytIDT/WLJ3YqfvpyE2SNEAN+r3gh3XfGXKnv+Zy6m9n4WfHGCHJZ5V0yCI++
5MezK+2d6sE9ETy0Vj7Cf0oYT1NQP/3E2f/p4vinda7+g/o69XcjRB24u4j2mexu91/Wb0zgHjy8
iGVEvu19NAfewfaIKHgdYBO0j29bd0QOFzG/ytGTQytRgl/wnr19OjxC8YdvcVpRMmIZT75Rsknz
U8Cb5AlQjoW3FgXKk5Yyt0tf+HTHT3P7G57zMbTuYRhwAWKBAcfv6pDrtHOr4ydoNFhSv7TSHrA4
bwlg/a2Y23ymm+x68gIFRpljfw50BDCdt07Vh6umhemCfFDaTBgsH7Z6T70Uk+PMUpvwxRLY1BOB
Ecs7x4vb2c+GZuSQOKeXIfCifnEqWKypFXSJLdthou+dm6rJaRElfPNqTigwuJDX9n/pHzOBd4B7
jfZzALFMaF88WECCy0LAaK9oUHvuGv82CoeM/ABWAoZYupqnsV10wzckI5PLYbsRml2+qz4ZV40c
YevGPcGQzN67uo97sscRv90qS1fuzP6riJ1vWejZD8JSF/3vvfMGmTK9yecAkgU8MyY1z0OqDGH9
ZKAPiCHz1fs8WBBFEWAVSQbMDed2FNDJwKTswppW8T1Sh6dhkzTFGJT33zoWQWxvuaxloZ4/K6bj
KxgCBScnH9PznM/Ns42plKGQph/RVqu0txZ+jIdAbh9THaNdrOa5XYmRdMHLb1Psw8LTRkGt5I5w
SyG+fPCE3CNxkzuzFuC/g3QDNDT1TuZ1JGSiui0v9qmNTppsj2ibU7Y3ThJl8BYvqOh1zqYW6bCO
LnaNHeELKKYb2lF/5AYVD8rKKkwLs+jWS0avTDAQrC0KiYIfLmx4b+8UvHx2px5QMm2X0CQ+QDXc
fwyYWWJMIaDrrRrjr0DxsO/IjNvE5DV3Rf3eHNfWG8GncDOBzb6cZnPPMxq5dNFbVwUD6VaqzSfX
eW7ihDU/sqw5ELnWR8xClKIQ0wGwVsuSGOiZvUFt6iX8WemHjhUL1+1e0LX4tzflv9LB7y9/eZNN
TdlANYTh4twQFdZ4u29o/CXCpivzb2U0d6iFVM18gRUMkT5cU3K73aricp56KjdH0RQbcxPB7dPl
WFcNHp97nscvhNYEe1iOvJHm3fUhbkM8iqOfoMi7To+4fxfcRGehsNc5ToSarZjIVMpmxQyDQCbh
zEQ3SEW0Ol/0AFakX5Wn/DteDBSjH4qj4l3RQElct35iMJg0VawDqwqok+s7p/H39GoxBtCq3Gk8
4Jn7ZZY2qJEfleon7eKWTWpInkCIeMf+AKawrOP5SaAyN5N9hpbBeimSluIppcYjVSAHrNLJ/r8/
IOiyxcQXtzLSMC+3erPsINKvrJJwlQKJ4YP0D30/5hJcHHPltGrGTU+qF9JH/XptPRV6q5yJKQGy
rb87O0ik9cjIXu1/12CtCSdZhiHi28X2mo8PbihIMobiPLSdoega2usFrVjjDm5g4FJWhXsrDC8e
pR6rT6TmCrdzFN+ABPl8x/dcFBWxtVKwI92yOgVBhk2mJujP7mQYCbmYadxWLLesIjMGcaIgSYzD
ggdMywgoXXNhe6iv64RzN2Jg18smLt2sH0AcmH6dczX9Xj729LXh2CZ6+4g+DjE8qDa8ldLwF/Y4
C88GtG8QPrr4p/COG+U6IlEpus4A7OJqMizdT8lRpXf7uVFsmUBhaLZeNfQhCyFvs5aepTt2G/n8
Lm5mYpef9bY+4HJzSmw0N5DqkcmSPVoFVMUycAH0RvQbhuYeGHo3avWl/9mowIN0jegzY80xIPUO
j/tcbMGMpiC/kfwTUGz1kKn/vXWg9Ky/EwoLBDHt2vXk3GDeU7GgJt1nCra3xLPGN7tvM+yoaHtA
ooptUVGXxlxiJa0fCKhUTAkcsLzQUZL3gB+5RZkekGnkCHYZPpaqY1BdONyM3BB5lSytPZZQd06R
rOpLAzC3lfPfd1UsQQSWrFvIEeigEq1Ly/SsrJsBemqI4fGu8WWEXhiaiYME0PgwF07Dj9c5UFZs
loz8eKZtRxzqyxpY6K09Kwnon2S1BVD7cDJqiDKczSB5goTztlnHZ6KFi+v00rF3KEDQaDkNVgc2
U5iGbDQQeyC9xTO/8OSfjENfZN2pR8iKE1iStSUlYZNQGPchafnIuvxSc29erqON4XA3zocoX8HL
bM1j26bXQLBr1U/d9PjK/ouabgGLH9xaKAW4ouXJrndZKtwTnvPFqXM/N3XE/MHeOhPlkJUfOdgX
UdXfONqjmg8N+lI3lc02oCgMnNCZ9DLbFIJ8PqUhy0qGHet8XtC0ztwT0Zty3/mO5lz3HDkjaPg3
Fv1dU5tIP+FvlD1gW2NQm4AW29FHCfuilAPudEnj/JW6K/aBZpgZRpLn2Qgm1r+HS14cIV0MejKo
5fROpo753QdD59STsMVxzPvzl/Ipu/12sqoCWMYGm1VCvnG4qD4KIQkeBPQdaezgfDeczJDnzKiD
DiDKlq8WBI2gCMrB99Cg6X9z55x7eAGus2F0JgIhWhTD3rDL5I1LoH/9Wp0uu7Bmb/b07XJdrNaT
NyBjqH/Iq7OF7VS/3wylCiKTYB4jjSDOUnUcGP3oQIp3CrJQiLtEOJRY1eo7ayEnc65v3iyGcLxK
G5eGxdcMpwjMohmFV5gXOr9isoh97DyJMDLM7kreUTcPCJeWi62mTNyfpyPNbwbk8Ka6JYBY88zA
6tcwZf5Mm3BXcsV+QTNElPHTwnBjmsDLH4eox1mGcFMlX5Qf1oYdrQZdlL1cAu0LR0fipGUAYvGh
DyNoi9JuO7o+IDfBujCNLQ22dGsnFcd4YdQJyPCqBO/7GV1QAJL9xJp6aCB5ukAKWxTgRk946oC9
9nXQoKt9BC2/AYUeIkqt/ZRJ02BZNyQfz5Nk/1XeG95AkLMQTYpVgpVF8Bbm6IWgIZ4+6IGKnE94
+2CPlz56eV6g71r7AW1NVQD/wOIGrf3eYbhfjnagX886dQysHNcsjBqrTu+tqLX/9Relu2kalbdC
h4c9Na0kjKsJor99YwdF7eMgeGofgg+bIjimheyztQL+OVz4t+YYLj78rvT6MZd3JJBEJfF8HUas
sqz4yps/U6d+cPCFRjdgAsI0lodVBB/AR3QRsBv3nB+tBppt0VXqAGaeZsewTcjK0m8/AIRp6pSb
tWgC2+N12zse+qh9mRzOjjMgkSGy7UqwPwl15F037oPwWj9gsRwdGlNwQOa6sJwtdQDcuNl+9Bpr
IuaO6KRkPQVFe+eAIIimbhBgN1xeoUWUqmeH/D8Kj8/JUpApzAxIZ4c6XlhRyjZfRH4u8fstw5zP
OKaxarGDfSNMPIOtayMXDU6zcusYCNqkd5LRPKL2f6s7iGNU47ggM5wrXhaxNhICH4RiweXIZ01n
r4YnVTclQsX1S1lnS4zA+UN97QnJDKVt8zQ5CkLb7ibkz+RygmdF6noAz58ZVaLQV7V9m0u5zc9y
lSOd8zSN2hQ2nOIq96rorIs/NmbCgVMFl4sQIN4jSSrmvfwFrtrzzYv4/j54ERDLGQzsVYOIcca0
RI3OLaaMkLyS/FGoXhjucWpjuERcPdcY7sYv8XoBIyc5rXzYJy5ytsFvp/50hNFiHtBfxYWK8lUh
Q9hLn+ww7V/7SzUC7VVOp/70RkQM8+lqtn3BwsN2OCrFvL0WqUsZ2WUJAkCoPCFIJDoKJaJXWD22
GkGM+MEG4mj6Jx3yEj36LNBkTLfP9W2aAvvwwaKldlvzeX5BFyAy9IqK7qcRGeMMZvGbMsn+SPIy
+5T2bK9jZdu91SaE/DlpY1I9V0+S3ZmjpaiiY0ywNlrYxrSIfhfRsGTikWfHPobjKYbT9wgNVeNZ
4nd3HYOU5G1qE1W7cCXgu5p+HPz0QU4Os78pJw9ye16/SFKYxmwKbnnSRdW5DL6FZ/M74ArJy/Xn
jGO/XLcj2GIwH1NwmX9Fp6XWjgmyPUVCVOeDt6ko+81HQGsbZXnMKSY+CGjGOWZvuy0q2N0ng/gj
pJqcAGDlZBopqxMcoXx2nt7Cjl3wKsRfUGLYZL0UF05s2pKPv+IbKoJdYvmJ1YQuQMWTuBBicSLd
o1rvE5BHzIhaHXSVKyroJTdKXpQiw8pcaSnwCw+XX7o/7I5TyCTafkUyjwkHjDGRUsvd5W1Xs7v7
nP906WAQbce41O2rSnnhC8U9YKIGJFUCac5jnTId7oLTewe9TfJkkjGEsor4WIJrIZ/A7R+4UX3F
JAZO/9As7wx+eI2ZGq79Itk8KI2lEr8k4c5B8R/AfIqEAaRZ8f1s4JcJ0bkIXhMAk+fawx5mT6se
mZuZXfIWqaf7O5nbF6+ilEjhooRXuZqysyDVTWAQY0RQwaY5nvPvkfylt77/dvkGBtnb18bapYWG
y6fBYOhgyG5Rs03Jkcx7Q46fXyopnxkrui0vGWyLjLfXrcOIYthsIH+xzgy2kCrhpsqqp4xp+WP2
iZpkrpn5KGcShiOCCheo8uRJri5wkEhXoSBFsyGiLaOeumLxzWEtQWLzJn5P06YG4/4Vx6uTER/F
TK/qBPoPSY/lNFamQHl83ZRIeikDg7uZSxai+q/P2qTBKQF96HtSLbuCFClKgpMs6M9TG5NZB3ar
rqZOPi6nwNXvbDkqTmUGasLiyxP8hOxl6YmBnL+QJJgpKJ4WoWUVQH9T+B0Wq1eMGDzkAsrj92RP
o1OCnzggx9t9xPF/J/+i9PLvvHXgoVldS8eXx1HwxftnNOgBRgUZz9I7FknifPQjHnye3MAfBpAB
WEzZVpTdtMJVt4OyQ1AuiyRMKUly+RQXh+vHAcGDJIy3CW8NPz5e3rIRhNbIbQ9Ojf8ITjyO/kh8
Wp5fio7thNpcuWVyTUOlmER/nQV8WxEEzuDUcMDiJwlUnjiZHO9XBezNpSEJr07uMkoIkLV4HA8k
/UIzp1kjsbG3wYSp5L5OaPTq9x+X7/mZw3mkD3mxajCMY7vjuHzL/1u1INhJp+iTRUNCOKJrIrry
fncvoKUAxMjDbc68mfmtlGeIMIjn0MElKvv3psMvI26t5NtBWUJjf22Ya4MePbAhkHFZBb1/Z0FT
VdtV63l6TI9y4wRiR/eIHTmDrCv1IZ8NbSzSF6CZn5YTqpVmIF046dTap4fOAs1ybUYI3JriQiof
vnfOWfRH578eP2SsBPrNhu2euMAmA8AW1fi6FJyMitvTXRqefIPOEH0wID4rkYEyGcMk3PXiPblz
UJSnFu0/65b+Z8Z8Ea2qJbSbzbvdhGwLwA632I15Psd11m5XOnh3QvGMmDwnBYgqzR6vU8470xnT
QHTmfQoV3nOu6565hIMIgp0z8X6OBGn6BCrHPRUtd9AdoXZpANwz6Fp/q4Mg2ZbB+VXsUErUJPvs
nq9MDu1c5jmCEPdnsAn/w4bkQT1ukX01UfjqJXNKoMw7FazDN5485e2tzBaWSYnayxlzkOM0t67v
ZDCwhAWmC19l4TSkjbwLiNIpetYfsvY/dHkAYshkhpBd6QZNO8opD/LXdCjeVsGOp8mCumhVe65m
/h1kq+HcI0/KXXpsPnrOo49YehLWQw/HNUwOM/g8FqfS2fSZsE1stqHuIaFGEUOuuVIyp1jeM/KN
+tLdsMxVGRtycEK1Teiqe+0fSzoaGkHTjFAOjpF1cvEN6ChfCIR99GknNBzmgBLMd1laZchJ6p/z
dbVtSfANz1656XzCTOtiwvYwmQkWJ0kzyi3CHZM8KolliYiC7uxxHCURvEhm8D7Txt+dPQ+RN0L3
nY8aovjTPjNkEL2L0gwG8CfIl1Bg9GKAwgyy//oo5KWa6oc6gDiGwOh06Ge+8PwlwikcjeTas6kD
q2nwA957cBkpkfP9b8hq/MyoUWMWwttNZ4c/+mqOkv3hEP179tv8gvHpRgpUesTcIBadRKQbGB7u
xFqiBpeMYp6GzT1RiMJW2/41yCNRnp3YS5HKwaIpuU4caXPCjrRd3luW8IMewkjDSVBphvfoK4eJ
2Z2cu9mssPECDaW1piY+oTUEXkpXPJId5udJigyNeg1VwVoL2SzvFOUdOYiUA8HO+xUEVjlZpCQB
DNnaY1axifsKnG2C3fwe4rwNvQCb/7HTVuFcWK8eCSU62Mue7ZkqVYUEuJrCysaNq81yrJtUPij2
cD4EiEBKoiiUSco6kE4sQXrAfkgC+jTvSdHOrlkEmImbbzPGB4p+A/OXMaeVsWwc3RXzihpShvvA
mrOTYTOjKtcQA69L7QypbA1V7uR/2asVbLJDV2v0vK7HZgRx+HIH3G7mjtC3XZY61JdEa6+rTBKa
ufYgABJWGjqU/VK9DlUo+jK2Zv89nJy3jtBqJsn0FzEo3is7+QV4CJnco18VLkRER4HJ0GUQ0d56
rveh6dIbENn3kYiIZovy3F6C2v3+mzyhmdY29lW6QUd0UXCCZb1torqNPPHZGxMjZrk8GXG6RmWD
Q/23jbSMf3/B4TfIWq1w5IRA98UpxMeqNlNEcBGIMeV7rYust01lraUc6ZbEcKu9jZrA23UAWCyF
5TsCrzKmimdeixtM/9z7jg4m5Wx7o7ZYbSiTySN3bhGRDyXWy0QScqCtYQZYG9pvdLBHIWgZVfgP
SbZt1/DX36T7yJkcRS9KpSfxv2Vr/AFHmwJJgnYCqLVQBz31hubH0DiZ8ZdqKTgKsne8sK28sp7G
unm3SjtZyLEybwuqqShPQhktfih8Eg88F3ZkwHbgVth1VurbouH+7HQKzK19MInpY/1DSl1O+LrQ
dXnX+TqhQ66EYpqm4uiM/vbRfpPA+gbmmRqVtl4J6i0XaYpM+CdFFQGmQBBGUWVv+Imq2usjj5/l
2ScvLRvxH7GCQmMHDtngnMyKpKr5QHpV3lReE9x0BO2Q/Ccf2YgJ9KuQd/cI+j3HZ2MQ3YiRFt+4
J+D+Kmdavc4SOsz50tkuptiQ5MYBQBbnKfo7eqOK6kzFVrnYpBNcxjHye1YCYvrmBqTPY7WbHHAM
oMMdfF32cqrsF8sjCbrg0vo8RQYEAzVquNwhj2A+KVA4/5mWli/e1u/4aAaeHLOicHdgP2Vtu7Cy
s3bCy/x+dTEJCAXLvrPOFT0HnhNyOD6vbAeZzrFkiHkvJCsCaCo8eDezMYkWE51o2LgEpcVSB+qV
wO1D5CUvrd2+seDxcWSDeU6j+Ky7o//vqKMGzC5CdmSczZsNzR7Lod93vwwMwC2DrTubawlEeZy0
KFpiXRRhwC8Yc6G8coXQsWYsABnX+bSDW3zvqqHXeYlbGmdjKnsrfNJ6MJ+MG66s/ZRGYVubRsfq
2JhRoYBqUqYjr5GkI55L9sVnA0la1+jDoQG7kPbX2UhjLhHCcAtYwtvosQhEyVcXRIxG5mxfkkj1
HHtlJ7xcAlMWK6lAt3YBBuo7hX7XhDDHnFKtMLKwdvJi87NU9Wy8wKFsv94tr1MZCnjNKAEPBNVF
QL6Ae9kjy4v7og+54b1qs2hD2cw/bJXR2ZKSyTP8/hSO4ba5E7Dm8Mbl5HcQ63uawLv/ql9/f6xF
0kwUcHNgjaQ7e+XAvjreyJc7nBf/3TfSgYi7VKgN6YrRktaE3ndolw3QSMLtkvlHychuPqkfFae5
eySzigvOyIh6vN1HYA4+RPygGHl8NvjJC249EiAlfK/DhxKLYJb3bZuMtOaxp24P5r4onksc3urI
3aohxesveBRWR/jPJNgDjXUM0S7gissaXjRo8gtMDYS6EDGvfFYvuUrH1axfdiYCmqqNmQVIeHB4
gwt1fihXMJh1Piu6p1L+qYAolLqLsprgxsQpRznDOJIJlJ7amK0ULXGFjFzlDXZ8zjV7rbgbCqew
u96h2TkYz9Y+w6IyJTl7Y8SFgSwQ/ZeEv7h5RWJcvLPaJ2XRrr/mC0t3BtqOerkooY+5G3Z8umBf
SyL52R0WeJ3mm7iQG+hL+Wl207pfIVEClqp9jPBJaVeVP08WNqsaQWkDtWj/BSixxHdhPy7ZfbvC
mn/0axanRLffm1b1q0F/iz8RBA2N3qrUaBZ+iY38NxkLA5KZPM+GvPdlmMgDXTeo0kxlq0jDMnyc
U2s9SNWPH9uhyA1MXzkD3o/41ooHDG9GnIdzq9N5Yg6BRzPmmPC60B835ZQ6He1p/P/DzdOJqn9y
wuXYSY/0IxK+RDPZl2yIpQQ0Byqaa16LhCzrj8bHjhM5w24mi2u4gOehi3UoPWNwOfzNnn2UCJJ2
m3MeHnASCRnadt5oOfwTqYvjd0l+duqKm1JlZrysmHK5enoD2gaIfOMvbdqAlS7ZShDTEsEi4FSq
1bO1x7ojEN0QJNQMpAegv82b19Xd2adAuDk2qbpR3blbrujkkYbSYV91jYgyCjMVD0S97D9lJgPw
UDw0KUga+GFB0e0188+l+yozqaS1wULpgZlnppd1gcUaXna93JyPrFK3CoGQ9MppjRgS0RqTv302
WP0jG1zBQU1OCPuV7uEy3kZISdas4yxYboyOHSG5Dd0CpFUAFzozpuaDew9mep069PVqgpeNtxTf
GvtLxuz0qUCVFgaaHJ20QTQa47WFOx0yfHDJgBG8tgAqrf5HVULDlo95xCZpR1oqED98C+XablIk
RR3ht76PktncL/SFTay7xH4ElcDxU4lcjtI/iAzz224MvuU8NhD4i62ECgN4TA4SKxzE/7sItfqr
oBYHKJ6u1+u9YNF0oJ2si020izexe3jQtqbnhcKLQ3Lx/bwf5LjR2TjStQBQeHgqveYlW0VYamdB
+Gc7ZN57UH7XBW1RBIfznwfRcow7u0nIt/3DRdPO9SSolpG1mBk2jZ7Uv2Uvl8T8rMs2B3H8uilW
MyZ7JZ7zwPsnIm18fMfiavXC1oNdyvN2NpWARD1rDsjjQBZ0EPrC6W7h7KCd1Qy8VfRkcvkeSZr0
kNT9t2bNncOipEepLfPAm4i4mY1JhTQHCF65b9Qgyr6ypwFuXWp3YT0+giJl+8dnD7BiqZGA8R+Q
7OI5H4URwJQXmQsw95RI8mLraaKuHqR5GbFkr/Tr1n+kkfUiHUEaqlNU+7bvsxHKUYoIgrUb952U
eFvkPereFD+lPsM2RAs5EM3Nvgdlf5gSzW4DSb31OtWFHZHFAJY2u5LGhLqz0JnGj2+h76uJXkjk
N+zkZMEysO82SRPKSyny5nZpncRQdwUlsk0WfvosWvz6/+rwRA3Fk45N6DpTkvxCmK9/8Hrs0Aj5
KmWqu2lnOnxsBVwr60yANE4DJziDTw/4uS3f7ylABy2pr3FqXD4fspFVcRRNnjbopZoeX9X72v25
pj+ztmlo6tvTT9CNKD8R82FpUn6v3CabR+Hz5ZTzoW/9hhdi1I5BG+0Dxg+dQjPSFKSQIJv5wM6k
nZb9HxNq6qiVhxInTTTIuYHBwQRvKPDS/HjZwIvfdiOS/kD3/jlVlmp1Z+Rm9LUJS8a3R6D5Owlw
BcE/KOS/zaPGgPL0HNotsS1LNLhmIl+B54FUZdfZbC1O6UPwImGtqpOI6nt2DctComCLx5wBO//r
hyGCiiW7UVnAnw993BgSyGSmXKG99Urfw0SlEu0wnzFMPSAJoq17OlXbbCgn22Wx7W9uhdlOU19E
ajQNSixRWmb9SumyfvAMRxjf9uG4RlsCF/bXnt1jgYZkjpoLZKB/sccC1b4VTKixZYO7vhTtqTGk
XOxobAjoEF0UlpAoDUNBhbdyz6K98K6Ro3blzeSiOYTVR75ensiCcrOsjpi6CmTUSNj3kpr+70GA
F1aOVWinHQaKs+8RtvrZEgR3NhokYAXqwPtaN3kOvGqAPm9H0c/07taz0gE1bMGsx30yFI7oZ30w
zRmTYw80SxCPVxRXHWZsgh3Wg83N4/WQru2Qi4dSZQuc5p/SZ/jk+dq0y/t7vsZzyf/byVYwu0zs
tgdKK73YN7GcSDsIvcx5dB9eefM8cctGUiu5vaA2RdK2l+2Y1FruduCcP+lOwK8RgTREgaBiokGU
ADQN/BIroFz6I5v1uHCSsCIKRIh7ev63eLQjLd4cex32d/6NfLZvmJOJ+RjgoyBoNAGJY88rOyxs
ykJPZOFy0dZgrbORKcu9xe2pCMgnrDn+U7DSK868ttDk8A4lYsS4h1SQh5ayoBFX8Mn4L9QjCuHm
alvHvXuKgS7TgNT4ghBYTf0t015m5I8qbUjAxz770yRo32h7prAzJHTUJydNLxxunFYtDz4f9b59
8b23i8U8mSDMT97cAYcBANCW3OawV9PhBLj7qBxT0njqmfNQVehYc9J4ah5YytOAswNoEfRx1k5x
0C42G3ws+MGB/nTnvAkBnASvwZ3PANHNhHVbkzTCVrhu2KyvzIjsAb/tQGxtBcHOcJyA+qXp+w7q
GO37hVF31iDlIYqImq7mh045etMhbJuF6xEVNTFShymRnThwD1m7WaV5+6ey1GHdC76HnnSQ2EX0
/WiCt8hyr7l7SXvZfW61guZaoQbUVVrR9LkNHDhDMY5jyYjtMyu8OxrjG42qD+1ROox+NadZ19jn
yhvZTZnTrEuFPEkYZdACkX8dXLXCnMbGHVMEjxXuwIeasc/1/H83yQubOiocCJ6haiUpEwskJfbN
rhM+VHnwR5oQaXYjejV8pDpMtNBuuFAADEt/Ekd2cVhdwCE3rJfNLg9itrzJerVA8qQ8Rd0BqqdB
tADixS5Bpa8acP9NqxPnrA0STaLgXeVmXocEIIBXP5zscu4vBSS0+fQJQ6BBaiuDVPjbbVgB97So
s5Uf9KMr5zDdFhh8slI405lkhGbSjvaJqHknShI/ADp3h+gQL8Y0IcV1HZRp/916QEKzJrYyqhO1
0haApEiAh32mWaak1h4WVRuTOQ/OMjwZArJSDZH51NmdRrUfDkX4oC9tiNbvJTorlrP4xcaq0sLY
0Iwa0xUvCS8PntogE/MdYpIhPt1Ig03jfFUnLzapn21iDriOKEY8VGR/e/BN1C1JJLYpGbflrnlF
jn2bJiPI8wNW93yx8dURNmm1SGqcRnZP8+VM4XUYGsmWCz5ztanve5vY74YAAhETMC1kCZZP6hVr
3oz/FQQca0kkSRQE/GTEs31K2q7Gpcy3zWPIqEaK8/IaIwh1F9K+AqEFv6QpuliPQ64ORRVUV+zG
lz8B/Zju6nqCHHMxUdPiqgBvzDtonFAJWc8pCAF0QJllDkwczxW+Nry9B8um7QhwapGs0TNO36sb
A9qvH7vXd/cFSOwT+oiIefL2ftlG1kaNn/6VZhG8EkjtF5GoYtwU+/bVD6UIEn+JUXu+zu60AA3P
WzQhfKjsOcOw45equZuqltUbk3sIdC95hEdQbu4v59rgh75TJMOPgp4n7NM3c2qtmD4ltSGCWTD3
8pPbgLF/x3s5ADz4QErzxM2z5jln06gxlFqsT0ah1S4rjsobv0eazeCroVwovv1TWvQEdJpYRlGq
6eKp6QPfQ+6nqQtXL8PxJAdxzEkw18ioyyJkII6aH4k7cI+4XcfVQOJRpkaNi6t4+UHB+ipdUEAd
o6zykL7Vnz0tSS+AW/Y2ihrOnGu7wReLcsXrVFt9DwIigrmdq42/5vbwz5i/6mr8PZjJqIoEbNTT
AGiQavOOz1EsBrRV7kJW4wgfcKZtLk75Fy61gjJtxiXHuQPxQW1it5Iv5x4JUsxBMVk5LEu9YWfg
J4kzmqQyEchuFgzXLd5QQZ5F2ypJXYfjn8DQqqIFmD6RWo5fOWDn/OeK60MkQP5zmdpnV7Q9HW4y
muCN11kn1YdWdDuAE4eq/YsfdGlc+eFvOA2kEpvXj1Sjoa0onf82JjVd5cDIwFUjBHqsOo2hiibQ
yxoIWbU7ZWGa9BNDFGjDa0lWJBzayf62Uf5fxdKL3seBJ5bIQkvTWPIlpqzdEI5hzg48oIV5fxgt
LtvrvAWIKuOV+HLXDbE5L/aDyiOuhWim5Ly/dEodZK1DOojaIGVy5fmLeIZMtazB7nZxR1zp64nI
NdgmYTNWQC600nC0+qCivoQkdpWwdB374RxEYocc3yJhoFSou2Uj8ehEKTrVbnReOeCPy9/yZiDw
1ecGrzRDgbXbbKr4Z4/J7etQTejVFJXXiFRpa8beOR0STtKSFyaaYzvPFtqNrYYdaG6KA5ahaAmn
U7ZFjzJKGLhjlE9HYUdmBo2iWVW+j42bKLN2NqofMYkAv819G/qwDRGB69TqFRhH57YtbAwiuUvx
gPSy+txb9eJ7ZseS2bLidT91R807Tmd3C6yO3CZoa9gMTwtQgxc6mgWycji9N57kdUyKXfJIRxt0
qHqobvOtjzPxl/eQ4qmK9NBoV6laDHcCF0OlLm0Z4qJBHw32KI/vJ9mgZNxerDmOYSqDDG1He0fo
7eP9cWgsTzAVZgkQdDbdaJTyasoXW9cZKnBC22oRfeZTYFSzzZJZBJ8ZDYuhkDI63RTngsUTkYZT
Eo6nBTFUJhS21fMweWANcZ7ohmhTG5T+2mApoCQZ/BwZP+ZCtqNwnKZ51d3f9rF5P5Bp2fdhXDpF
AAeaBdg+pEzDinf9LUnuloxzJb2pBWT4anLrCsf7yO3b4xXHsFquUZ5pwJNSoVszOg216jx3ja0M
8DUOShTryeX7pf49TmotRMczxrp5qYynBo/A0UB8/H+5dC/a+sxWfHi1T1fhYMDH8oD47jW8uW9f
/iW8OpWN5MmHuiw4GpSyhrpIUFR2jLFQ+0LZYa2Mogg7HuKuPZkyb6ssTmqHWPmpECS0Fgwqkx5U
RcqRd4oX4m7NKPPIcEfFT5h7tO0QsfkIkVwEX5BWgXmrybWhR70HGY/8vriCoslMHQ74tTRw7069
MYPsJa0LDHakdmHoEx8lsHQ0dYMq1Bvz6T7QkUGLYBWkfaQoIMzD7NG5jVMvJThAF+Kehc3PpVc7
n9Jyy3qEGfXNLFu/mapwWsqr5BXiyqeFHNcY2H6BB6soeK79xgyGkLdMoDvc0KL8IYyuht0H4oXI
v0+cmpkyqR9yNip7ts8/Qa7nZw/7B+yhPxfoPecLspPi02eZbxrb27Hh5f+1c9p7JbXYQF/OUc9q
Qj5deaRt2XdzmGW4g+NztuYRHQldyvA2+PfhTIgEMm9cTwMqX14PJN6rJJm2G2uQjngUHEMPMZ+a
7bNKRG2SD6Tjl37x4RTQouXC4GwOnL/kXvinZmn/9OjeFcmumdETNQ18UhLZzvMibWX2z/G8SNXM
Ck2ryOS1mbpE40ieZn9rmLniJLBHzBt2u3U1uOVAuYEbvuxULyadi1n6/8WnCCprvaJ3hfObgj/A
aCbHvBz1pSgCAmXnzN4O46f2RYPUzTcucgQVn4xL6zL23BR5at4BSs54FVr7KL44N5JouYOqa5n5
LxK06lgq5iLr0+rRCH4LSMlAMst/R3w5sF43/Jv1b22Eu4j+dZ5HELoPjWl4++2PlErlc2a3p6jv
H5nyNmOZOZSP9+oBn39hpe4RMlM2euQSKc0PrU598Npmu4krqTRUXLYl+yXgl0Mzd+2G8xl5VfnW
W2nvIPjCB+E497ReS8aqUjN6sMhSvhbnceqUXRsFBbpY06EBHNfttIbc9eTaijHJsG4JqsauAa/Z
optPWQpB3PSq3ZrMSXmkXfH2+GvkrElGP7vGeEc5BjidBXoBYsgwRt/Vqg0sDSwpGTj0c1EbR21+
HWWwUJ6cLxhmjh4bNBHBNmar/k4U27+Kg5iBMwYn6OT/8FyT47k9frYSn7VokJj1CzpnA5qpjSY4
w5yeJi/Ocl9xIz5tGZcaWtszmUrESIyIfHMUCyYU56Q7nZtkJkEyf592nnOiaClsgz1+O7FB1jNu
03VDFvjJKw0Ywi8lzQJ0jjrivEZ90gt1iy+uei3rTzlFZ2Bn9M7Czpa5o8JnBG6rr5+pZgGyiBqs
W6brLYdQbP8QK5+4OYREbAi+jjrR3Yx6y0qWOxSDgBg8SfQ7QKKNRjS8Koqxl5zjmnwOsH0sJ1l7
o+4LUvZwaWJ+wTUa0pxCILq9U/Y/C2s0eDAn/DpGuCwsMeFmiKLBuQULlPzElffLNhTCWR07p2Bo
4xy0eaKkaoZau6DnOyyMcfdkzQpddqYpj0stf+cPaHvsdD/b1ZBv7Fnz5F59YqklX9VDdjLwAKjv
Ptf/jWc7p00L3ygdBqlKvC/r7nejdpqncUbi9p/1RZwEsxUgEjELN9+ayhmwAXU5c7aOK3aNYenY
cqu39hjl+OpQwpUwHVHdFsUlYkdCiX35KlD3D56MjZYAOd3JZ1b7yGTQYVsSoRagRKfsck4RB1Ku
/fU8HiIp9aaHYm2xdk2XAra4DMY6eUKmQPYhgDXai0LO/RJy+FwsgwPzcEbGcUDBcTYC+wqc815C
e1DQcMHptP1IJ51krU95HmaOGpZBElXfS3RizAmf16djeX0hFBFN8AoZt3715oqOTzIKD6mQNCSV
Bz79jZiSwfa8CzsTfzzX6rypQjrFGwRLj1QzSOl/MeqUQfaiLBajX30SYKaDOhVaOw12eSQs8YKQ
W+e20ToJbTDaJoiynMo0ylzrpYzh4qYrKElY8mH6Y4gDqckOXEEDxLkP53J7RM8RDku62r10XGKq
6O3Rae0YYNUL33A03YQu2T6xxRSCT0g52xONKSY/nuLuQR0mTPJmbDBacrbeFjb7tvHsy9xo/7Uf
+ogc0NpOYfSbajzo4wk2QOBWbGh8+bxyMV7H/fgZxHCQ90PgLNECBvE0HvDSLb/JCGhlWCLHjx37
Z9066DxCtJXOSpiu1QtgYG3Y5FtZTRoOtROiJOc37svF7iUuPUsSGt51J0kbI5CQTypp9MCtwMDW
Ifo4KB1rqJiAH3fho1lqgFUTx3r/jDTWnIYG2gDV3E66+fA0SSn14D3d28rFpn0D7FeTEUjNy0qb
+MkUygguM3Jx/72l1bcuC5Xg8LFj1g1/PUapK3Y2r6PM0GLR67TkgWFtENawCT7Y2omid8X/0w/i
+9G+xGJ+fwP4/KY/2QBQxEgqoJMJCNikNguMXvgh/TQLQBevIQ1E2WdywuT2EU/t9BtuR/V3Im9w
QGXHR2t68rWKEb1YbV2KpnqfXoQnZ2r0phM4KZUCUi1s+nDoaOa33ADXeiGgDE4hjOsBuYGlSpGw
pnRVPae3X9LgAlpiAyE4E3JsB9r0eKW+OzuUxWYwJIj3Qx65LA5AkC4h4H+Qerenvxp8XKX7pJtp
MV2BeKmXy1Xqq0EHFTuu43f/NfZqK76u7zR0s3H18RCH4+i9lg1FHMiT+MkXDNJ5Ej53zsv7TFNn
Gj9U7lhA/KwgL3wul/PTheq/joSFxBE2N58Dw+RKEcO+XKXcvwM1F4SjFa0thUI4YtkcJuq0T63J
3CImYsYG1wHqztaifPJSHpiBL9RC4HC+siXJnnpQ3WAr0HQtr7jOk3EaZDfRgvbhNefjJd6zGbqr
DtVlRVxT7cz4Zu8PZsMeyo6JV6k5/8u4VxrqZqR1PXZ8zJ/GqwkikPKaAFDMhFujP4EU3ubKxZLv
xDAmuvSK7ilwUCGLLQoiXu6LlLcBDS00qObiyzr1TAhAOXRogpLOVV39PhqD3Ve0ua6zvCH3CpMk
8nMUe+p2oGZHuY/cT7rvIYGB1HDbqazOmeCD9+CnIOv1waJspkyfWxGXgfJh7gR50wv8q68/XvhH
W4GN8x7URPcJfdmjTNIovfioYtW8fPa5edLdqtWtNOwD0ouhX0fbzGD0j3ZHinaq7eVw4YtZotyW
CbVpgnj4/BBsUra/cAxQ1BQDaOc4peb9shJGBlCk8we8DlgYJj2XM3WVlJNCwIwK91uA6d8+wIGA
1XbAAG5pMIp3uj7CrPoBgRTwB4h1otabMufZXYP/2LQc3+jpfOPbAaZyqhFcqeAhieOPNfGYeqRW
m6JQS9utCK1KVEuGhLrAgiE4YC3x0bc60Sd5nD32dM1fuYsoFxgoHVCHkh6NGqJoRY3LKmQwYHJ6
Qvc+xkltTOsPywyaU7V2RUth4C9A1wGv1E4P1UmuwDVC5AAGF/mUKudCmc8nzV6nwK/DIrWPu9SS
4aJNsnEFqVl3/1O/rGpfszeem3Otp0E7A9QPKwJSAJEKxUuqhjm5Rl7zyHubPgaNTmcZQDjUpa4S
FknulTbwLKHPWDzsWahOEdvhGN06Jz+JlQz4hpznzbZWnVefHAfxDrOUcDkzVR83LSTUL99DiPA1
XQ0Mg0LLZohIVM3cMT30tz2viRYFkXbFqs7FnzM6Puj+1zMTvLDaZizrb1az2vQTuikshcZZ4H5C
S/0x8Idi2ea0TnztO3LYpCBMtu27vRIOre9zPdtIGrlU+93qVEMqNIL9g22YZMEAHp8nloY32doj
9s8R/rbpTgkmA+FQLgLaRax0YTj7KvxsNGd5xasS6J0zHkIo8IdkxqDkSPetpPeCRrFktyYoAE47
y6tsksjg5lKsQfJ6fOcrsuKU80k7pX6rKnvm7gMO4UV2oF15z5uXKCRSC51byuts1gAfggesGNYE
Dx2jDVI0gUZ0SMPE0MaZ0GH1NN1wCIqGYLSPouCJAOImvEqOVmqZpGzR+SQ0LgLEiZmAgHyEePVJ
gzcY+IENI2bNwYF6iJNzzgakG3MBONSdm3yiv9PTMwSRlFoWYflYid/VZ0xgbqiagZN8lnZDML2r
+k88lIWKstpunbL+C/UYlk+E02cAKsSUT1O2xzhFaLO9Poze3VIn50IPkikMwN93I4FppH1HlsWk
GKshoSTBBLBMaPz1Shfn8r/UDyKU0d8qMk+Uit/omHhJWFA3Zv+ojCs+ozX0wR+SPfEjqRdCyTri
bjvL8Vif8EaoQuV4JBNzU1mKfRT/99soh0aMNEhJtI8ZomvtQ+4ExPN6OfmM1H1epqxxjr80cIla
GbWv4jG/sG9yAeir9iOel8Xavmewd0N+Fp6+7ymXgc1X5Zcd3BIkcoTrAv7bOHPcSLa+5Z4MgEXv
TrbHIhIP32p97/gklCaMtLSF2SUJ0aCRBhltFgLaobZCO3axcoTNpVzX6QIhdxjutuzo7ICmb4pR
G9gsWNRzm57/rF9i2SyQM+FVARru5M1/PPuPEiXW/fL7IoDW7qqtGl6/FRmgHyS9T2MvZ6Z2Td1L
4wZNDc3y2ukJE6Ny8snbQ8k106Ko79qBz+c1Alw7+0GPf1sd3/plW0Y6JOioakwB++X+nv54Gs9k
4Hb+PrBpgir0Pzxesvsq3x8gJDPFz6pK2VNHLW1fBe5wFX8aqCgixBjEhvlDTkzTbbqVfAfp3Bvf
R2mTxVXZjfhwNe8HS3RIJSh0C+wOpCZSTW3knG8zF3bhjPePmS8Gfu5J/Y0yajupbYwG7vES/xkW
teY7s+tgHB5yUGL7k0fY2UkgHD3yzrOjGkn1gI/OVv4tCBd+sgmyi7Nnxolnk3dsPoMPe46oMjfr
HBsybgzFhYHMQCTH9Kz2SdWFmlWs8Pm+NjuhP7IKH+xehTEa6fioAyid2PRp4BrgK5J9GCSeHFWL
SXOvJI8fZwi+Eb7UwiLebAH7GSeQ0euladqRRRkp0ONnmIoq4pNV4YVDJ4rSRPu9ViPG+0zWuptm
qP1pdu0f4bzRI1DUQIJgWbtoH5010ui09Ng43pg2+HXehc09YySkp8V9J19OdNHNAGPfw339I6oR
f3N89Ww/pFPaJ79Vy9Nn7V76iqk/b3Nrps8DcEqIJs8vocNaxbR0weMlenJ2TaITg0Kl79QZwe0d
zmBK8LK9rpDiM0+S2SFCZwdUVv1CmylsHLDMU0azHKnGsWwqAoq78CJgtsM87e01EM5bioSmM9cz
LqfglhdAgyjVkQ7bzlZJFqOUksfTHfPyTiRjFrifUMfloVLoWM7t+3SQ69YZABRL1i79WlT64EzJ
ZcAeoE/ip6mSon/jkp4mEB+xHGgSRX7Gsq5Q8YKFWaRnZxPaBJ2xwZFi+yTfAStWM2Rt8LJiqBBd
8qQLMO1AqwbASFjO6Tj8BxGnVf3hVv865K8PnI+gD1GUhoGrtEkIaxLa+knNGO8eoo+CvwNyzbeG
Xb1N3QgyA+eUzq9mHPh1WTA5OeuxZQg241qtnf8goD74zlXepDCMSV78NsYm8L5Nja3fllFO/eAR
rwjMr8Wm6QEuZFEXrCKtwwFukRXyb8rI52CWsfLY90PYatKbxEno+Hjp7eOrxw/6G9daSAzm+gde
Ltd+Rt3zlXiLSMDuU1bNCZ9CSgrExhI0ref8fhkPdH+vjNpOm0r1yN8nBsQt5Gw89pFhBJm6AN+g
uo3bIsVeRAUK+yKvKIpDUf+jWx5F2dtRH18j5jjNN5//xJ7WpWQ5Yoyvo1if6O83JMVzvQ/FUl0V
PZPQ7jFbeBt8jODWIYHFZUwaY+/UjgYY/hL8fMUlzpeZ+EzoEovPe8garjWdULM8MPAjn1MrsseE
1VFJ+FvPho+v5fOtsHr0kVa4RZ7UKyeAmnz9Tcbgrgch2UTZ3ZWX5e0XfMKRTU2Oej7Oh9QLgg0o
B1Mn3ObUCwfA+VH3VnQnP1eZLlyChxy5yi/zwE60ZlQHP+w7ELlxDjCBVJnktD2Gq98RugxQeeng
J1trEHfLHV+U74R6AiwkyDga88pt29eedB+DjGoCLABMWKNTnar6e+M+DyrYJDYlEYgLKqC1hFYV
pexWrDQcIOnXwegPGddtyfDJezqORAuybW3IS0Qhux9e78vlPIcGrfuvb/XaPBqjnuHfXaxYasjh
qn/zLYnRdd6EHFZ5XZDCYwV2la6bVvHYcc615NmXH2qxyXUTm858cb9jNt4kUkEgFU1Uz9zeajQp
68pgtVc6avP0D+NsrAF0oiihyW+8ssitQvSmMCIK4jQMzb1Z1EkocMS43hDZt+rqb961TS2Nj3pC
I1JOYbIVgOt22fAdt163woU4QAUTsrWDnk+UX1hJp1BfgBwDDQ16QyfisHczYvc7vXKEBFqOVHiE
yW9wqiI4Ir0X+CdI2VSZYVCq0u2EvX3zOcASWlyou35EKmn3k0M6U3UO+gd8kLZ3P6aZUj6jlf13
HdCsbksM34aJNt4GC16tMWeVLKvPT8nvkLs2BjnAG4B8oOIhBcsOVnozCTldODsz5WzV1QkrD6Ai
noubx62zEVaw0yCF5m81iyGyOtfkVgJgF1nmceIJ62wfQmCkOlhwLGVRvwxBWar025J1gU1PwPub
PX3nmQPnzaBSf43RDy7BeDl6m214s8F68k6gMt/9Ls+q4FDwgEUmHpc+N3tfh9SqnjsGvV2NYtaD
6XNJeO6eH7VvbnRC2ZsjBBZlLV+lO3/qeQRKmUseVCAm6d1DwgIsoWayRjVx+1pYHPAfYe+KjKl7
KvQOZbCunWLcglaQ/S2xIIt6TEicDPxnCESz/AUzLEd9R78CeVDnUV4djwYz+En+X0ZqRaVW0oaE
pZkg8y6491m61cU/TfsKzU3aqtWkOA8yhVYrs02SjkEOy3Qh2SC8mrWW/dTbJRi/vU+q/seRYDSr
uxHDLRZWv0GjvYmz/VktJPMrJzfgTtINVroEz62oAdb1ohkYJQdfuJWCxivxN0m3EReeDm1zWmy2
IAfGMVeP/Wj7qwsJgAzAzTAcKMc4V4sPzCzHoZysPHIsMFCfq27wENuB5GfaXoOCrjdjUB8iv8QD
IV5Y6GYQVwsTpBOXG32AjOSS69HJ8cwDwMLQpFpaC0EwZLicwAfRN1Nyy0aPpgkypWBrlORrrjFt
PoVOGeJXKdAru6yFHjeYgBgr8B7w7DExNh2M3oZqX3wZ6qfMXxjC2fY53b5w8dAgVmR05ZAEyfok
0ZI3i7ED+NF6qdTEKO1KOXDxL5ntHH29OEDXisECop/qWV8zsD+MDxgN4AWMDjqpF09P8PPXbRPF
iPQ/S7TT3ZDoVnWsHFlTwinRJ5jFOvf/A0ohjC8Z7XDJANIDosOH0XYPQn64t8cJ1V4dc3rNWqsU
w779BoH9aOfUAOM3L1+YTYPMLG0VJ/qDp9Rpe3tWB7hdGcmX8OnZy2rpVkSwtzksiH4IUGLtLXos
pJRprWHzFIelx9fssW9ZWjW+Cgt6YWPNwF1yibS//DIZ1ajs3z+dXY4rEiLq/UhPlTXfFuoLgpJR
zI2lPLFVsBkPDLS7nu/2xJnCecRIAuSbG9eXsACv6AFz0fSpBure8BKeZ0hAuqkvHcRLhZHDFsw8
zvAH6t+/M5WQh3cjSVD/Dg1DGQDZIRgY2J3lktk+7ikKMC01OVCWB/phrCOYIeSons8VtMLNcJ9p
KCP2pJSHrVo8MBHwCBwnWLXwarVnzADnOeC4/6eINVcP5f/1aQT4J1//KqgkwbctebqnTtGBnOHW
HrmeDPyqDjSDWxngGKBhuW+qtxFfVufTlnZrRWM/9/Qca5Fd4Tvfb25mgJ/3VKrnYoNXCmYPigoB
dEuBRYNwIpUkx7TSE31auZFyQvDyCIcupCddWQEoN92KW1fyKca6y1LQt4W2vfVEZWYAw40OAkA9
LVogqg02pWwyuWZVxW3O+NCw5GEne86ALVmPGLTfUm7tmvwnRsUPOVV9uoGUcTvBB3QSmOw3tSqx
Txi0ANr2QxMpfQPazNLrsyrxVbpDJGt4UgOlMmuLQjXeugvDMKE5hKN8h7xvswc6YB4tOScraM7o
di8iTKGMNcHubPod/LWeseVMSHvFms8uwXki9M0LN2EyBVIaRVX0NDm080iERvuuHtAZbXaw9Qvo
b1jbYj7HoIo4tbqXko1q8OJhSLfBLUfP1E4kB2Ny/bXBqGKUvKy2xY73PGrsqN9xaJEQoM9nzIlO
XN59YWwDMhLsQ/d/KE01gYHmI0+AtLD2Fp53vDw43uBSAXQwAqoQXR1M7QTUlN3bDC61vKZknzUu
SMUGZ/fKw/LSB4FqPbwhPJwJSrL0YElfa0/J8ep2e+ao1dWXPHjytyPFCstIdKBqRGUgLyTp7AqM
x3D6K26brWOEGkj0+Q48DmyJTukeWu+zRP24SXvPADQ/bPvdePHJHmGRV+4lLsgCxkFg0zy8bmyv
8zF379gPmkVmnitmqzG1frByYnelW5VFThDJOxlweRlTj/KBPYZxNFzwDx3pq5nm7Gey+1iheQvu
qsoDCsG7QD/Aw6W0lwDJo9bLtQPNgGPzRQmG4KwsmCMC+5iDq7CsbNf+u9Ehn69OcGX2NELmLvbH
VYDLiuAji8fJEbcWW57/++qjSBLl3vxSo5S9ja/txVyiMOuU3HHk43zeBj/s23lnxjbDEckoJgbr
iv4ecFFJLDaGyAtfLNxZ/Y7DWqlrKKSMmOm6O1KUrNU6v6UZLsexA6oe2sm5aFtbCNply2toW6dA
AzxaY+9Bd8OK69w3TUezo3LBmjn38kn8UBk6EysQ6pXD1LCzU/oy80cPT//4RioTp2C/yUSQfh6g
CQN6P2pmw/N72AfezYzv12lu753qSnn7RnOqVLFqlz7GdLvqVubr71IlBk8W+k1J5eLEC8OXeD2I
0fThmaeSxl2GF/CM9c32oxdjAdG0UE8DxEjZmXlm4Hwpa2T8WARhBAbR4z+pTAEpPjFWVgUAfKTo
WAIpTdA/rLeoXVBR99E2L5h6vxKX58+PbaRiXihKiqs4LqHA6y5+M8zU7G7/wyRZv1JodpR+E7k9
8gXmPBJytM+UyE1iw+LUgX4C2656APy3yQCsnXMShRUBlrzKQyU4W3I2xpFItaujBbVP8xaXr5fR
NZLjwjBDA51AxxSvNq3Gchcoq++d7TABj/LFT6kER7JMX/mOnHXBZBJ4Cdij9XliYOFSwg55+Rbh
4nuoSi4iO3gVhT075WYObRcIw6qL3juiY0gARtwPT9iNhlTPJ74Kv6/uuhxk335GvJd/cu4CmACH
PkejqX2Bxb95B79pEPEpiynFxgxjX8AnD2LFJEfeVxQQH+BXlpLHP9MTY7+Mte5yio+Paqp8uHtr
OeACnz+5MyV8XcwXXZbBHOYMXHquBJuHWTZqVq4fHlBQGUPkyAIhrYV2NpKrE4x0LTXe18O6H4G7
gRboG47KryLTPyZT4DaieUera5slh926hlwR/B7V/+6AnQXzep13qexRXo/jIj1O2gGR2iCkWlth
Qy5eZK32pJhoM8J63gJiWjVlOHbDtDv0cjBr6/Z4oSMg7D4RWOLksvi6Vz9JcTWeQOuBLyUyNS+p
jFUc6CDjoffcWLxzmI5s7/9XRJeYWCM2fyRgSzPrfwC79ZF8tmPGd51Q26ILbRXkVyA+TpuSKVgA
OS86+he2rQVedaofNAXT8nQjLQDIGfxKrXkEJjx0ufuxnLnzSymCOgzBN4GgPP+eOx9ELnEqNLRo
fFoPicM8wbnNqyyduCGcvZVqRuIGNjCxNVhIDu60BXIOWb37IuLQtURxLSODLL+b7JgAVksBCunB
KyHKmD5LHw1Ew1VKSdQo4h/VmxjHg/L3Vm2TBFKZoAIjAlce5cFSziiM9KdhgiA3fOgA0iZn5BTY
syf0jH7lwuAUAFh78It/XPIHdElW0JkmbSuLc5m4elxIuhvqbnqJV927A1fBMOIlbNhLtTfx7c0S
3cA+mo9z4wgMgY7V+mE879wseEgFB73vCFtkhD1ppvqMQqwuW5D4HGZEUnSSTur8KVJjgQya07Wb
0CCucesILX0DSYK5PBMj51HUjfWYdCPkODz63oYi4olSuhByaCTVxVmdrjpI565NIKyWhbHOKHyK
PDzC2jOuAGWSW5gEGAV40kogGd2RQXmCCTJsGEIVF4PT5zgah09a6c+r2aD+vFkG48pAUAcMAwtr
AYbbhg345VnncGsOQUCSxU/RTQ+oNwhonZyhs5h0CbH/dj127jC+nHkRkey8e2ElpZbk+cHUHWtA
HSj767/OIRuDTJVirl92i0lrZ/3FzeJGS5MhhRWh17NvvCDak8dx5qz5+uNRAcbnzFxrWMt/ZbVU
gF1FOb4LfNw/djisUcjd2CCdWNeYOxdGj+rm/rIjOec6jlZ6N2AAp4xH2GdeMomqpWXCPehzgm0k
BJqDFkbIxArw55VlsWmU1/6ijq3RfdtZsFR326XbC9TNKEhpf0tGt7PqHBy3kT4MTTPSUZxse/NW
ZdX63vKPytBfdb64UPyZ8/iZy2lYjvykKqxvGDaI85cVjqlqGVp2xnyZLcG5gGVN+XD/bTzucO8x
UCPbi4GQjwVWqcNNdkE9Uk6C57g0mSk6rnkT2WiV2698LnV+2iKNCMzWFGnmMDpHGwz1HVJHy7Hy
2feIqktss8KdR4pDfXywljeWmeumIe8ATueSPfHGe7TFszNa3SmqzbBlYI467S27pJ4L2LQQb9WC
TFXsNpb55gWKiknJhLCJxnO9yoTKZn75nHp80DVy0OcEjEbPhPHAKzsn/Y+W913+JIrj9xK5SXO5
OgfuhNzvV9D6BsEzmsCqU6nHUBpvvBgJWHR5nxlLUJi5KjgQg8MPw6Nx8zQMzHE8PPr5jjCvEzu8
80zeCuT5HwRghO/VRcNB1nc5+HbLHuI0pgY+t5DJFB6JrI0BRawdpPfCK8Rh8p9v0jRoYbZBLijN
JI70dYmlCbbJ+Oj8Oh5BLTtXy9AFB+F8vASL8kvB4o/OYTeFJ4eRCnUcdxeN/m/oKyGBAhrmZeKe
i6/O93kT6GA6uQBWfuVumqjvtLGYmhs5b51ueHCtKMCjbK43qh538M9z0tpElLWr+k8orJAfuoQa
h0CRfVaWhnwn7D9oaZk331fhb31HuJ/MikFdPnEWQxkN2U2ja6ohNdL3b99oAliEX2U1U+T6zgUT
mQVGDdzbzDLllTqu+pGMNCv7AesO3tXBdtwgzLfQ9Q5aLLOP7eyc+ttX2SL8K0QxSbVnOQJvEYvw
YSCTiVpvanDmDc0lryXXV28S6zsHtzIrt5wJHlLE+VmAQmkti8h9MtzbXZb1jGcLZYCZ2DtDGwqG
1cY5/laNBXvr2PmuoxI3zGbRdmRA9F9l34JOwuB0tCDpMOZOv+YPFETB3oR4ZhCtB8E4FTVSWiEp
NWYUuS6HdR0IkID4kYeDNWlYtJ20KoH/kRqJDMMlFpbvb9w4VTZnZVR9DYRoHIkH2x/aXI+sgAn8
GpthYecFmchtwt1OZ/eTPmivoyyO9RRwXJpxMW/uc28FAls3hZXrqg+ePbwScbA/Mq0S60u5hhHq
MErpxk6EdaaecqWNpC7v6gafb6bHXahzEVSGJgY4j561hL5o0e76RtrEjVVgIEAnREzUILE8E9aj
2NnnTm1DDsiO8kC1iATDKI4uMPY2WRUwkoKyLxOKZJT6BktMB+ydBYMGmHkBSbBBGBNu7dmzAgRA
HdJgmTcc+3Ko0yKiHcveLMC6aQc5gKShC0rC/FIxMrXzbMO08sHbpmm4YIUY8gPmv+vjpQ+jLxX4
ptqlox2iPpiBzA+8ZeBXNWsm+WY1RXkP5bW/YEydD/X6Zoooa6k+yfJoFZe9fmM8qo+PUvbHx5vp
v3pA3lRYKfy3ekvLmW2x7cpWKy1W15m3KcevtpPbqcUHSyz/C5DvbfnSFGPhh33RmHKkvFrIHOfg
oU6vCsFdiEkpM5p0rxSo+dcU1CgHPXA/I449oYjQkvrq88T/OaWc3+iLCCU5i8JEYrJFuKKqEpu8
qB9ZxEgY8QuTKVczTfA81840EoQBkYJa/rNVqALOif0x9LqWRILUScAqm/1DxVk0ASCD/g6flqKT
XM2B/yWgmvlU3nN+MrdRJEQWy1akIFnSc5wUL0hEoH8F/L9jDoThT9+a2WbCu5DTyx6apesGRpfO
i02LvtPECfPsF3WVL825b1u23T2IuzBOAI4WU4ikuZ3Va+3ZstyZgdqZvU7FjZlQ3mH6IMW4LVnD
QpIoGiGA6KFW2kHDIYiGHpNN0xpxmWyuHr7lyptRIHACMfVm4RolxKYSsGo+r7FHOvJAauU826qB
DL/Je2qE0+KXrtY1mZrNRgre8ez7qxuvwYlapwN5GIBwzpvRFv8aID2eueoVjXv54GCAmzM8gQli
UwpkbcKylxFBqppUsxe0pSV4tfwCCYx0CMdv1+LsyJhgNc4lA08+r4SaMT+ER+FY9flJN1rrTter
dS5IOJ+/MASgXQ5QxaQzM7e4M/s3UKg+an1LTjEoN22MbZSZDqtmg3SZiwr8pVOJPOkqBBDbsK9v
dlOo+/67WMnGqjWc2ANeyM+0C7DZcHzlrHr21QBwU0aDrAsKOdMiezT16TNqsHkAjbQtWZbONhBG
M5MZcH9T6InRGIOV2P2gL2+GXoyGparWEX6qrZrffmvizuzZpCdZpXwNphyhQzuQrcuXGoeW5fbS
wZZnlNnYURHq1d7CW+lw3XKWiyacEsbkPtf5qdVdwYGWJ1t9yolZZR92pNhXHYO+n0KbLfMAV6KB
HVKCb4ijDwqaCrFjzqzWWQWXqEgkCN99tlDDXaMQIRZQjgNstxuVvKNgZsbHFLFd1BacILJRDB10
dCLhOrBgoVZBioBskAAdEC97gmBCyJYe6u57brjDoLMv3MFLhqlgeRElSZbaNOOdOdbaric4bS9F
M6W0uKfgapCN0psRJu98XzVU9W+YY5sVSkvUKdv3ffXmDQhNB48NTqI9i1H1wBNxSNJt0u8QOh/5
A5D6oUe7S7e0zLvc1D0sMW1ZCfPE8KnCi2pAqDrZlaA5HcTa0bCTsRwSsx9IeQb21b2HOx666RsD
iM4fE409K9Ih+FF9HvH63F9y1WNVIxN4hIX5lCwdKz2SHsSOx0WKO4BXp5tS2vKvVvTORO+DxFKB
8iU/Ju6s07I9zBfuQVWqHO6enA03x0By5XkCGFrRoUAfKDGW1N46j5nUmzl4JogrLHIDj9f+xrl4
G+0jl6U9WYk64YTTXDl5a6kR2/qnpUak5o4vlvqxXC0MotnA3wgccjjqGCSpOUxMaD0aXzcmcGHg
mCBAQqCxl/SvVNH+2K7Vg3zRG6I6VHhjciGd/vZIX+10mYgcYJxW2tEf3ARrsmt0RyK8a8Wlerdy
C95I5F8g2q7z4lPN8wjlvTLBYZz9JHazfjpaaeCHI9G4K96avRPveZmMGCtAUZfxmJpRMNH6YW1U
EopfJhJ5lKpuK8maBnvPJ4na8IcNECwZ4k9azwSPIXKl/I5PvOx8u9KgSUMA00zGfOYJhuTv0rea
w9a/YIG7tk7QpIBCPLwiqaAWTS0mPiOUwIllQKuBTJBRD/6LJdx0yn6P5fhbpqwvTfhXcCwNnwfk
Ad0vMbFRgPifyvHY3tftNTnybsXPpHnZ4bhzXFTeFsjuig6Yi7R3GddBKKlvM+aMOs1ewltMx8UF
l2ODubNesTq/md1uPMFmd5gcT5ZR0p+OMild4QJQzkWYaCbB+bcf0QUthaP4plCHC58emt4R2CTl
Xu5m9H5Uvrif+Lr4JbdK1+Qyw8BGR2SXCTfCobtAfa8mycl0lVfag34+i4mgOIkdaatUQe3YYoch
LVYVuEDsMNIsCc3sRKAevQVhEuye6XH4Mdd3dKZzx/z0GtPjRPnFCK8xDJBYrXMx9tTltC3oUyFg
7nsDMUptbHBszbJ1hwJxBm9D5ZQNs6QFy/kuPRXJPDsJqy5ysdNQcuEKVQp5jNClxHGPsjoKHQgt
xdVZ+ATgDVttcWC3j+tyYHWlexiubhMa9JpFDY2bpdX7BLp0qo/8DLKkvgi1SDIVaxiMGKhBrc1F
YYoV3yH59zMp8Z9DvnUypG9hi7OHpsjtz05cFS6qbhZcpT2rCfCYgGjkeKaM6+xcVQdG03IzqJBF
lW21arQHeddQd05d2y24F4oMdYz9uxom7tuNO9rkHexyyocbQCxDCaEUko/SBbiLa9aiz4Wa6YlA
lXyh9Yoh2YBvCuliR9ssJfwByPB6nc2ZVkiGNdzEs+mM2cMaMQoB6N1cKo7dmIHLkmmIx79txeOe
PRMEUF7oIGofxsjwRTCKPxYsPsIaDLCQXCqh3tVW3Zr8gObqWGr8JB0ZThL90lNwR6U7XCKgPbAd
apl1YZButdvfIzu7RuHcLgTKkRt2K1uZs2KlJXJV27xXuQgyq/o7/LwmYirpieBXLE3Zy0GAcGQZ
iz8PuY+4ZHYBvrvy5yixI1POtnVsTzt68eWITshYAJPOTNztXbbeVvnG0UBfCW//j8OF0ZW33HE8
ecMrMRpMYSXtug1LULHwrHdG0u6nnGG8lO36vCH0k0IHi9UnuTVJSVrCNgNBNCe6nrshhYMc3bhU
mU+MBvYhrgXY7q3xILsfB+lrbNw9896xmW7t90OiKh76241N2I2fn5vret+ZfQvdx7RZPmVzPh9e
j2umF0oBGn8z8k0XzN7AtA7I2U3cFPp43gslwZdQSYn50fv1KktG98Kxjmd7rS6UzB8uKpj9TAxW
BL6DPQDesW2JpKn/Uz4+OhE8b2B71J5zp5x6iJ28A+ChU/2XsAkWNVfS3bV55CH4oHBOI9VEJNoK
uu7yY2b8QdiZzP2x3vk7cxvrkDuoRCJkE8Rk7C7PqKeCtsDr4UUnZWI7YdENnjn936vtH+JfUW9G
9qxi/LQTWHu5cbawmK2TR6xvKBIqeAe7B+SvawcEalAWwvZx/0ztzYBNmE00v3PoeHY9PZbzEcPu
+Sg1jrPAWBO7qcYfzZDhibxJHxqul3zlzjszKLCY36bkbH7IfqxaanQVH6vwyKAnQVAUXRiqkpXr
pgCupI1IRbIe8eJU8j4pDpRCudzCLdF96EcQDCNVxpp0+IhgGjF4AZ/bHeWw4iLYPccYLzTNwti0
bXRFiH/gtxgvDklX6SrDzXr5G90c+eonLJNn91OXzUoaNX7ZgMJP4T/O3QIDx41zUwUQuDmporQH
id6GSNmunaG8ES80WzJWY27dS1LAsJbrVtDRcmvXwvWPmlnrvhG3b6YFYOuJhTfHAAaQSlhy+TmB
ATyNaY4REFLj8onJxVfWAEeuEynT6UqewH49w+EpemQvSGJbc5nJKKQS4hJOSIoteAUeZwhlzqoQ
tJyJWO1Ca6pKp7zJ3SDUUBzqBNF8JxmBjKDPcC1Nh71DsqZpIyGmNbtw3VBGfuvaX/+F35cRhHOQ
LS8yDKM30lp8Dm7WsR7AhgSLEdIXC+wniHeqUGmGIXFe3TE5AP05lrdO7VHIN9jMPZUQFTkaX75m
Ij/NWqitzdYXLQCVeR+Vsoqeme7qnieqXkS6eQcx3yhEe2ExsMTzLcsa/KQy5qZ/0PeZiu5OLlJS
prwhYP+GxULRpr9gApmIuLbpVmG+lAUMYFbT2vU1vjMN3JYkYAkzHYeLr1V/OTqK5jInofbSQ65H
/OfFvD2NPmMVGfgKA5ygkf67RmkEvxsX+LGzxOC2uuFo/8KEAukqttnNr5ZNDC8QS2GJxBAVcpFH
QjnFY1y4ftUBnGj9lzw17cRhiqxyYl1brSNehJZ3/3ZZMQciOiCtpG2/2cahgHO1KgPtns9RBZg1
sW2ChQLUcI8YeTEQBp1StfZauBNak5WtnUV7GOu1a9PA3ZEWghKCsVq5N48qx4EgptyOXWPORTso
98Z+eYtx92H1V4V5LHmUTFIgcCAbwZwM51zddkMPkGvDNh0rCt554/MzgmnrIgo/GId1BGsJUcQZ
yq6M0SYHc3/FRY+1OrpKtxotf/T6pkJjDMNwrGBMmiVCF2WVvish8p5T3CyoL9wVFP1wLpQ2EAu7
mp2iP7Ke0Cc+4mIy/HAt2DrDU5jodj7bZFzWcQzI+wmwNCng1KVaKYtkhRVyNbiUDxKhacWMy3QR
CpgyQ4vgSKDmbhDAk6G7WPNWUrsp9ZV7TQ/HjCc1slNJ9qDvAJ1M4rypxtZLa87Y8l3GHY1W6d9b
p7iwravDivroR7Od/rYJImtTF8rHnLDt3DlM5EFjwtWBVjmqe8tpVWZSw7LQiC6P0bgp/IAH7ko+
NLsvKhPgk4id2LYuhjBljWF2hZpfWH8Vbtyp/xc9qlHjpfpLJ7U+/plmutkV4qfV4FqqUNk3sAgC
byZl7bSvrATZbW7hFyFtQ4HbgJP2QvhEqW7ZYEkX2XrN8dCsmnWIINGr3CYF+Zhk1zekRjpFys5g
NgIOJoxEXbHBuyA2tJPPkyL9ClxszrpkHzTaKPbhHGJzTj82KeILBIA79m3s++X2b2iAx+hB/FC1
L/PlSywCHJ/txxbeWWcLtltBDecf5Xsi7fr9xk6JUAZ28pegRm+2ig9ia2D9T0db6+7j+PpLz8SO
ZN5FHcQ/cRulSs6v5WA0lKtFPut5RZeBI6p/41VMrKLQ7lRrXhCtoCqKKgmR+24DREigddhPxkIB
ZJAnO0lupvl2kXU/KDpMovKfaQBuhbD6lQwzOwlOCFv0Jvt3SHuh6/j3pe3+23ARuBxIyx+sdL7C
nvwAGLGrJeo5wz76V9qwzlEZq5EwWCvbROFguEiybDTctc8w9CrKkOXDnsbSHAdYX9S8HOd6I+Xh
iX1VBcINWIZiYgjpSSbBUyaGw3diFKKy3xYBUbvL2PAqERCIMejCyXlWZRpiAoKThsJBMCTYBAio
uDvpcBzd7waUzEX0uvh50ernikgjvHhloPgO4OF6NreoS0wtmOgDCtIdzu2I5+U6JMonEdE5AIM/
IznvelzPd1gi6+gNAC487qsDeVea9Xk3hPuUlTQqIxldWcI/WLd26uvQ2bvhaYhcFiTd/SdJNylZ
DKIKFOTjMENSqusCrcBPexXnoUyBNmywDIG+ckBntjiCeFjsTwqnN4ZVjLGjIRRvGnYw4esFKNeX
BWZIrEaxjHRliwbCjBUgZoJqOEwe+cduUa9YvqbtFqSCk/ZBI24mA3iZtA5ERyl4o4sf1sqNe9zw
ut0ESIYtE3HFBSMrzFBT0ltt9N4BiU37hnlz/vpPr7fIyx8jPAvlhszWWHbdq/FMMRDCbIATWdnx
+BIh/wbB0x2oA0LUEXWkyo/GmdPHuQZlbX5OXUXDP/BCa/uy3yxCX0fO0skhYXoN1EfCtOtrRLq7
0wStgqOroOV8hiSoHX9D6CwIe8NvZpUxRN6aQKr2xOk+txM6/cInwC7USjXiXyH4D+9ew0T+R2a5
Ue5cBw6MwQaRqbUWryenp/EEQTh12uQcLKAjpPqQVy8GUaH7PlO4zWPQDzx4kSBVWwMwF2M9r6ry
HZEJrwT/jjEJQoOE1m+2LHHxOq7CV8O0RDvxedYvxSFvlQwdjY/qXuwuJECf45n8Glx3ON5Fxfcm
fk3jbHSXpu/ZjLzxrMFoZYCTZCz9sBc8tWagt99qs8HAEIh/coEjx0jag378FSX9ve0ax6h+c7Gr
bkAyAmCaB7t8OOqpAe7GEfnyzTxZtWBvKqkrpremp6IHshdb9NcgG6mH9sSeWy+0oPmEucVPmA6i
4XI/i1rkNR+j+rdaJxfcq44+7mDJ6nVb01vuxQUj0qidA1KIYbhs+Rz/r7Ntatj65r7tDd/8QJvx
zZr+VEn7AVr0YyVLODljpKf4GaWEOm4xGMA2g/vl349MPtsL7eAYrEleLkoUMptfhTii47vTdf4C
du8asxOJwqKZiQv804BlU3K7IoEZKKXfvQxlQU7wTGeNEUAojltD3BaN0UT3mUvFOQxBlR7bT9nf
kOqWM3OU0Cj4uLGI4/k6bIcZ45gI3FXVbtYW5RZaKIatjBiIJSKHh0KAQ+nTqQ0StOKrg8klNiOl
0iAT5AHdF0bYm6GrjOT+7G2N6v7oarwctLGU3LyC7chDS/+Pk1p1leQ9Ivi3TYXYpixAmFfBWNI5
xSyzqujqNSZhNFrlM2wyxGRDaA94s+YTFiGBktvsem4nrnQi3BuQEl6KpH3bATA9L7sL0Ai127LF
hkyJqFyXi+8vAZQ957MiVfypPqowdj7T96iPvvcMji7QgCHgwkcyVH66oPXJ61qjk7vO4hlo6JoA
ghVTLWZDHeKgHOkR3zfvqZJpHrMx1z+09eDWnkEqXQ+gm7lRYOxqkpLHlUOyeYQzZahIiQbht77s
7foxeGISjl/G+viRDvS/qkBOkQru0b3AIwl66DSTId0AZz107ZywfU3w/Ltxav1fJ4FRerPgmW/U
5KUPn5lsi+yPINKbAzfWSzFf4GgIOHNrBcENOfdVLGJ/oUga2y9UBc/wZ27IZOXmiwSEidi+dEmq
fdbFciQYXlzIqiQ05pjNwAoW/TxoeQ8rOT9GzmRQKA4P2FOX9DGRy8DzM0vK5/jMRuD1ifQ18KBs
knMfEdisRbwPytBJ+hx+U8xK5MZgFB6N0JabUjURSOtDfL5LKwK3468ZfjWKqGVZ5Jqrkuu/tx0f
BGhAdXjlhLNY/VoJ+pgOUAzhEf0jrAx94B4xqiVsM9Qk7FCy082U+YiL2W0RNRmy49R2BRgb56zd
e5uza64T5R8WJMPnAJJaxUvY0GEk9dxv4iL43P1jjLeg9vvkXjTD+y9pZoEE6bmfVaVJWoW7jBQM
95O6rDBol5aAdBt+n/HS90J/F8mT0KdYHQomfr24n1C82El3BmTZScpeL3lItocqCYfl11pZtUz0
Ak19SW5eH0Sj30lfjCJxzetQxnnIvJlvVQ5CMVbN9RMkxqHEIKe9T+c9UV30zLMMZr9jJffj08ep
qMlk8NDxF6tQu+YpPGIMFZjMkG3807OiRFtILFuY4YoyZiN2gsdKWTjiuDvUEme1uv5bpjvdIQDe
hzj/bkrw9aio1+jAsizF0G4/CGYHgZCr8Ms17vD+U9m+gn2lWpY7q/ZGa/IuNGpb18qJB6eCD0Uy
4F1FWyKoZfmAnWSsCqy85uwoRKGhcSwLbyyr09Z6vLxsTiuuvOksCGHHIxhSWkBO/LnI8buDR4vj
2DjS+TpsBlLsESYpFwM8kQG7ycqmiEzvJlpJ10lannmgQlKRNOJuG3mJsKNIKRijOlCw1fLg0Msp
lEoELYcYWFhVfh1dBeilgeEzJl0Nu2qOaAA4HNhpFf3hhv0eQh9pDlRfNpKTqrAvzSnlUwR2pYG9
PUDNrEfuzEDqdIVOVsdAlA6+u3WjW/QBHqfYPDjbSih00fhQEw8OX7SbB1HsOp3jvc4AFI1Lq0yH
UzrCPweB+cN+2n9ixEAg0VnjFH7UOCJjtGUXjeT/4jnMZCSyGwJ3slE5PgeXPcGd31AZeo3LQK9B
puQ1IrPGr6GfA5qLTNDFIhdGGOQmls/xAL7TzbHHTWuxE4QjH/+h9WARx19Dn91nil/7dwoqpiSo
n8rJ2VcdZ2MXHUgDaGXu7EwLkqvKUceJqYIKsUXzjMLttPWOWhrd+nB/osMtmo0EGdv/iAGZwtb1
3h8Y2Ii4NynYzlvzaZtazZ3BqsRKp9s2DTrUrCbmM6DHw0X7SNg/wvwndjT+3o04GSgOVMgWRWVZ
UOgjqT6N+RaaHT5FT8b9QfSzL/Rbko5Jsnxt9XVUKEMlCEmjroxY6PO8aCc28BHzc+4r5TDrfidx
S/Mar1Dq3kwQcTGYH+Hykflt4SpX6OZdlksuOuZoT/Oo+OEyhs264z3LWGYwan41Sx09FO1b8qrS
MKw5S9lXP+WfwFDUmpo4i1MsKMAvejB5XrL/3Ag7wH+bYDje0Cke6EH12h11MB6NC2Rlj7k6CoiT
NEXY9pvftULzlEmG58QFpKITesfOpu2tF7shXtTd+yjD75i6E0hCvXvRBVUY9Qz701nVghz1sD/x
QhzANiMZXT1IReSgYiWnzLO82r+N8Qr32XSaoSAcoVGhThQc1L1UGWapMTdZDEPJYXlMwn11Gh3D
CR3IxPcGzMQJJs3scMKdLntOMIqp4VXdbyCxvn8EAL0wEv0TaqWsws/XsP/eyrQwbeIBfnl606GX
3Fij982pUjdhbsD275g28fL0K2/kZ2eW8KpgyafdQQ6JfSIW1XvKkkUgItulTGfUg8vc0/aD1LyU
39HSL1piZeg2nFAPq/w18D054ud+WQPjNrXGo2xUqVJ9clG4i2IXA5QIQ6VGjE/EM9tUtLebfnoi
nJ/xPa9kpaLXhLgG5rUnjjHtw/sOJIj/GsjL100MEFB6ekx4RmQjkUuhV4ZGrXMDU+OynYbJ3a0M
D4FZ4sASfJaTAzlA0hTr39LkRgEW4iMGIl6w6L2xbM1w9YD+HGFbcL73k4NiEXlrosiY1qG/pgD0
VbXxEpqTVeh+6wd3ulVw4kvlwTImThZVQXWrjz/ssXSL5/UvG/tYbEq+Pjgue5kb3wOTNJ4nHAm2
x1cddxlaG81KOTKIXMBIVsg32EKcSZOjj8baLiucEFoq8tpJl83PVUErIXZ0TIO4YdOXA5dTz+f6
jNt4rbt5lGPkS1QIr6PwGIlQ205LiR4cRP9U953gd4kPrvssHGa4+3IMCdyArC6qzP0L7TfRPR2u
SALkdJu029m46yZ5LLFXhAqHpRuiw7KtWzIBP9MPu67wH+Uzxk1cNDp0YixkGSlUHatutKMIST41
Fa5MOzYiQivKmPImZdzY3TVJ8X6Hk14sJDzhxOPsCG/s0+Lg62kUMDatwYyq3XlQlg5FfFTVC5kr
bxMH/4uZRQVWv6aaxRrJTm49KsaA/aJa3a9oLm8/ED8gfxY7yHAVc8coM79B3KUHut8XGZgOpwUv
zNE7u0JOhkzLHFJ/bqMmLN5rg7FYXoPIdTtPQ4jfW+SGMK0T5vPcIXEObffOMmx1jUZ2m3tzyz7l
jfgoOfy/6LJeWji3J2uEGiUeALFoAZWEaEAvZJdii0PqDWT1n8s0HAN25d/NTvenl9UepvZzQ6O2
hW+x8L4tzDEueAF9yea2g2rcKs8FtAnG689Qrz+IfPM3a8V11J3GrMHVyOneWnb7gF7n26sccY3B
0r6raheFSpphGw1/se50+oRbBSb++M1nizj177in8/CRKmPyjtlbt1YsI82CcZlQBHIyDIXZ3JjN
uHXWBAbay1gdP4ryEFvp/gY4PVGXZpuUuZeiHyi+uOz/9TDFr6cqF1oBlQ/SGlMJfiXV+V2l69Hy
13N7eG7r4HXm100pn+ozLdUloZEd9wJ9zsYvuALO93/4fNG4z246f7fJ4h6dVg5J/EbRlC4eakb7
A22SrSlElmkW5EF1Y9OUYT2gt/se1iddmN5Qi0cwW2XTJgAyaDBr77dT0AoPcSvT2Fqv+m2XCMPG
XYfGxzDl0tA/Ket6MY6Pr7jTFiAzGtGOFX6w14MgZ4Sjqaz4uUssV2KaHN1yqTLGetppywOeBKI6
Y0bK+SSZrpriIAZaC+lQmOXYFImT0v/h/Oz9ji2wDy/4fWBgwhE5QD0WLEy07aUIYPhkGPUA4WsE
xuyDQ7zydphK3T2X8FJEOEaI0TZj9syZAYn6fqi2jK0qmQ0HCdcWzAYT4++mma0KqQ43N33camBH
wu7nUX0h8Jmq8LE/JkqwKe0dTm8pAe99zbef+7rUkc7Rdq4j93L/ypV3k1RL974K9ahEtvHeFYYG
459uikSgFpmNRvUmJy0gLJ1ehtqymBf5HcrkAeQxHmtGss4wJ+o871pbkXknPgl6JXqsITZWobxS
cryfMS+tsiKktzYfWAhYk/ioNMhpUaVJB7c1fRLHFHbjliMv3oq1TQ5VBxgeYECQi0ks8Qjv7dqQ
NR/F4Bkx8jmA2XtaBflIg7w3qlB265tiC4Fib8hD4rEbRi5yqIp+HTpnpPHvpwwzlAMgKdmCEvpp
knsR3qBjhFcUK7mWxg5nq2BGImkwGqB9VLj2KXNWgclJ4STdrfU8yeEp8hFTOjRiKxSqWY6wzMX8
qtOIdyIHUtbUB/INSSIKwceN2AeJ6Jz1ftCmdBu8gmVtFaZBqhtHeF74vT5jso0+DXLvvFJ5Coz0
nEmRaE/PlOcMlTz5TVGWylVi8jv3UyBwUUa3SFE+WWTRewr0N0sa6d2wawZWTx1nV+Nitz9hgz1u
wypIwCTGRK8gCdz4i5gSooirfMeuPRx/IQ/xMGYul3clYAx7cuaGSmrkmD5QrRtiArvqRzw63Cvc
yIap6rC37C55rCjSEVKUwlcpkQ0a4j5u93ruzHwvSMqizrEBrkScwMpVNccLJs1Sfp/LW7dsX567
5hOVD2BNACPh++UfycNO7oy/Y8CAgpFG3K4h3yuZG5nh19ZflIZ3qxhpXlC/Ms9SxSjH1gzUAANn
FXwoVbvoFEaRTGuUPbbqnntelqVShZS456s8jB1uQam/uAIQwhG9fHual80ObF3wgduBw7vnZ23s
M98kvUHqAKKH1SQb6du5z+vWWn/U1nPvGcSYGcGNW2U6VoNzgd2hpVSk94r6ZGfU38dmAFw6bvG/
ovokesecJBLztmM8gvpn1CM7UQhfab/VkP1D45/wdRkt34OI9wPfRwSue1v7erkaHskqLPdPjELG
SaRWIWLZStp7+0HpJFN94askpIRnC+d4/HJOQdgBmL8LYsdY+wJdazCZzyoJ/Kg4LLVJPyjxFAyX
cO3yeDtgNK/1WUi5GUuEA1fDnOV+VlG+6XziSlsmOqcKRe+eR7Z1fCY82KJjY1NCNb73Mjw4lqvy
lCf11AnRoxevvJCzC/ADP4JE2GR5RxEgA0ltHWPx1Y6zZiKRINQsyYhJTqstQRHKa+oukeezHtMT
vNU2gdhpSzZqIZKpMgCpXmpe0XJn2ImDLhdm7/qu2v2p9L2pp5WXcr0cUXM2FIuv4SdNvjhGQa3T
aood8tAhgtfI2xNF6fTDFri7Pdoqso91bHo4ZyPJz0TYYaKBdcQA/vBKKkRDxSfhMMA7RPgNsvVJ
fPMkSxj4X2mxXrjy3Rx3x9k52/kcv2BXPNIuGYgyTP7mIlviNS4PtXKjtXVqn9tVYU3ReE+z5SVR
Uj9SM1sNBYsyTOApfZbcWU89zTLZ0ibNKFVDwxKCxoYSepx1nHfPu7Noac+9LoYg887v8s7oTpxY
85G3K0ovDAqewe+EFL6OCU9MXh/GmuB3Js/LSxyh/f1K3yzI704j2cOH5NiE7NIo690hN700eeF5
gd/NbssmLcI67tvqBDxuWCubB9sh9GYsE0JrqKcOdKqbYEGkMQEImKTedNW1pz7/XdLt+tNjacZi
WD4KEYuJKgS0ek1uP0UuUt5OJAhHIilClFP6lVGrxCxZ5gGBry8eCf3trOmyXYEKROrSP57gy+5J
026C3d1WscO1bw0Erqgqdab0hg7Z+PpSe7uwAnbO6gqghRxyyB+P43z4tyzTSD3V4M4I9auSpVvJ
BV3Udv1YCXn8Npkj8ZckuIsIKmoql9/xNaXcf/UPlmCcAJ+2kLaiRS9pjdtAsex/Tnx7ay0Ar8eO
yztWliolJOmWp7niDfm4eVt08dqD9d87Hcx/jQygh2DZBCRVkLrPyogTiemMNHC16KzkZfn0S6WI
aeu9wWv33Xwc/eYDpqnLAuLJUIrstuilCofnZNcQePTwonaHjCep8RyuKgX37CRkE1GngFCqwSe0
z1vFfR4mw5/qEI9Jucdz+cSo8e5HfjobiomEGGwpAMAq6u51LTNeeq9jVsQ/O2XdLz/OfTS45Zj/
RaD7wp9Yem4rnx4yY41oAlDdbpB+HyksKcLU0rGN0IV7Z5LbBhy16oIqD0ga7ulp6smuoQoAQMC6
QfCmFu7UV1cHpRLaS5+Gi8EtfZRMnVl/sxv57y2BSGqJDwdNGs3OEy0UhpsOof1JQ5Y+uaw9yRMT
N3KVsu9YAUUeetfCrQIFEWuPjx0lgE02G4TWV4V4RdMIrv0UJs9t7ehuieOBZQWyS0k7GUW7j2ir
Ct8Kg6PJbWMZq/bbs/Mf/uqxikVDdB1tmPAlKvF2omjbKezF95S2ur/YhUF6ayIs/7afTLbDAweu
PavXOG0V8Dvxzj+y5OguEyiOCGpnkputKhKmxdn0t4lS6/xlAagyoSKxjAiiDGJKNmFOG14CgSZ9
2jX0Fhl5hvcJW4WLpemKV9zuJ9RlpPe85UmtyTrY3ePoBjeu14U6J7OTgNLlCsH5tcsk3JKXJ5KR
r77zm993r/qPrnHohxOITMfxHIdwF6p/7YIw+egpIT1QoDDPV0/7SyD0nP/TR9wS4gAZQqh1QCSx
mdCcLAWw7JrJOp7TssSNXID0Y9bOfjRXKTFlbJ9/7pBh7TdvBzfHaBO2HCg2R9qNp9f2AdEZ37Nu
O+lIRULwx++ttERAyKHXAneQ/ZV3Odfmno6y1WQkc+rpivGZT8InSdrUuSWyq5Fbp5e8SvWv+7dy
H1xNifI4lFnceG59h18e5XLKYZOvYHtLW+dyE0P/223GQ8mip7FMU/hTtlYBVehU6FLIPcjcZRbX
sdKvaPRKfMGrK8jn++VSF/JLTkHmLnfdGlzC/HVQqd9sZeqlgDp8rvS8rzLjg4pMU1zOiB4Ndgbz
6OE86sK+A93Sc/i+JN0QjojiIyDq027SwAJj1bjUnfAJeDq4nP9CDgDLmo5rojRVJA/Z3R9tYnW7
nKa8Xn5bW8YvjcrUHIwxmv5cBu83upR7msUY12NoNUo0/StQqBrUpUNYQJqenKZM8mLVqHOshhvN
8vuC8HFNLFidC1702vb7xE8SAzV8yXF/M4pWbvrQNIFBuyIKyauriZVMv7bOiw+rxLIk6Bt25/aY
QQDxHIMJSJHpB/AjzYe5SAbBLnuryyV1B5Pi5CQrqname14MTPlV5eHNLzWyAekt2wTK1rPztl7/
xX7SKgqssVvWyijiyQ2ITw5PI/oeOUrst3ASS5WIkqTxm3rtxLzqancLbjYm27PsVrtb+ZVhBjxS
yneMzzEyGqwa2GucJfA/QdMChLTek/l/gaonTTkqD1YfXa5mKVPgRP1A+WzO9LmhRINYy+r6C/d7
kbD3XFGtd4OH4WG4P1K0CUjuceFT3UNec+rXRBKYp42fYAf82Vn/cknRvZJSKRhEFff956E9I92y
sFl/PAX5knu5iWooVNj9udLmUzVo+bBJwkqptMptciCoMxqaJrN5g+xNRyPk1vCr9OahbMSqG76H
WPcPGKjzmMNNO3YoPDm0p9bnLzzfmImuBiVyIzypkOfUZNyyR8OqKTF+XRexCpH53W+kmVTMOrsy
f4AH3wqDPUjVGr15HB3MeR47YA5dP5G+eO9euMQXWo3UQc32+LhsqyBHF7mPDqJfcFEDqhmfugfu
lgyVh4XVMh2hlgzZsRT7P/lgp4P8kDhvtye5iwr6V3R5R+rzcH2utU+R1mwcEb2ezlJH4fEVmCim
yG8YhCnpbvWM3EVltHJUA+BszgN0hQRV0boMTw5363flnclHFe3VhYg8AXwoSnnzEfH6jHpXME+z
QDsbFeXOCMgxsRQDySNx8sP1ft/DSMaF3ozYhb4LfAoKuSX+IkRM241uhXb6Wy6Dcuw3owleVnS1
9pml97T1eC57Pu9pco0nyXxuZfnBwOvCBA1yRUdyh9KGpehl7eZpj9I/Wdx6ravIzCdkyr+yFbej
iKXH2zXXcFU0NjWv6ROKMW/6HzOLwflyHIBv7awWitpx5+EJjANi+DLiQurfH9FwlagZ6Whu7fm2
i/E1ffrEdjQIsdJrqPoJTABoLmM29puPh37DPWD0EudsoNGTxBXn8w5v+y+93UXi01nO8J77mC/d
IKYH9FOCgNmxmdn7f3DdLASNu2PRTyENmn66v1ETxUAIYlLEubRMOWengC2IV85RWxkGD63/9aCZ
8nEEOFfu3yWxttWRwEvLW7mmnWxqFV38gKnma9iAZ9+2szkmvL2iGa7OlctiutJrBer8H24YI/ST
PlLosHaQmINEqXRvpaU+03N3pTu8D/SitcevpklhkKMdiPPppD/NqilwB/1MtcR9Q62klFDMWdbC
Lp7/W41sr2AEUSSLjzeOhgWwl67Nm9fmUHD5TP19UORpJJMbK0/iz2QxH9S6uGgeegWmOP5601jT
6H02S0/YQVtc/QQ34L7m6sqK3kYBECT/6VyONuLNbcQbisM3zkAXaL18N6OUqlTUxhLQmWWCyizR
MwMPZlhJrgSv3xLvTjwBjM9xivzuYy+aV+f3IJ5ux6IJpXAEa7iwCyxxXaP1gr3WOU4BMHg5dukU
ulbgy5oGzft6Mledh6JhOZE9dNdpC2bjn/roP4mSPJ/OewMVQCreeZM6oQuGg4pPXShIrw0xwBAu
ibY/BQIDxYK2qB/54xyO5XBZwSMvS37BIDlBvW7PVroGtXbAdJ75YtfvNkf1UgUBKcvNpd+58Huu
/6jPyEFtR8x3tzK7IVRoKrT3Sxd/0md7zBRD8XtWrz8SezdmNwW3Q2h+zQ8/Y1LQ6kPX4Pqf6h0W
ZVylXvAsRWSnYEK1gcEaYLBcgGOriEbda0xjibSU6+IsUVgcxSFZ5c/aB7646NaUN+BcAYrHHzo8
3xVxXzijgoIkNf8H00zSS5AtVdkIPbX9eE2D5zGWk0rwkrFMxs2t2L2aw0HYLu2SoI0XWp88Mr7h
y9Cj5Q2W1lJ8SgpD1fN+zqJ9kdqwtQqW5JWNtbHNEHSn+woZiX1UmTZ7J7eT4L+uZRXlJfTq2vQ3
ThUIB7hsdNGaoi1ERLvfHkoqYyu+IrlPPsuybTBagOpikQ36KEO06Jue5+g4vU2wXKhV0KVvgx9E
tAEeFp0oGEpvB476Tyev/9NnuDOKWmem0xHbqJhc2JPFDcaC7y+CcokZU7T/2a7M3S3785FJ+3/z
pUbgDZEoRoNQ58fMqfFlnuVanQBhjIxvnpwqJc3lBdsqMEB3kKiQ7eoIllM5bso8asmQG1mosU6e
uH2L4BMjOeGApE9WIcp73rjm3ivW4QfYPEymU+3eGIB4CaiXqGIZFMWojMP0ckGQzmCwOsufOUr8
ywNSGBw847OY25gcXdJfY2w7FHjew+KrtNblUd8tiQAXj/0JvzB16GwlKVILDF2eIC2zWqkviOtW
aGFcctfg962Y6Lrm+MFKwMyjAxJ1iGGHsXJKoHGduXLkkLAfiYZMjkN95IV3mBuMNiY4RK350DJy
LrEOqFNBsuxqPeIFCE4li0vXkNfwQebN5geqkbeAJFdvK+6wmIoOA+lMRKwut3y0yFUzDjsP37qS
Pjus1JEFXhEp91UVU1iXE+SF7GAsr9RoWc8Z9IzzvCzlIWRf2qaS9KnqZeI3xWNoP05hHDtMIsNc
E2VXginDNYWIHOr0QsR4nWIMyzvtwmKDLQFkq1tvoJAnyshTfKH3OzkTRIGpsqC30M2Y/D47jEs2
IT98KnMq3La28PV5aNFxm98DDCufJGJMJIB6zKeMeSx1uYB4k98LhpuEYJqTQb1e16/DQ4UWI7Ty
EdVSn2rbUVuriG+iDHxoAOPgxk7OgPxoYUuI6U6MARxyMxIMpmmDW8wPjWJzbW4eNAETsPkyEwXc
SByb7g9d1kvi5Bu9vh2LNgvqQ/c8pmHj35BC96DE1QQGEeAVvwrSbIMx0sOcWnpsD4Y9bkPM3vRQ
1jEWAJPihJWEWPbsceCUJwTj9f/WYffyQbm85C2ueQwwF+YQ6t29g4bW6FThUcfelq3ZgN1TnF19
Q27WllZdOTHJ/gBBu/lLs8sSVH1TtxxuEM9wBOYc4SDFCRpT1bgd9bA5+KgHXsMRYa+Cykt+lIBB
qsyKpFNU2+NIJJOxblY5Eue/Orl3bfk3DDxC4EGeKznVKIACdJhKBu7VNg1NmooSoYInFxeuO0lB
3X4mnzmvNVgXupRXrU44kACZqWSaVT4eUYMGjQ/1N86TbXljL1bdTkPKoEr7VTUbyJmYF+nIQvcO
1gIa3UiOjHAK79163cRWz7G9fFJHXOq7fUBhi76YeH6W3eQw+ujHL3OD38DaKd8w1BqT39W++Fy4
xZ3s/A9B2DQwNelqXQqkPqVRkLCS7583sBz5bqe1Mhgj44NN7uREkzCZw1GcdsdoUl0PkaTQeEA2
6E6wiEeRIzRRBnL9vgpdMkIDXFbdSmketu3/1/mCPcfNG9YsAGE4U56eEmWvITsUkS8aMrh4ZRC2
CmwKrSDmH9KeMpypbsIYoIK9AUguy/W4oMQOoYzZrXn8w8rJtRRBujnjAGkJ6MfWUrc47tLfQOBa
cFqsJcgL8uW0AEspQZZsAsV3tCXaDbSFPDD4XqrTY3hPbc9XQWgOcgSs5M9prex3hg3pLjOarOcP
IadiMcGteCgaJK34idQ9HxuTIDeV3mFPMxrB/D0JIWaVSJPyCQmTcD1V0ZhDJri0WwUX1UxS4mmP
W8RY4Cq68h2Od5fB4ejRSnEk/Z3f3SHEo9DYT9OUwwxbkO7icD1PBi+OhP6tpj0fD2Fzzx3zP5Ae
znHaeRTwaQjk0rb+TL9eEQ2f9ik7p52M1AryN0YtfbuqxSJGH49Hp9BIuP6zties2g8PqDAdTc3k
4tqvE8cMV2m3kEg1Kyg40/SZbdThv6kRdjuR2CtjGDF8uHGKqmPbFHkdOJM0/C+QJ4b3TwYFlOkl
3KCDaUwaCMR6HHEhGcO2g40j+lxGnkHREBQgT7/3coIrnje/g2nYBEHl/Zq/zAvS4pmxQLJnSgSG
ZRZtxeXwLCffW7y7mQpEXGCSzkkRdNEcyFZMns5WFd13Jsh2cmjlabAB44R+CmF8oAMzmNSCDQQx
pwccxgLoKzGcfaLJ+YRo3G1o8CMzlsBpAX5yMLX+WBSbUPbC1BfH3vJGpULOBc5YcnXOgU/VuDCm
nrRAGU5pdyyRjUOX4n6mXuAiLGQw1K03awkRGNDMsn4XE8tRuggJS+dYyh3byuz3NWuCSeD7tAt7
JCZ7HstLoW7T5Zxy42Z0R+c7HLumVyGqCGZDBCStIwRhA/Op9eEzsYJr2RaarKlX4CiIW2X9cDHG
I2wKF//32B/9ipWLNyopqZaDCd0eI4YwJjYode7PeJJjunWBwcsVSdSzSfGu95SrU8GHy5wbpurN
R48JQ2acYFoIhSNOwhdLOpIrN131ytpK7sCfdtFFQkNfpbyeUumxW4ULDuPLN5fkgQ6QDq2TIoUF
vzeHJRZVLiBV2Oj9rTYpHd1Od8+NYg9FkBnxLiXbgjir6OB88h8udLsKb9D/ijYWFyXR3tNRJcN1
pc3UlViTSdqedpj4CJUi+jI5keAINVg6ps0Xruy8zqZtPbtwqpPLmMQc79fEG4gdCpDK4ZXHNCfj
ulDq4KDVBTmsAHyoFJYqjEkkMCxXQ5cUonSdZlloanZugR9IHDQ/hVFEWxUE06noTpppFZ78+LKW
mK3q/oKbYUL3j81WFnC9ix8gdquTgaegK8rJqIDSSOVyKI0tXIdmUMtkfrI9DIJsQv022vq/mrHM
AXS4ehT4h5Rzb4I6lzs2UBm6AxjT/zpJniTIpK61vTXtrO8KVvkIyIw4UqrX3YH6sk4jMp0NFvsJ
h9e4Ksx2mrjtk5/OTPQJThpOhkQwW6I4VTPMwU2seOuujJvFcEnwC0g/ecEFcSSvF7Q5CD8mAFDj
hXLWyrdLuGGTC+B2aG7kPJdvGdxWYGpuhDSntlo1x44wd9BVKKfYMHJnUjMUfojzyUVjQn/TyVpI
P3db8a8z3nsBNS+d/idjSdS8LUKjugWKv7yko4BEauncNlcr2I2YCl9YWDBT5G6iqV4MlHUviuRV
Q1jkZdfcgohUGGEnqNx9cqswUaYjsfKPH8LN6MT0bdTxRvKh/Jauo+yJEGxfnXhO4MzAujbP8RlG
SPCzFIZydLlvxyM746YBowjctAI8G8F7qjZPzlgYqOzYrOIm96x3tkp62VDPglmWKzUs8JNq/l73
RZXQFC9hN91ZxPr375PbclprM3n1zugshRB54V+43AXoAKXIE/CP5JLUuRGu4M9CiXQubp9Z0F+8
XFeQqdG1jRlK4jNqiT9VpJTa0s52Zcus8cFfbJh0l2qVAL2TKWNF8W+UfrvOamHjd/0zsWsLXThW
jh7ZuMNpNPP4B+pUBmYdDx3hX9ppzF+mjQS3nHd6JisyswURRKz6OoeVVdvawz3+wrB/vkPjPX35
S9u16z/o70ibsq9cm7mlIdza5GO8Hf+oQqxfRAYvgZH81+AjalZGFGEGDb7RSLN17J8+5efkfOU5
vAJraWYgoPKhjepa4YU3HKUNLwbZAZ0TqnnxB30cej8aTg1lT/UZQo/pS82KJiSxqiXpGbTMCJAR
ZQkBaFKDe3lK8jHFp6ey4bzFoppWe9YgsASesfiTaWrsnTEEuC7l4GuMPNMAzeF+87xlfsb4U8Lf
MJrSUtH6TNyBrzw8I6pNMYTif8jHUPSQAmFzvtarMcJ79NyMzFKKZq6Mdig1O/MnLahUUvrj+5S6
HyW3xEGdf6adqtVKdKnU1TbWmoLkTn/kRH3FRzLyCug9U7kJCgmAatmDply0eS1O/PBXPXSINdYe
/deKJzuixbyqiOKK1fc8XLkpmpQ+1FqSxzMF2o3Lj+SwQiTI8KvTf4MBa473Gkxv6XwuhW66EY5c
lRXuwCeGcOSsUzv5VB4g0di2NbF8pLu4n8WnMZsQYIzyduZLNdvp4N1yPsoqRzXdHANoDqeAFZpx
7CJUGKPmboZNnmiV5n93NB3XNcYlecZoMwGN7PSY5KDl/RognWkHSpdJJmDc/mnvkTFU2uYI9ZSi
zCdbt7PKApQI/geM69rAKTTlH9P9CrDGPsTO2Rg1h2T3Y4RZJg/gnXohKe0ZkcVZC1My3Ex4o9/f
5k5rDWW7UkSKeTMvxt/xn6+55oeprYPTxUyGu5PpZU+qHlvFOhRNWCk7gftPz+JlmFW1FH1hVV0P
FRp13mOk5GBcjU3LubCmeMC2Nd2q+1gf0hlNvgzlfDS9eJCZgXa4I/cgOjSu0bI4sX2NyhaCq48C
yrQFj1wfnLDB9/iLO11dmkhMHbpQeQM900+yYKTMulIAutPfo9sPWh43XqsofUVrVWn9GzKEuwHl
W+jfsOArBXXvITulav+LkTLGCaWvq/a7YZSZMfNs6DXQlVrIxLUvL5UkJQxeMjEu2cLmdHYzm8nt
rVaQaih42OR2ccmp1TvCkRhoYrd6zPmVOiIe5QFB+8U1XooduiL04750NECQE26w3P9jU8dVvTpq
PNUtFVqHeC3GU5BorXaC4u3QC4Z0pR/AcsbRPIK6drALOpYBuC8ErHl+QXb+WAhbMcxl+7Vc6p6R
hGZTrIeT6IhdL6f3Lf3rVlcWFrrDCaCBjVOXDXDgmEiDf6LPEctGkk3rcg2nMW3LMuEb4ZL9Qyk6
c+oXq5s7hqEOAL/iZvwVAg2smRMk/xk1dyvWMQHYJhk2A2qtIQDP7d/dtY0Fk/CTOGo2/p5DhjHQ
wyGoevq3Lck/4y+9y3rY4K/O90/PHOGG7gOGKKP/bEk+nkUwOL20vUrio/fyi+8/zLf7UZJU2MqA
p5qLRTI0bGEuh/BIqwvyAnpswJfR/kwl4WvGkjxG99MCMsi9hgy05hT/VFkk2lN/iss1+vp7QBpg
t+/LU2a5B8CYbEezw4IncLTTcM3SH2mIAjzcVFimKo7+RjMa43dS5no0LlffrTj3d7PLhH5oEquX
dm8A23eD3mUMFvcyF53CUlezhf7xgupx7O19CeZqyG7BYHe4IpcxNUjywEHFjs0jWI4DhC5ltRMp
8ZuccQwkzbfYdp9hQn3rGyxdOfhUyPxuY/pyodKpFuRYw5ny3lUIMziUoPq8OkTq9AKGclOwW6+5
dqhhzVkaJwTrdU61c5BLtMgMVgMVj/5gcinQalu78kgrsUtOwyDpJC1I/P+hz7eTzmmTQyZclwmg
PLeFgcSlHFjZwAJI+AMINATdiCN0+97o55Pu4QbIn+TnxLgAFJBbHKEsBq3s546C25NBsFtehP5t
x+qRdZtOrXYXm7XR+9YKRI+iZbintIGkgPwzyG5NjB9UT0d1mJO2JGEf7A4xkwwfWLUjPu2ue2HJ
IrwpN/nrgk7kYt8slDmjiFAtYqEnf3hnY5jKGxHceWBne3cHAPzUE6I4YIaRzG8dkSeyxbuI0j6T
63vlIUqhVHDjVOMdKvwyla9ccS1oHopUOegLsSDrbG6lhNv+ysBqeBqim/AfiHhXZKA2FWZDm6D2
HN5ZBeY83H6M9XuoddJ2u7Zn22XoBAZDvNLCRvca79xY12QikkVzmmPxRLq8ScSXRkAcaGWNagx4
evjejbD93GOVPrQyC+HTir247qaRrpLw0nuWfCpHv5KE0Zbe9G0Hi5w1fsrVw6rZcqXMHEi3IZ03
dm8PsaV2zqLoI/XoL1JQbhnnKDB2EeFsgoDJGH21IQfGZRsODelw0qvy1IdNYRgUHx5eDEfMQZwM
m2/vxwgpaJUpVogd58Ntdt6aV9+fBT2DxEEVJAsUw60aRKXrFUlt7XGl8ZKCCX3ou75MfE4jvfw+
feZK70TtvwmRaOiLHUFpkkfFDFeewzzmXteYPZ9UybejxgsRp4S58C9oTTG12bLcmiqStOWPrvdT
I1/4H8RSgRXpXOzlWNbP9rcCercXMDeCJob/BSCvfP0NuPc9z/go3cT3Bp/8jdn92lf2SqUv8OL7
fSdoUZ+IY/J3Fsw/vtdO0KXhm/ut118GXDx/fxSibQhEgw6w7pyp55lmliN88kbairL1ML5w/LLY
juuG/5itksowHU0V1uPvtF1F7CXmKyKCrlPHvEKraeUVjWcVmw0KX5GNSxNLg4w0ezW4jzXs9ySl
XMn76xKq8LbShqDdoZp9dhpccK+76HJe1G1KQoYX97IWm9q1ty1BXrofnz27oEqzcYxf9gtf/aer
KdTsMiuXlxWayoBjPLWG3H/mMk6G04oLv7hPKw8E+26WRZwOX07OPl17aJnR1kF9H/q6K0Ru9Vdz
OuSNo+axaVRMOc/IwV8ykl+7IIhlSr3Xa5wU3OhbQFDMWQJhJ7jnOs/temb1cqdz31n+AnOWvC63
VC4nPIa4U1Nr7fbTH6/sZPRVvrMUYIRn0UUDKP59Lj/opfLHNbZie7QLqYEG+/Jv7VD4RmkowsXc
maQvDUv1MO7juRE8vS/9XtuJqpcnOMH7R5Ld6jCdsqnyNnyZgnArNhVAAoSpZxMFUiOckMjdbHJR
nOyGFZAjFdNkT9HtH7zh3nJ8m4H6DcwAcWe690ane2Q7ZJl+RjAREbBKdFO7fWF/HYagJAOT0ntk
BQJh/XDSSXCbYZD2j8kzUQC2UBqfyVimOLTQeqOrn5H1pRUNI5ObfyUsmiGm7i4grJMs8+KQt6N0
Q9ENG3BBCINsZYBGnnf4UaHtCMGiZ4oMUKbu1cVDjUQ7VF7dHMUYELW32V3CwdzyEC3hzNGePcLs
BlsFyrcHhCsSHrlKqQdNQTsJ08CV7nEAY1hvmUfCpCZeLnVx8f87HLuUiEz1hlmpfleo4ipAXn+W
eTsQsg7yHFeZAWfYrZYeg7rmFihrHGXJjDMp2usSZ5+qQuKBT814mbNUEejY9GoJExUqbD+0Giia
PSV7pVkCnHCTI6Qg4wL185I6ksxYKaWbmCUlBYaqdXt6e65723Il0qc1IWuYc7FqaaYl+SCYTTp8
sR6zoqaZscrLAYirZtZdTqRHsPZUd0xiNvce/yhkEeuSetcgn1nfAO6Xivzx12+K1ezLj/SOX64l
/BX5iRX/pZ7uhU2laqtOwyNMYwwXB46QfH9ObmBCRRDahUTa2dRPYQRy99PsXawAiDcrqX74NZ0z
f0qEqDLrC0Xze4iusDsFnwjvHnEkByLHhqDWx6H7ToYnlltHuJY6DC6Dhn1cauEGfhpQE9Z+31NV
8MhlnvR1CZxplx6OK62nVG/Z6Ggv3263W82ooMpNoenNE/IrrqHYduAIz8dvGfBr066QXTIYL4KM
ney/7ttKYeT55GeB9u29iNqXkip3jYqHUnIbFyVCh1+mGUGlnuaFQ+pKLJh4q6p3g7hhS5SNZl+G
sZtgnpkkz9Ek4uM0LiFlCCR8FPUgek8uoyMO7pS+P96FIQvmuNElB4eV1ved2yQxskV5e3PmtzH6
Xw9oR63JmPJW2kznThrjZoA3z4PBvyg8nrgvu9JPNRVenzBwmVSxeAKfGbjZ1JG+j/VJWXCCeWnD
aVkO9pl7k9ph27k8HMII5yWVDv54DIk9QHjf8pqNEmKqPJ8TwlIMP0u+Eykh0TdSkwwnGRkpGV6V
yG5IY3/0p0DMzfNViPrpbQLzjgmFWSi/bQh+KhmS2SIWXHkAWRUocIwuJZGAZGo6BLNoyLHxl+qG
YrRxRP+oHEsMbzuuGBttZwvOAbtNq71+n5OTxJw7qiO8xo0NOtpY+1ySNjeB8edk0eUucji1zNxM
vCNmz8ZLxvyn0sAtj/tingmis0zoPUJS+fZG0CMIbVIMUCs+uEkFLhib1nwRmcoPLy3F/eI7zzOQ
FcJGbgMrVVm9xjvy5o2rSrCLTJGS1yW55K9ghpdcrHK/HeGa5dNpv95xijatywUsACm2eXGGEhQw
BDw0ptLIpPyHq2+Jq3E+GHF1Sx6CKjwApQQOb6Bb/+cs/CLhQRHsyrrb0Lwh/BSVTwgdJBrge55Y
h+V2Joi3vACaLbyPUQAJ2NxTltueAHLuHW2ivP6NJxIXgyBWqUpLt2K40+584lhlGgKtNwYU2cWq
ZUYkCkWflEXXP0V0v6ZV1utjKsDGV49CEQCukvBn1CnLRQ3prLYv/06uz21K0/Fy72tPWzhKwrXe
jSM5pwp52iL5xsP1vR/9ztipAavrIZ2GKw2OszLgQzYIOqnm9y/0+B3Ax/K/dWNWlx0cReLqyYsG
hG22mSleEfTVT08k0/dDTTkRSs8ikCjODf8jotrkWVcCTw4rCdfP4m1Xz0h+cG40d0zykctkaTU+
rLDCCX9HbamnqWCqBoDdWgJ+TEnGvKrf9DRSlKYremKH68fkvGDz57cn/jBo3I9J3XhknHRGEScw
0Cp7g2nv5csf499g0xmjvvZu82a4oe/1SM5Bb3+KObFkenleT84mdwZ/qZU9/qmRaNuqFQoSYdP7
kGHulT+iYppahKodZfA6KyaLwrGEmYh+xeiGgSzD8q99q3WfNWRRaxnY1coZvnQVFcVQAMuoxDnn
jpIhDi78WfjlMS7h1jIw+hT70OvfkHuIPLwposnWniNdqdvpA87fwCj3PtF21Tt4nrCkwkvMP5QT
szInRfbbYJHrD1gEiLMw5VQ2Ia63nDNkKFqFH3WqprgtNrRZZ6WyFBMv5a1RnWcS3Wg+YOK5vWR3
wA+F4erEjtUtMncOCdnwSWpw0XY8dkaLSG8k4bl3BYDThh9q0LHXKHVfjEG2y4+EWeOEKiH8ND6M
+4OAKW2LQtGmsKhcWkZ3yBHaoPZZYenGtP+mO/M7e0SmMgq2S0SYsuvhg95RpbRAz6G8tmgN+OVN
+0bnFE4eDUJHepb6/IaZQgzvumCKhSXaeKN7PoIrHqB+U9sGpQqrETKMrPghMSPfa4O2oT2KaFG6
QawZ5DLlQHmBPSEpzKPqd1e0/+OP6rYahlUERPj4NlLtx77BV3xOxsXQpl1fANsLuMLh9auaKma1
L7Q0l9YuxkaOw/GgdZsJxszf9ioQdgiM/lbURgAdc3u+UPWbuMM72UG03P+h33XancvFraKdOC1G
qE6sqO21hBxMGVoQIGQ6OviLjTmkYyhrNuwwXZedceL0jcOyRrZXtBn6myX2H3WjPg0/fIhOZQC5
HfOVdY5h5oH9MVtLZ+ELPnm81nqsiHEYVeRctmDIyaA5szpw9R7PEtzSNgsU05E+lxzMGvYcEAGa
ID6s+bndqhE/Oxwf4pn7vAvUf3ED3HBsryL06dzFDplGgOgFvRAfvlPip1dPXDwQMZ2d3JqLJAkq
lhloNojgURp+4Pzaq92WdVzWXEZmOvNqkmh9ArOvR8dIiMs6Y1sqKS8gHRCIYMydTA8kv6QWOG8P
jCP4mi9XqJM9plfv/aP7Qri5QLav+Keew4YWfWoKkQlvUt2ObdNmVQUbBxYNseEXglDwjReqoK5Q
j2lIDqk25UidKAhbM0KgpD9wfYymtPcVjT9DLNP8ILtJCGyh/UlLBvi5Y1FLy4Vv/9za30xbjDjE
ACpxS0THPQayKEpxq1Ls2GdfLM2/HKEQl8gyBKMhCv0PpWwpuX99HbMAmrGmMawWPFtdTAB3oEPo
mA7smAqcODVoKhqVFfawAYJL/NFgI1VI+ORBV5PlTMHkLkxrCgbUb7rvfFCZrj3FXDpb7ig3YGPr
UqsIqaxrVm2uX+sHjWjIIAoEp9lvSBltmoV364qxC0p+jIzmtPYPqjA72n9Y9KosY/DYaeox1RYz
HOlDPA+IOrAansp4Mz1jQEqJgKRxrR6PVDggpaXYwyP6MWlrZDtnzYf7c0Yx2y1EKoBq9V+W/mdP
AbST1T/opDh1fkxyzHMwvA0zt+cua6xTpiBMJX7wAPiuWg/cdDuOP5dX2Xk503p+bMRl5gQTdZdM
0kcMySV68nv8I9IOQUIY9D2fa5S53F6/ohhvnrLYWp0d3hzQGAoC6QrAuV6wDC56T2RLliJ1EPev
L9II/+JBXd/ioWKki8GB2hVGSVl6zaatve1BflJgj+SB1vaQE8XT+Cb54W9Ny6riZ4F9fOhaM8Eo
JpmrcS7HtZzSgppqyKCMx63Aaat5CFwLtqquy1+BIEGXXpGHiZ0tn8Qy46N6T4ebaM7GGYCToSIW
vv5q+6xTkyazhHr1xpm0LeV8wRvo7ZpfM/heMnEiz1ZcetgugxhyMn5v8QOMQkPea5HgQeD4zLHw
psysMZ931tV2pfB69FladNqecSrsUnQEF5j9JZ/a2KxmO1/Ann/nA3PF3C/6v6FeNVHesvQQhfGm
gPOpYXy7zxaNw7fayR2voIyH+fWdF4SNR/Pta1fZUYEBTFYsMz1959QiChCCfi/QVF3DEJHEz7z5
NHg+yF4Yufs1GcStAZsbPTACRR/SRzBWK8G8WYEfK063+cH+ighU+qvictXCPXdPcSsR4pxBvd+E
oJGvzUoZ2QAp4sICUQKUTnndnY6YBrzwOsG6bp3QRv0oBYVR8UpsVUa3ZjVSvGVRmFnw8sCzXHro
J5VsXWFy9SH9nomThFPUX1wSovXyKy6Q7UBzqaTbQVIPWIhZDndlBPHUbwfOze6yjt2SFcOzST0O
4DGvwUZSwWlDUELQynlT0O6lATrA9mGglA+zWQF0KB3UhHJWsPJL5Tunea+n3Bg9kmFbu0PdvyEc
BqaQge72KASfKcZyTuV1er10pe18Y2qMH7DeQW1OlX7n3LSpjjNnUKAtaZa7fKDjNUYWnOK7+6zm
KaZfszBI4KSI0dFo3Zpz6gJTfUmOuaK9qCliLQjqhamqhu+q4QhU0sS8Kh/EAfCgzrIcAWjVT6vf
i3H31uajlbsmdbMNkr/C+eYz9XEa2CK09Hnj9rC15LUq818PA/sdeVLu+HEWHHn3aYiERk5Ng7xm
aftZNvzoYo283wXMhDHItAufyblI9whUbGCvYi+p9NeZ7g7xWI2fFSIlYzOd+UhkzgFp6RTl9Vyc
tzuCQ2gudXpY3nMdLeopTwGJR2ldCHbBHGtFzFMhGXwaEW74xlljIyPMG40lHTKtVzqXD22kYtJZ
JUdwbnN6g3s243hNRl1MjHtFkNQCXm7GhBDLWQ1+dKxpxrQNMpY4Ur/7GG4yqunzNDSyl/3MufwM
mKCupyc6SVvhAk/PrbJSBYXpQY5U/OnSUobjk7Y9fyRPBWKuJ+hbftruAkzC1dn1tTbmK14Te3dU
Qd2Divtsn5eX7cnt/hqP3ImXsMHfxdJVQhoouFJpVbfj1Pk4+Kva5p/j0pQvjIu7yGeJ3KS9mWrg
+oGD4XW+gOo13Z8ZjL5ju01EN5+fCabDhinZ/jgdn9cFZLk0bsGAjLJ3OIBWCl2YJwkdUiHth8cr
Gjz48BpXjjDLFKzrQmbld6EGB8jtwgJtQ3DZ3cA2pqYe5FN48C8PwN8dNyyzaa/8QGm9+NkCxUcv
ErK82e14byd6c2HUy8z8BqG+0wsUvUdbbgnv0Mt3DxenODBInBX2OQIN6Vzv+WeBHtLdYmkJ5Pk0
qsHsBRp9YeIc9CugUMm2RCy2yOtxyZs40eZ1uwG42/vULdI9q5dKuuJAJE3Hjnj4yMrMABkjfDGe
LVkDAc1r4+YgF8Exb4NVNWtxOdEC+3WIyDpegZa67maVtXj7sgCNjAevpmyJ7f7vuFTMS+SBKuPc
zroFyBx7qcMgdJaWg3gL0AbXr2cFJYi6Mu2igpNWlmQ7dpJNSieRYvMEVz67mqa5RIpoh/Zw55/C
SGbWgsm1WkKxgOkXmIrXbY8Oow05Zwtz11QtH/MdJ3rleDaARv37VdlHQMzGuj1FNwXDc4VVmj/Y
QNdrLgvyDOzeP4nO2UiNae5qUMs7NQ1nqQzUrK3xrGcsnWb5tMJtBWfWCsZ4T/yYXY5myaOq2Bgo
QXqpzAKxvGZ4ElEClfj/60rDJSTFaP10rpg2Z5hrogLhsf0FICnteVqM88ktsf0k3FNcEyyjzeGP
gTr+ZGt+NegMklGC0EQo5qKDQb07AVidXlEqHeNc6VgT+NwnIdj78Gic2OZQQamzxuh3dAvoXHIz
+JgVSUkKW6bYAHs3KVW7CQN6rpF+9VC7ke+SkfuAXFiumwYgWgQjWyC69gS1uOVJSPZnJtV6qqWl
0/UX0MFlz2zU+1qimBEONksWHZNlGZOrIJRneTNbhfgSX1v+TYzVg8QQOQpza+nhAeaEdUDrq+Fu
9Rz594MlW7In069NvkB7xInZ/5jtmSLAyYzY/Iimg6qsWLykBPPrZRBEgb50rIjBwTY7xw7T9Hv0
1QkyoAw8U++viiCebbCiwVwiAag+k0E35/95l+ew6wox9T+d9CYvJwToxMfLGosdAc3YL4GiifIn
ZfUKG8pS/voT+Dg9sd/J8IkMHUcsmaDx+z0Fou0I9d6BCZ+u2M3xdkuElDC4pNvCoCWBvL+JoDmH
wz0x9CALHHbPUBXCOuoBvLzjvj3Oxuxx/oFAFP1Iz8nEaZd+e+d5lGLNYsxWgz+619y6GdvPJS7M
mdglcCiKi8desOhljPxS0yqhgYAWpeuVQpTnOPrFGD9ROekxIGUGe7Gt9rUfHqXGy1NtdOsJ6cPW
p0ln4t3npmWvcwpGAyrikJcngcnue/SS1SZeYN5SNDhjJyCzsAjIt5kPaC6oRTpqQwmX+ek5GguX
ZpLnzj6pLT9/uyOLZ6RRZoMaRhJ7FB4eHBytvy7LYlz51PXsvP3XCfOMc6GKE0shet2Dc4g9K6wV
rJsR4Ty2Csscolqwd2QpByXV6nevT25E4lBMc+jOkt6gxu1HPmKNIV/74bLXv1i5llZUbRE0uiU0
gqFcxHelTH03O3opNsI9zSZFVfsAzpwU9GlTFgDi9Sg/WA3XuEqdSgsimaUs3fL4hyGX79kTvXF1
84du0VPQEkbbflRmJwzguJ5MNwtXMCFW3DiQIEpSdPRzn8PNF9XXwGdyV6hNC9KTZKYkmekk3e8V
LPxBbbCl9VAce3LAJB2ZC+dJqLRBlL265sXnfynrmQkNwaZxcvHyCE+/94kXwuMaf5DG9STmZbRo
YV5YUnveb2hHbVLxRnK6IZnv+JHk0BY9Sz0gEnhRuZwOZQeniYOqKa354galh2gJHSVrBweStge0
aEBRw+2x2P9pmceZnoHTvPmJmOl8oX8gQZuWoVTYj9SoKPwkTJdtxCuTpWn6KFUCyN9YBdM9gna9
S3bkoubPpww0GjKSt1hJ/yM7se05h27ZUa+DsPGXh65rCXMAXnzE5SD7F5kiC8MlaOqZ1XeJku+n
aVl+wldtAPuKTn+z4vj3RYUwH3Fv3yHCSTg28COQPB8m080g7T1U0Ygw4wC5DcgN8p4wN83KnPJC
JXQJPz3boSqxg9XXKtLR88VSxeIGB07xWyK9OzulxEcqt2o3RrVrw9N+FeHF9eql601Ihin5yKAe
EgiJHudhy4wEWMgLACjFPz42lWx0DRVjHNJfzOyhs/3uDGzJdGbDWAA6CUk4bAdRBAxDI1YaaHR5
RrJMjYZJ7kj153L5icZ9I4ayKphFo5lpJnc3mDDUSH+xpt++W8Y00qOT7/aYFw+Djar8He5a5ZRp
Cmo7ToCV0UFun7NPVFo/f7tQU8RbEu7cW5By6EtTHD52KOpKQyvR9mIj/GF+RsII22o+r/zmkoPz
kg+TvIej3DM/2KPhoUz+F2AC/Y7wugw4FTo4115iBtYc1dow/mMEtXn6rHYIp2MzOr3A/AnTBuZE
rtIGretaPB1ppdZNHBl4TQOedG9b1s4xtQW7V102iKFU7s7kMqI97QrzhhL1a17mIUC4i0ee4vvk
4s9zRUHKy7LTZ90Rp41C9aWa4FzzJdrvZkLBxxm53IsGLrif70SukT27NBo442YZ7ecwYLkRJT9v
3paj25qxtEY/iOR2gWI/WNNfohqrsAp3ppXrNTh3g2YaKC4EBWPg7JGvkET+zGbJfCL9cpV3qUaN
VyD4IvdoBQ9LxUbtdkH3u00gF19ehb7U+eI6LgkjTtH/qhPNRU9MGXdCve6g/3GMNpWwRr0BnZKn
YXkkrzjKhA7ag/lBOoSqTkAZqFigU5UBpiLKyOLjHxUzvKDLqfoNzUybrDVzy+NAiuvpDUArMTVV
VfdbqLQ52sXlDAvr181QLrvj8QBdS3GiOQhFlfjZhMypu6oXiKb5nnD8dA0uZnuhDw20bD+jQ4Py
IFIBoz3QtsRmbwbB8lnQ3aU1/3PL2ufZFvRmWKfeZQe5s0zUsVNFGLj/QpsMueeIPYkgxL6+o2dS
9PpkA4ih+XOGIGi2+EamlBdcx70J17fhZarobDTLvVBkkyAfFzVCIbLDlRgi6u6X5sP3TnkAgfH/
V0bqZpxbnuONX0ctzS6v8DStuQLl8wq3e/CXPweCsHbSxAQez4YVcenBuF3kf9EQfFf6iFfmi78w
Ir51+v2gXKGSp2zyBcJv6GeOJiSE0rLvb+4ZJAmYoe9mrAbizVIWIdZb82m8Brf6379+7FmLvjrF
odLljMYz+XoxF8gnvE6MITkNhgpmSG1m4NV7a+N4U5BAjkYF3O+r4lAfT+E+LRdqfMZ861kofgJY
qG0PrgMlvL8yHtEPSrYQ/OnCTPq7Z+8Mzr7J5WgqNqQCXm8p92l4sQZpXOEi9NIEX/K/7M3jkZHz
Ko75AQEp5dJxcqKDzRuWj/vhhNWHda6yqkPcT9G/0wtlgPeKSVjGL6UDauoyMmYjq9oxtZAvsd/t
d3vmrjOt1JbbPHEwzSoaYgIETWvgisaW8jGdcyAJV6lTb62wVmh4M7r6Qs5oL/e5JqTIAOT2HXn2
V+Rm6QehKWW8RGH/dLTbkXHhKfHpH+YHMrgsTlRoln0+MDMBL7FbFU+Y+Grog2xi78m/94ymnjw/
W2p6s0bVLbTARr7eKDM7Ycu2E2+o+WYxBoxXqKc7EwI1zMh20IobNPpz5l2cVySwdaOx0flpqTGV
0YwoktHm5S3DMjNOPhL9S/ykaK+ND30ZIEbMPUtEs/nF0itoBHB6spLi3Z32Q46IPN3a87xWfY20
crtIumej34O9SUZSdNKnGD8o4Af9Ir9O3alhyxWuPOhsaFISI/HUTZxhwghUVn76esIY3QVPD3EO
K1AE5DJ+boK6XRa417WLKlcmAp3loocnHt7AkUHFREeP9hpVt8lhKr3kYmZm3/5mvfh3OQPldtOb
N5FGTa+3TIUIAZl+kc+9NECaDUdmein+36Ip5tdvc4pYlf6I+KIjg0ZISjaG2ZQdpqXyShNUqpCp
m0O9KwqemOEmUSIAwnggZLQdr19cAXZ4sjY8UEplB7KolJMw7bwjxqJA4Zz9t+K+Wcu701hvCu/C
33+vtwWzH9qIvQ5ngN/bVsthiw8j1DDt6MG5zB1wYH06yxumOnVPBrpITofoC0SjUeBEv2/wg255
1HQhxG5shTUNFcVJe0qF24IY2uQu3tf8a1UpdCivukPtc6H3foaTFRrjmoqAB1Gup7sXrMxJp07t
tkqNPJYLIH3F/8Nztg6U6fXsQQi6eiLCHr52szrFJJwfXc63K7fElWdlOBmJLYIgM5rCuwba9HHj
slIJOi95QF+6Z0k7qSBuC864y0QF3DlRELIUJuoEa2vL21Fju6WrebaqzqvtpEBC2n0T/UoFsQB4
xgVXVkRs96xo5rjJIaQrJgCF+I+DOoYdDSig2ZJvHEh0zZ6nsA1hHFGBY0bcMzg95O80wAHz7AJH
hzQXiHp57Prw3/nDR+oIsprDebZe0X3lgpUCjROFGiz5gAvCnP77EdAtO70xbcXPURuLePqlId8V
9+Olypd9LxnpqehGM0+UyP/PN2p7/4gU9ZslGSapWXtNFEg7pfscsiVNsxIKWy6M3oIFXdGV4Wve
VKigZNaWua9QfeGQn5WL/fnwoM/KXW1r8pQA2RZv7RFHVScLSAtpcIkbmuouUp754SLSse6Le/js
vOrqYiZ5gt8DYv0KytWDEDblxmk2kP8Aeumxvy7QNIH2tU90lwW3/g5YFacuGRStOIfMiDyFdh6H
WwVly4dHLt0KDpGNYJm0TRALHgpy+qp7k+cdJZQCxK8GxizLNXIoGs94v3lDJ+7N/Oacgrqn8CJp
7Lk5Ipyw0MLWtqiU2heomE9uzQb46xJI7RJvK3YbfWJXf4HA2Agj4DQKtk5jn7hcRb3lag4LonXV
6MhWlnYs9XOBAIv7opXlIYgCmkJW+m8W4Czqu5s26vDHTL2FFWMPRQDdxnWvr2d3vBjs6dg7abDg
9S24rwFIUWk/NBHupXav3205VAHgNcJS+6ucxlHob2LSby5iHLz5jwvq+AqhzqiVUYjoakzGRDHA
U9iEUR1fwhwQ/jjgiv1988ryLUdyir7MZNhmQOL8ZEIEYJk1OMfyV6iTvee1kXmotYTp4TXJ4iXm
e4E9iG7x5Xnt+QJng7bsZSpp5w6jdyqKHRiO1+Pfm0HdIQih+hkjlDnZKOrotEpELhzE32j5FC0e
QytSYqW4a8ev4f1j8JEyBv/LKTMceMaluVfTAd9rCyGqdumtm4h0Xw1Elc5+SKQZwHOjuNjJ00F8
QtjR5dnDOb1P5YvUmwgCmd7hQuTXZJNEnuhfWomHLQuTxP3HQMdx5uxkGNgQD8faSURieC9nW1ci
soXQJ06FQVOOZ1dSoyuOYGgQCHtRGNUrh60fpbmamE5tpdMeBcMgXoSTIoph/cppxM4stZUn0rHC
gDkDhYaewgf+R9P0JzsLXnCjoPOTvaFl+o8SdYEa33y8c5zBWazNkwW/m1OCSPVbPQAKxVdytW3C
5jVKezawTUV95ednZjl9mRUPs3moCQjzcPPO+PRlUzkjS/oBKkvTag9JpwwH3QiQCSnurU5OHaUz
9bXaks6asC5ZCTQ/DteBDDm5YhpBgmagwE1eqEEf5C7fvWisMlqmhBoEkO06A1Bs3ATaHa4DMRq/
mLDzW4bfn1FbpBJQ20SKcNnqnKpY472WBxs4PDKvdaE1a5U3Fv1SArgONa7fw7sUcg1msM24FKyX
qSiNp/lk+D2XbyIAryvQVUABVqNyVCKinqFKCiMvzvKNPiDbgVdB94V1Ca5HXcUiPhRBjmsqiD9r
LCjInMJmRxD8XSQNUIvLAwKHhSA3zdnRlX8DLy98r4HiSle4SsAH/dMWYWRgXX1WfcH1K2MdH3Ka
UynchYIRiClFHGWH5+OMNrac6PXHX788l7z2M5En9KEs2FLjm5tty1M0SGYvKWWobSY3s8eRAxWi
WQRDj/7c8BiW0SW1JyklNBcoJPByiADgG+O2DY8KdgCUBob4rnZonmwrIgV0v4tFLVXull/KPL3H
hkiufnT4cyfRy1SxZNnXWrGhbJ3GbBTs069RaYJPH/K9sc2xESC7EGmLC+4P5ZwEZVyQcaiqKklD
Mqhs+8negn5fTA8CBK965qU3U1WGfafowMF2JbZ6vPB4cuPknntQwh7hLoRpxflpTVtGirhJJIv1
3z72NbvmM8tI2jh9nKEfosp2DrLARBRXJI+jK7Ik9CtS56zbPuoWQy0MTg62KnAaTeXTVoaTLMgi
M97noQ5AaPKqfbfhvL3SXgsycuDh7+euPz7NgV1xXDpI8uKjqxUAV2qu5YJvrUuVCkuT3BGAXMUO
bS6tfpReR1AuitzZDsxunjFcc53dSwcl2nA2YtZkEIZqeU2pCjtNznxtSy39i6cKsgB6hi/aCvdt
W3QbpuN14e6oxbfdlmAL9jR+32ZmisFKmDRqsVsVWZ4hLbWEb/2HCejAQ3ulBncpD3uf0M+SGlbR
V64N8nytOVm9EDZOgDfRmrLRe4entTGms5+RyNzV47Sa1AJrsMFGsY2F/reBQeG7y/NlvytdfYEx
YjDKoelzLkKrM6MGO4tBqX4gOELkSC9fZWpth4X3WEcTLH1mmIoz2ehhQ/cfLSXnIiQRG10STRAI
0JZ8HKSxCITW2NdOBpZx89Q1ynm823S6o5CwOvXBKWDqTQ9Uws1wpCdJ1/u4FvQTRahF9nMafm3j
UoxjjTcDmj9nbVsnbbvaiR4dCbDjXDpD0VIi8xPBwOYuIkXqlbgUJ8025bPriHwCIe6A2PGxDaXz
XTMfHQXKwed2TYLw00AI9LMvczrzao4IsXtP2cLQGjg1KySWKQkVzTPW96pB6lE6Cz8aDyH4OC+d
ESEEwHDW5DBAMq37y0XfNI/rpzQJCXdfarldrbBK1dpRgg4j1gBdieaOoszmWASwC7K681akTc6J
b8NgptfgMczCil7r3eRHhzM4g50AC7N/iW145fXDWzG5UWY5U4lUgENFbdMy48Yn/5paxmGoNeMV
9pnP2JtEc26aLFNkhE479bJHZDSRSeQzVcto60xYLbCElnpSw1tev+vE4PehRMB5gfyx7UXgZPSJ
fDNeyMEVlDd9fOdmm8Nds9FZsn/QulS/6uaVJJDtr7UsJZ5x54jQt4/L/ejMfsxlKz0gvdWWVFER
v3EoE0BOKO34ZhpdAshdQGkzQ8dRMiO/QXi76cAW0ki4Cb8bUZ3h8xAH67yzi7jAg73s6V5Jr3N7
sZgz9HepqQGiqCl+Ez+0fiFB5Zppp794upOgi46gkpRbV1yWSdAAdcGVmP3F+xMxUyWV6xr/vf99
GdYXyhWvUxuCpJtBTcHR+8ZLaRPqQJxkBqSct7qcy6uhI3tI3tQqq/csYI0OAxBhg/QVhuDAZMCl
NgX97MB3VLY4bCuauvKhGCGm4iZzYqda/nq/mNf1kQhOkoZB1NSKKGtyI7f4ISN8WEUx52gLbm9G
Xj5IoUZfBLaVWGkHQmDk688o9mD4Poj3O01Qwz4HHwFT5yttGWwSFKnuK4688IdQj0YUIu2fi81f
O/llrp8eMBQ5hx7Z6DM2xohgCmGSERs+DGHTPgTMg/RbcPDUUm5Zj80EIZIxw2Twvxd4AZdbos94
KY4h+BiWFDioe2DGRTEgQ2idiRcTdKjnkh1nXhU/5py+Amg0pYPtjlNF112w1jGYYq7b9y2iQHv5
Zcb/3i1b1dmpW8tp7sPub4kaE//0OIk/2fWfa1B3d59/AhGuxPuhFOK2Utd0Cl8IsUe2Fho8JYyi
o8vWzvlG3786v1RH/fUsogkAtrkm593sEnLvHRm43IGQpAvWryJbzcPnzjL4oj0/cj90WgRKPOyJ
P6GG3H9ldzKDJWjq592PN1Cl5a9VQzMj1UNQ4I7+dOHotp9xDKeXtPmOrwhFAQ3n4p9vJosvjLGO
PqstWZrJHSsW+AjLFtxzt28vik8QA+IS4mKynAxdAgy2G35xkoDiW8Ujn8y2Bjb0hVhRvZN4O4JG
5b+/nJKCneFpewTPnTOngTvT4ZRuiT0p8s2l6bMO/AHmdwkATTtTtHTiRxqbrTH6w/MEQtjijoC4
D8BoFQ+B/9ZRph1LRlpIFONCPCmQkbIOJLdemp2rfRN8dlAgyVOvPe7U8UqxVi9NIGMxu6qK7u1p
5fesFEFBV0brG4sdcf/fXt9LK2gdwnEinX7k5aFNBvKCehmypcBqKjvSuu84m191DnsEg0xIhDqa
H03rEIi0m5GkWPj53CHQ/ElsW+K00+AwYtYMJ7UvQlIMQPwknTdWTuQm1ya3+TN34bb4J/sfcFBC
kq0ZOsOFT88g0FycMyiKfw6SaFM9tlTIkItVzQWgesRzZRu4T4pyNDVpxIMxdOU3PpsiJCybglF1
yYuNGDBaqnFOOP6Y1M6DDykoqVBDdZs6tHnZDCLlTBmiODP0JUdLH2wmIZPWHw2QOPJVSveHRgB3
LLATUVb2t25xrmd7QcX8shrUAQ8mp44AL9qvbs1TohGl77rVoChRKsGG2QPDGo89ym/MC4JMAaYq
hXJRWH3qgoekQLsoQA7yPygkbCDpJHLHPyU9mq8gHborRGbceQlvCaOjPalKrEKh84RSGEC/NMUT
HD2/0J0WDJPkZdFQwEokDpr5YsFOCL5ynXjnfpI0hHJOTWHsDpvpO1KVpz+bNyfmdf0EPcaHMZWc
Rw4hyZkKPDdTUkMUk2QYGvojslH7z/VFvX439EuxM8xErgdEUOU3rliYY99QbBD28hJGEg7HMuO0
0rsyjtYH0jUrFrQ98oY/wqJ40KyRJ4hbbzHBZx3nXUxSQc5gQmiNULtrrdKTYoSZWZuez9OfH0+T
si1OM6vXRYHJfUoGDjoGDxyulTPYLMmfLUtBXPHyuJL0AKzeiZKz50rzPsQg0BCAh4R8G2y819Qt
hsTZVes0DRz4zXk0V2muNl10k+EJodJ9r+Dl1TYB27nBg2fecyfo1XDsde6F4ae+8HIQJ3rKzIux
7gKg9Q3eozF7TKCHBi0OtmGh8eO+3HAkxM3A5dNNfGlY9YaPYufkzcdJ1Ug+KCFnmzybqmyag1Lv
/1S3c7VfqMg0O70BAn3LbF+W/ulPQ/hqqldAh9gYso2o5B2vpypvvOgRXTTW/oxXi6rSRBIpYLLq
NEGbL1HS1MalO82HqjaZyQRDRH2xbUNcM56yUZfXT8+b9w65h0Xyz3SLTtA/BoLpnBwQwG2ZOeJP
GTcATWR64RD8S5ZZuL0coWQTIhosLRILx4RRTipz1hbY65w2fQq++hnDN9wIcQL3SBQsOHXsy874
tyZoeWt9vDVN7kiJqJOtlj72djrswDB1YSPh16wjEga4mjp7c2gJ4GYEUxxgJAkJ/kr9prJf6BYG
k0vRNtlHZSSxUcfsDakUdy/OFWXQz3FAl2x0no6+Ks6YqDAK8eQRsQ4jCf/JN5+hMjJMbew7RGNk
0rfZDVeraVObmysWtJJzm+pVVD5atOPek9w+SSRGHIF5jQYsHFDC4UmNqhFXzTiSqyoJjSEME+up
3FoP/jHTpIlpoN7TKBL6XyaWMX9DZoPjX5awY/66oNz0Jhx7fMJ4JutyxRv8cSY1oxX8o9EKyBf8
GPzhlM0BQcVhJ55PtAle2jQMe3hRFVlooF9uy6b4NxoICz78gmq0gw8jqjToOj5WxZI2zYHeJDrq
RTTuPr6YdL9JrHoy3Zkof9rOgRrgFvgQq0wrK0r1FljXOzG1q+0TbAoJeHAMHIZYQic+2mCqoMzc
rDxYZtwvv1NsJZJcBcbZukIQ1ZVxrmaBGclJaL0h7FVzDy9uas8z9ew+e1lUK1htJHVLQRPHeAfp
ypeIVTAS05aqD2HB1xhDKuJ2QZF6wCDKoXF2BtBZ3uj4F8200cjJ+b3bQoIQazdSrl4lko8QnnL2
Ix85IlHQjyzlwnhi3s4rlGZllLlAFCKZYrz+T2ZZfUCHlyPcNsWbv7dczUqZEYQt1d0g4ZidS255
qvNvZh3D6+S7sBsinmJzhJN8XBGKHhrMnVMgvXx4R2IxEIQ8Why87aJeaCSyDpLYSmiFn5hFB91t
+SN9umKbdN8kxkFHhEWCAn4oq4o1TSKFX1UJZTnRMfIMrmOIf0ZOncJCebNwigAxtBbUAnt3Tv8h
Xmd0OOTfPP+7dwWjAYHf8pU3nn1H/VX6N3TLSW/zJzlrqGmVPBTWezE5OpSU8pL/dQ1jdzcxv2eP
edJkHX9GO68arzLWNzzXIa9XBAyezkU4eySD4z19cLJbwgs0zaHwohEQBsxpagU9sDc9SF3mRMh7
IcyNMfpkKMhAAHpW11bDZeEW/FB7pVE1xO4L1utkp8FV/2VRZq7sCGBOExlGefpKL0ZoFhcQYHpr
kgnvsTHEgtgTbYsUUN8c8W89kZv0nbH3SZvB4/oLZeyWaMR5j5kF6kat7HMWSrhxh+Ss7X3FDsKz
hXpHT7uZ1VhA+oFcEpwRX8m00RwK1w0P0ZOlVwWDiSMjfljciqg1udSdV4m2tAjMDeMybTYaUi46
JEyv1MZSP305YMhpSTJK8b7iu7T5T+TgAcWgRlCzC2eXGBY+OIfcXXzi5ZpwNdOH5yc+F+9oMBQM
mWVmkinJkZmosq+ZJrPsULCS19bYG0u6+maJzmywCBcc3fyNftVYEqEatCNBTMLmR0XCraQyvYEr
UzDQ9CzVJujGciPOj1+ieGNgFZy8+P1qZyBr6d7Z/Rz5bBHh70XG7LHWN2ub6HwH9R418U0Fh16V
T2uIC8zViL5SoQldG0aNkIe8NBE/86eD3l1E1MhVwomnui1PMtsX7zSZBPeB7ruKRvEg6YGdCRfC
jxC7WMFVNmiBuuEKArynamqzO6WQgkougEE6pEhL28zqwOQuPBcXgwEHmgXlGQ5l3lUvRlvPc9Yp
H/dVJ+N7LL3sdLKJ4Zdo4Pvm4Yn3oL054XWTRGg0qHSAdtOL8kUlvH5TQkyO1HDDOAmeRsVbCDvr
uE7WoTNZ0o5q1y8jjwrqlNT1t7rnfVppQayucvwuyu0ysA4bdhgIYLjNC5eZVXqRvaaRx8dh2/9W
5vD9j/T4+FuH2b7qY4nEt78GQLNnLpNg2luaykQuq7EGL4tqHeRSDmi/eavk8FFM8suv+MzpiQL0
bTcuviz4hzs1U/186RcanYPTqvfgO7JLTg+Rn0vEHgdkdBAFd1AZaqjjVSbNcPWzt8cVVFwyxohW
x4qRi2K6eAlw2EjSbf9BPZRAc8JK37sjDupLJjHYypI36KbHRy9ZgQS3J8yW4mZS0bMGgTZyb4V0
MdznCE/um5zMKxmhuqH0dBoCPK9XwKHVIddxa8xODLFzjDWC0vpOfyfv/7EYyZRJcnQl0pOp9N0U
JLPQNYOeWldOcqGaPet7PAUmQwQ3ADc1SS2RBBcGcZP2yWtTzRfBiAGRkMyoz5VX9IXm90PBpo5L
k/JBmowS5dI7HvYVE+jVCuk7O58hfXzhB3UAuV7xqG03C59atvhO2b2LwRt/7JY9mpMbSAGw/DBR
/WGS5x5qV6k5JN9g9dMfGVzhf0DkNgQdI56KDUTHA7rOzeVmzW2EsfT/3MGEpDFFVrFHnN99qbsp
ZoJWW8DcsgNtU8gCP8hBV7tJtFWp5RmZ120/rkU8tkhivH3fNNb0xG03f+B20QWYAuE6Bzt4SNt7
BJtGKLYfT4IiaacsDaYWlvTBTyhPEj0fOf7Jhn4OLKlthoyxeHyfwzr76NGgvPHhar6b+LJ6gkIt
B7cVpOGt3/oRPz/WvwQf7DO4eQI3NSH9Rs6V54BlRCaknDWXPOTd60MdZscwJxukx/IaK5voBLmb
VCsmv6woW/G7v+YxwXIh6vR2PdHmd5D1MpvsEpNfj3Ns7EfW6ZjGBEyFoY1BCjwmfjY1HvAoKGNu
Wcc4GxALog+meuCWKGAvGFYr9SoKVwj99nvOuaaLFTI0tz9Vd13WDIF5stShiNeuR9JlQeYDGinU
Jqq//5WmHRD7XkC9ERzc+ilrvA8MqEAzhMIVhl/RYhfIYwvjBOhyNXCRk3LlQTLL94YKv0nEtlSl
nXDe/bI5LKSIAwfTpSOtFJUw/WIvq/7cZkkzWjZ/wlHE0Ro2OUGdV7DE2fDZZiKMXWA794rsf+w0
1n6Mkfls6qMKqMI3aLwon2c6QzTZjqJ4F7JPxmL9OXCeW9wOyIvtov5sIU51WDxU/b6I5bOLkOcv
Pwi4I6h+XHKh/b1ftNJC9VSQwQDEGoU6esMgoJmUXZnZ2/6+KFMqVYv4IetamKSzZqbRe47rZNRL
PhF/jXEUVlpx2WkCrRRkf/2rMRkSsT6O2W+t+3rvsCy0q8J96cBdSxE4QMtx8OlLh6/AySz7KaBa
MWnt3JijWPeJ0FHY7kYVhfalWtluT46e5OQ6C5cypryUCJAAoA21ePSRzMReNzLodnVUi5BU4kAz
guFOWRTe/sXGrB+5kiAU3N5kc3nEvCGQ03OIPTHFc2kVny7MTrP6CsoGqAOYQOfq+u2x9zukdF4K
Vwf2laZHUCh+6ckEUB5TqmZEOG8oDlB8xo2H5a0QGkbGdTQxlgFC76NKczDTbZ/OJCtBLKyPSPU2
2T1IwLyRGjADzUwzbpMbjLtt9y0A/BFwalrQhUzn7z0+bXR5GABcKRPx/wuVM4aqZtRDIghHRSGu
tLosC0MSBAvWBuyGrtuFsZQvl80eV5yS1+eA3JQgCGgZ/Y0TN4pVRM6xH0EKesWUmYiPemdx5Ngv
cJu7UjfrX9o3NEGEYQOgb0+y1J/yM2waWXxxhkuJg8k9DSJM152ahiBh3jx0H/ET6WP6vR+IVy5q
T6Oz/f+9QufmMJUVibpkJKsKsPZ2mkP+i/4tenVcxZ8mIxoyRcXquPMEJLVuYg36k56XviOgK/o/
dt6K1Q6Rwej14b2th1nmyQRekttUG2mc8YkhGLJ0j6kylxHbltzW6j6Iuj5V9hxd6SWQ/Jbop7IM
xB0UhBjjdNhjMyKR1lBO+bsKtY8U6NpR7+isM4u1U+nH2erEvMqMuatAkUDQ1MMKvIo+6QKXvJ6X
+8y0uYlUL1x7UWM9CVWfWIB2AIqi/kzQevSxpegE0HANKkXbFulepuhafiVsq5F1+z5hf1kZVGUL
KEgTeMVzTIYtnlZ2Y/eR88Fij9ftn9kJqxaOhS3vsh7UFiXmcHjiDPqxFD9Xv+XGpWxLV3bkNJCc
vpHbYR+TFSKX3du5TT5h17WxJftYwe5NY5WyX1jEO6W1N/ZVA9/04QPGumUfoRZ29txZcrQGtxcW
nMhdS4z0ZUS3ijKq/sxJZ7Me2MiZKvJEcHiH9U+DooZv5iVYeQ3fiJrl7atyoWEVHiYKdgOViI3K
P7U4cM1EmHa9UrnZHIGY0+Wj6hy3sfAe9OORw+TVpOF7T2TlFLfZ13T/704qFIeng9I+Ubr4qfAc
Z+Q0qVE0WXWiFVXvJooRfubKhvAXzRg8zNOj+5/fGvCRWRGp1LDuQIFl+ZmajjwIOUpLP/HHMNN0
JKM8Y0+fbJ3SjOx2PiaJuNy0dv8A59pjS/hXlNO/lx5S9xGTRHJPug1Ig8HbW1AHCJpZj2DcCPbD
8guJ3lbhTBMd1GSXtDyJttKB5lIgj4AdCqbcMId+TMclRgROkZd3he+U4OO++08mGXLR+LJ/4kkT
V2K3gYjulTkYeJDtIVwuRR8LXQdp2vgMygMpQoDdfDMJ5Pmffvn5R4ZM6WC7jRB/110x8EhWUj0W
XxnZAzz/gV9GWXChHbqhbFPuSs24+6vnNusn42WykZAlDASe1GLlJ9Kigqjwhc+k69Opm9Wfn5+1
j5Vgg4DqIn/Ed+s2S/DgY7xrr18sWivSMwSw+ZCjuGTFI65pUn1TD2VfReybWRS6UajqANFq8oLy
6dOu8RlVORqpGR30zFB/E7hHJAwSsizEf9XzP/IKvnyALcwcxpxi+pzet1DMY70+pdrW4zmuWS7P
1phj6Y4dr5X1PMuMUHWF2Ld8Fo7aKrwtC3Wbh6DmKEYA0znaxXZT1eIh0ppLDm2eYNVdl5PwEevE
x5sWpw2iW53mtjI0O+crsCNcdHbmS77Ib78VsRoJyq8RIB84f1LvOrmPlFLaRQHWz/l2eSrRuvxs
Pn155I+R4QCLswVccgojuTVJ/URzlJ5gIlVdA17bZBLEDOXq/4KGeJ+mmDcHoSWZjSc4bYtXeeLR
R8mGs558uV5hHwK1GBXq8LxEJ/uOLFYN3P0PbDENoSbGY/ORsL/XXqLhnxtQ7c6bf7/WWdrmacPB
obisIqJsSLlJCo4zs5Mb5MI9eHIIIx+KNO/RVfzD0KtXFlpulRP39M9aL9jqbOFwJZkD1DXZPHCS
p4Hj403oRf7uihMzrozwZUQm3QCg18FdmGDrcIW432XkfovXJK/D+CzBfur1f/rOpVo48CqJb7TA
GqNVLIQ8dErPZkan8bnklHVoS6jEYI6NPfLtmkH4JjzrJI9YHVFQZgr1s2Lo3ffY1oU0J6MmK+cA
WdDXV+WJe961SR0KufLvelhuo7K92CgZKvwRvq5lGK5SfB6FCDYhGa6vm8E6MuiQpf+qHo5Dv4jx
X46fPwzdAAyHpynZ5wmrlSXm9lCZ3JovXwG7QEaj9JXCgwP7PgKENx9htD5pmMUiUoFZDEPw50Bj
LGS/ToWB51FGvn6F3fSuQ31Tvj0qxPWPY/NehjAbPnncW4XTxiQ6DOAqs99Ip12DwJfEs15lmYHQ
0ZEkSn7hB0tASB8W8fN5Fqv4/InQMUjrutMklZJIT0RGb9djLcXUd6BglMj2xFHAaGs/BKoOdA9A
b1Azz5njzT17CRFlafdnTskLyMbXfUZpTXTW44ln64159Zuw7KIiquMBAOjc8MSv7eY8/TCdayEa
1X8XxHERfZ5z2AsYI3gpb5nLcXJp3H0OjSCrj/m1ceLwFf5tp6l8YNyiyvXQicj/M1sy9eyAq6J8
NgJGSshGJK1eC/ZlsuodOPXqk8HRRqKTcqdaIqnP6C/bpMmCcEhq52WSdjYhfaWh//CRJNagkDJQ
xBztJE+6nd4X2FOkTpxgULGRkhQI3H32Z+hnWTM5dlhrAXsVFGpkNQSZIhUEhuZEX1aIxL+nxXiG
GgENkyiqiMAnMdFJXRuc+IG5SXw8wuqx4n3mW7QNHACaRSE7U5MlZDAbIaIwmAeHdmlcSuFCpMai
dpetkbRADK0Gf0Y81Hk0rn4SzD5gaDZsbGKSUpKfeG/gvpcwgvt1k9K+31Loy9Ud1FfNy74oEAZk
HuSqeNlhXLEsxyFKqJYe26GEEdMK+7U9FKfOImqDLrFE9kCn9CwSlJEVYfVt6ZcKifBwOnZ31tr4
2myY8A4brcaEwPedFeHBykGfI3UfvwZKTGHMdIqlCfcXu1bZ832FT3vnd6aXB8NjGIdiGkH2ef5Q
mnAx4wZM4jWj7WH8+yx6jsQiv6jVGwhTab925y6sFhc6AX72zsKu/HXE2UnPNUD1x1lfwUjN/x+H
oa9gWsOyeLhIk2ipQrZWX1Yy07mY2uXV8R4uqVnX45gM/JvwScwl1lb+tStepUw8pkp24VbcW3Kr
q8/UFRG1ahDm2oztKRhC4OKCnwjUj5oilTSp076jin+zbvYjXs1SQL3osfxoY4dNmyukXFRCO1yk
44ZGrMcXVQaKYofBVyTtl6Ic3PV2bjD5EBkac/tNXCE+PSUqE1dS0/lZF09bxvC39mfSqDNldzD9
INbhsGN2VLABmJinfdklDv48xst3vLQD5IDuBs6zyegiS5IL7dKC0WBNu8ij/Gtv4MgIQWwayLON
21NJLInq8ApCDgIYmPpTg6a9huDy9QZtOPrpI1ly0Q5oVsUadC+ZUBF0qnE1ulBdf1CpPKol8ja5
PQTWbz2SFzW4Iy+4yeeNIx5JWohWvgrOTPFYmvZ/5f2Rsq3SKiYFM/qF3y0AoT9np8sFUYwD5hF8
PtyAxBEdWcDDIC91Jt4ha2M9siMewUoJoD29ynmfP0bWLePv2B1azBPrvubfcSRLcX7eUeCGGF0k
CTAXAmAdWzut+a3zdzFCp1iycaKuwX/xNy3uMX0huHtYFD/Iy/IWkbWjR6kxL6wfNt+437bs74bL
IdqYkis9xLJn6mFjUh60i/gqJFCUV5mt8p4N+G3CTaBqG7un4JgodCCdSPh3zn+CdtZAybLGoCnU
IshDI9Q6QjNRG7LKWN9txw9T36ZotXfpTtrJSWtv8TI63i20l5FmShnGqPQZEFZFQUIiJi/H8y0B
2OjqRFjzd+Btikg0+72ddzdvE4MLU2KgcEqWg8R3nN+vi3FnATtbRQncikEvGwcmVd/9OGdMcfEa
iaOVy3ziTQ59dnGtq5QIYGlY9A1oyEe4+a3ezukD6vH8M3BtWDhuqHmTH1kbLD+5s5z/T4OVwdKc
frANmDxgXhU7P5NbQVnBEQKPCF9IymSVMku3mRIA2LoxRZZSYhe6CNYTwuOuR7ZDIOaE94sZRddF
C7rGuujLuR7PWlh8Yyn/9DFcEOp/s0sR3400X7d5RbETrK/dYvB+CluXl7DImWFct9zVtZPHLTed
zH4cGxldmUPT19M2aSQ95HvWCUB96f+J9EoNxXl+rUWJkaMzJ8bnJsI4guRSzjZtiC7kmaft8Tpd
AvBx7CmY1StoIssDFUQm3ERSTuYVvO1Kl+iK85iQDuYTA2kRuY1NHT91YQI2SIHTBXTUoY1Gj7c+
mDZGyRdbWm2AMWFmhjcc0BxyKvPaHWzEow373of6WHBS5j2McE0hRKHJtFKLdtb/dNAkNuk4OZMS
ve9C9EIZXbdU9+hjOrouipho+lA0Y6nFou3ggiAviDzvx87/AF2mmqLW3Iez9JQm6y7bNmmpWKvA
Cqe3JzpWEY2L7DC8/O+oarp8Br+AhEM6W7a+8nDsn6Aat1PzaPy8SHrlVLIuSvGBkk9UYLfC84Q5
UoqTNb1OOHhrjSJoC8LKyYhw7EBmX9b1tef5do0Pb7naXqr+OTWdiAzeKeawvarbpoX9la9yFUss
PBdjoRpAVKdlojJv+w0xYqlkwnXqCp2SWjcTGOe6Ah3ikCPE31iH4hqExTx/Cff3ssYmSes2EFgD
vf7BNRKylshB5QRnKB4KIf33L1nL+UtUW65czG/Nu0NQhNBA2L+y7Yx7VaHatnOMItrInwVOi5sI
/vIXdKfBVPfdtcF3i2CTEyOMDQCNXNsQ01SGJ0ZhkrWe399WIdjE+wgsL4ZhuXrBjWQ5mnHKDNzW
nCasaDp8cBkgzwOehAUfAqkuPGIcJsiFDb/gvEw7Hvx4yS1lMSu4On5jvse2coD/9RfkcmNPwdAV
bCGH+TYGSSaa3fOPZpTofKPsevsEUWQ5h1BCnoDJzPxea/+Xdv15p+WeVcO9SUnjclhEj+H6AzXp
ud1o15+WdKj1w3MB33BYEoGIyE+eCqF8OE0fEDFm6izpiyTEeHrzPBH2s2WFqQacdWTJ1FrdkYtf
XXCGCsPlpDF2MI2VhLSOD6h3LeWXte871B3L+d36xf4HkoZ8a1N2D9VY5UnKYdx0X0Pxb+ofKnNP
DRBDmUzPDTiV04USSkSjYh2QbhBvuWIK/jM0XA/0MNdcgeUZcyQ1ynhyed7YHonFF4QLByeaTXcM
tZMkyLOsA7r8L7L6ELWKHMeq3XpNWjb6qrl8/PsxHxWzM9FS5fm6+W+2/Kr+7I2T6Y9H2SbVrExh
vYRsSI/bCSWOklqf+Mdms2B04hREi6IvZqTA2dNHSb9YxJ84gqldHE1iLDnnnLG28NFSe/zsS2QV
Ez2qk3cc2x3OjWdZGeTmLAB+kOc5gj5sSbgWbkpwhE75teszqIt8IJmr5H4s4cuwWOpJ17FtA3YN
FCVzoxOyg3vO5Qb1wapdgrh+3nhHGc907rirFi8cayChNI+0B7FHkEn+iH3tpQxOhtvpiQH+kcrp
fTr+FF6BSG453Kf5nTvVKNwGW/RDD3wab+mAtA3bgC7wIa3gVO3YGBzMycgAvzuKIgUznx3NV9Lq
yHwHjeX11l85Xn0n8pshpMlRiCG+9c3Hb+9K9egpIpqrVHLr/Vl8lfFQtdG2aOMcIYBegasBfpAf
Nt5NVnOE30V14GEvJu/Z+dIEyCQgJN5y9cn9n4Id/pY6rTSmbB7x100Mrktlrjnt8gtHqSo0yyzc
LdWNHOakKoUn7eomGwIanXdyLpnYzJLnW6n4gRJ74P/2Q9eY5nELQOBvAsI1yTC4sHHtbZInC+Ig
ILVe/c54ynbmCv2aOJxlz19az07v3H3mdGezRZuwYtByscsnR34FGj69bMMl9NwJYsCHn8glUxdS
WmlZ9RGFlt8zXruxu/FLzZADV/xFLDvmWm+Lx2E8s/iEpp7JVVudpJVvgrmZqdki6r3M5a2WI5Ju
RJpOzIomVvKJL5OJbhKl7Wog99lMkzTAEl8ZQNw9SbXuYNh3b8jTZK41kEWRPYCYm1vZ2eu6FFVW
MF3ouT2kzjtCtLB5MyHQ6qyA1fRHnaeY4oXjJmxn7zWGzr1W4jCqZF7qi5MjGWFtceEgGewqi0PO
mSMv0RmAGJt9Pa4r0jv76Jk8ZqSCFhY1OPYIlcrQxB/fxfMvgxNafDPud03zPL97JYBnxlKRCdig
wClrxnxQmzn0XpwPeCnTmX4IquUyHf2gp1pF7XcTtHNSGObEdPqK5E9aQmsa3FVzjbeRawAgHGmI
E/aIZ2FTjCf5xreEny96hAnRNBcDmdKkuu7IcncFS80PseG1an5xFBYmK0vG/YwwRzJt3dyAnRkh
1C5xsJyZ7nEkluZP/tlmS9thGWK2R/N9DLRv2vmx9ynhtwoDxaQUnDu3SA6b5gC614IQQCbkWSDQ
cFTFL8CH+8bV/qfEWcnFpJ2Z5WiMuZiF1u/R3sloKErz8kbaAjV9Swo6Qrq83c05cZf9c6Ibus18
aAhxXx+m50khqGNI0BaEN6zZMBgumfaBr5i/mxnP7GAGBrlXOT/669ukSXjIDGcLHgXYm9039x0n
3NyN8pbF5qTQ7v3kX+2gloFgUBn2lVPNKxFmisu7jNm/UtMeiHi+ZWblIB3LEphg/jtlFFxrDJCF
Tva8eSGTtcsYryJd2c3jlhgpYcSuNss3hdyfzLQ2y35s2uMmrztgwGksaha/pa4vdUM1ro0+gtVO
4YI66J4WpnnRSDkoYzkivsLQrKSD+6vLgz6f+1SaCVdh+pjqrTCmdoJKDZBnUeqSVqIM7+IdrS5e
SLAg+w/FrX34jlE3k2HpsCC5LOLtDuyai43sIIX4/TVBU6NDO4fJqUDh1BYd5NN4KzPYltbnqOWT
kGXg0EfsfhOH93ZuIHeTFyOS1nOQqFYZQ/ToT2IJjBwrOYvz2vCJKEd3uef/BF9Ldtf1kHOAyEhH
jdJHB5+oeVsZywaEAJusw6y3gkhLXJtX9sFyrVvriI2234oVqkVarTEuq7Pt83+puZ0WNP32gnwv
fOIjrkym6vRE8TaWlbJChjeTeHWd/rKHpV82U0VIi8Klo2JfxJN0q1FVqAnB2t2cRhE1JgkNyLYD
/HX4knZovF1TmJxW+1u8j0zOMlsAI6MNLEMF/hj4EXTgQK0n+hveCo5jpLxtvvG1cOW9HU+wJHnx
3Lr4NerhE8sM8H66Iaauw4Ev/HakZYYPbyWYgYNPVHK+3UoFU89lWxHukCYdbwh9zwTcCnNlmTG8
TKL62dL4XqiLnDBsgMSBWAJh6dRc8lG92ewRb7vr1G/vwfDGWUGfElonWFhJszFVQI9nLTOFE9qf
a7Hcz9j/FbmdJBd+ttNndppqIzoY4ytActAZ6NJvjgpNXQ2Bg88/6YFZknheCzfSkdKTcTDxco+i
K+PygArYVpcxMh+GWOHq+IHgShpgLOzl7YU5KVgybiPQEh4nB+/ID5WL9wwbXCFUL7FfkpZu6TJt
AyxZDKbDTtzie/jbza84KmyvA8t136uTAR/5xeFdoyWW5JiesmWnUZZfpzTEzKOaD3ZXBa8MK+oR
mCChEyYaIv8si8PGwIFDYslnOssAn1Sj3IopFdubmOhUzDmoF+7FshOcFHDao1f+sykmUkP5U9jD
ZddtVfQpovB4x8RO6aHVSBMOrwKVeWfir18OljdbdkUGjp86Z/U2hVkJ5ywABDfDEmvdOwSuVFFk
52hipv0hVXbT1TUDTFmoAVlOTEvq+idqZwZRPTGVQuNjJvRre9sbk2ZkLKEdWrZN3RycAMCzAbYI
JDKGtRLoyAHlEtLyG1hVma0ke59luG2jpwbk4VVY6o9BB2yPHQpyKyQeRizqnQ5mOlq5+ZFXr1W+
DIgrYGuCt1KZq6Kmg/45MD50dmtIKqJlWpIkWK2bQlzMXw1jA2kvkrCihs35iXI0KQYoL8XzbzyR
Xq0qsVGJZcA77I/SsSIbW/rQlElejtVTLfcxS775NVL0zeALBMJIdcasI+KLhATcbPjubjnpzGL/
94qGHbWQcaW+iIq4OoKx5d1dkr7fnu3N4tu3RM3vRCivocLPrXijjULml+eLNA3aXvUyKv7jJHMU
/LD3GaoblFB+TgHjNRP3SFJUnLcJjtua6/ByjZw4L7EKLYr0af+UrpJ0XV4zFzJ/qV0Z9YlKLONy
OL9Ifv3n+ZBiJIxEaT47KH/dVKMSrF8g+ZCWqtU6O0st4uYg15Z8Fg3fWmqLhEyyKIl6DUTtHLd9
Hc2CvFsdB60RAm1EMt5jxDiV5DaZH3PHwFNPTwAkr8GYD7PULDq39eUzymzP8r4CKaV2LwvcXfat
qXb/uydzKGVuqoflUEgJZPCyyseTwGxbn9pm1hR82L4Aea24MVX1ZvE41jYHHd9cyWdRAyEUzWEm
GKFMYYgaR4xSX9wTkRTHUweOah0mRISMhDDyCxxYehcToyPa1OuBxjmIHMXk8M1syStNQWwcxuHL
7Q4Yxaozk3v7FAVWUaCQhhOGlmqQCCgKAQiSmyxIUAv+TbclGvINbve24L6X9LCVqjHAh5HYAp4w
dSvqjz1OxlcZat5XAYllXF/HYHLjdmRzBL2r0odUp+1VIl7Y17oldUgfoKOEtokwFTBp60xo/IZY
eHNmYTj8WyQbv5lv8ax4wTdbCYF4jM1CUc4ZWUtLaTklQMekDkqrp+3dsFLX0AQjZ4YytGAVfnGO
8ausUmdqMDVFc570mM2WUIGHp1U2B/JrpmLKxjkJz8HccDO6Q0Eumlsg9RefHWM38LeFFdCyE1VO
NeMr/ELq5mb8gO8biygoYnQ1QcsIDgu0ccMdW4gHAyCGti3hiU/55B3ioYAzYvyVlrn34bgdGBI2
85oBepDSdG1Gq1zE0elJvi+8jyHxLU/75xULETZ1GuI0i//PXIuwy0+8PS5EK8ec8GfUw5W2mN7E
hLbsnAp0gH7SniQ+Kb/PrYLlGvGYLKrt7m2BXUoUM6Y2d2hVIsdffAn/rAXKNjqCqWXJFOPOIxo8
YThsMRB4ZsKKLpJ01SfpQa8Pb80JSmdnrn8M8ORcJERNhf4MkUnNRKyddC8Mtg2iifwrmO3tO2AV
7qWyfXCM5qm7GyJYyaHtArGffvq65+EkC9J6hLm0JOLXg0pKkUGiqv5KLG16OGUpOXqFweXjqeSp
4A5m3ZmcEC0Gwa+8R8tlUAdpzLmxVmgJ4IwBlNIxhTpU+TXF2uAY7tikJ97mLY4w0pCZ+w3mC2hs
khKt8TToP4Jw56Xm5LDdpwEZ0lKIeT00sKkSD+O1rXXmySX1qOaVJAsC+VueaQrmD8kpsKIqrhj/
RB8o0LTKGON5arGbJCK2ZDQvhArs3gp5wbXtrpTsVF3KkXwIiG0XVb9WIvs4PkCZOalNLBzNN91T
lEbkKxR/e3+gKZU/bIoACUSIsFl8yk3R3scHG92y6XMKLUwijK2wOzc8N/zODVeUUhSxT4cp6Jh5
fZIyRQGn6yqU0T3MK6V56sCNV+n/sfMV1Nn5qK5j3Q2cBjsS8jzSMNSpPFntSn7Gor4mKzveg2qV
Fx4FAenaUa2232zzupJr6dTpKNM33AF4sdUIn7BobWquyWNB6BJjwJ6rNVPFYnIkvhB8G57BZZtu
KHY9LdoDCKkHEmL/8xZU4uNaCigRStAKd9PoeDvXDBXv5lAf769wyKovK9y00fk7o4dTWdUD5keM
yXXVoflgzVacy2RNhkdEvaITWxPeuOOeNUfjmeerhgMw5IkAptNID7YJ2FL6+nMYRDi1RTwriRYF
SSgPwyBZYPnlUIDTjxXq5+B/jroOxL7edoMLEaiZWAC/m2T5ZJamxUrnGEcxneChplnmCgAtjnDO
lDkX6wKAOW2Af4B0VcT+/df8T+Ear7o5x9bIOp8C0ugBb6UgJH9BLAGaa2Jc1kOAcjUkzLavqJhj
5GGMBGDOhTtN0Mk/V9VQTHJCPlkgdQkQTuK7biltxIhjIQm5sz0s50kh0fi6u02hTK6WsE48Fhnc
MAsryW8IUFS4wSCoeZ/Yfj/Ay45KG1xKdrjLco4zOOFKBW07tIfpb67g7FXGPHXGWkZ4TxKfJDr5
1aaY0hzt+JVcpJE1BRLi2kt9PAR2zZpxAMdHtC+kQn/VygaI35hErtt/afYU83sXwuURilIgL8yj
eBUTB4M6O65JkcJZQK2KVnjmiRBTs7s2V/gpGX9HsPo2nzUU6c5DK95EOjXiJ6rwusVw5oT7uHsX
Zi/F6Gmt2im+bnWSO+0UHxnpnNmgwa91AdKWAZEi1YYHXoYHt2AYRpptCi5Rh8Y2xmacauDCc/08
osSVq2lUGPMqfF8iTXtjuef3NBNQ+cx76/4/H+BsF/CnL45fCvMxIth49rScHADHeG+0g5HiPFgi
e++FMwTri8hhDxQGkH/WuinBBt4rzeEMMLcA9tCF3uV0tP92uVZM6hn42otzckK+z+k10AuCXTce
Yt+KngZgP0Xd67STKiObFjrb+jA8bK9Zpmzf8T+hqh+hmBffcYYqQlUx+s7gEj3Bc5rCiRk9r2dk
c++DR1vPXTnyc9HjyoLIxmHZehuar1jiCt+htkDERQKCZSRuXLOr7rexiAOXtAVVt8v1mgFhD94p
fsIB3Km9b3hULRwTJLyzm7WM5twWDy2gPkJT6VkRZkyzJ7BenZ1kKNpaTqvTAuKU1Ezr/qUxq2gy
9YoPlJlqi9gb8Ajx8pjG23z2Wi7tYn8AjLxwUeOVSedd1qriR+pA1eEEnIESeAsCnVL7CPNoHN54
ojAWiVKXWwc3s9V3BaNEhxij9nTiZiv815XA01Ws3Ez+zRPh4CLOmYXhvXVMGlfKGk1Poi6cfhZp
qsHEO7oCXfi5aC7N+yI36acKgFP1oGbay116fX88nQy1clSNX9fnL7jWOeF/993m749lyH90VGi+
P4nSonRXhBmUrKIt/i5QCbrpr6SvZIwqSWQibDb5IhbdoxhTi035urIb03eUYoDN3037/Ao/gc/K
N1T5c7o/alPT8G/WrhrakBRc6HdQWXtxbKSNtHiEJs/3ANn9BP4UFW7kqlOATEfaqZtoE2YF0bsh
8JmAwwll0TjNDO8r3E1TFUQ2T6EBNVsu7/KJYUHWbBbYTP0ZING56ecFf8Z0gjZGjQlCFr54xU6I
YHljiloNMd4t5D376cxVqEdTmn1+/oRJ26FCDgIn7QDbZuxcNyBy5xLVfv4tNcCuU87d/lsrSZAQ
RpcpFNGO7cWes9X6qEhxMvMsEfz0hFt4zTvwwZkZwWDs4buFghw77d2LBwCihMUmalZRg8xWj/eZ
pRIrizwotBDse9nuN9H3xDL35OjTMrAcuKe6W9F5cSlFMeUdcnArZuRF/gomb12yJEwBbHa4d6sI
fhOvhPBtOayV8tTYFHzvv54WUCVi74wf7Ng01B/8ho9EsPxCyTnM8iZ7UiilZniWq5AKxMQfE+P6
8FwXKWVmZQDpfLES9FFnRvEn2zrV0uQg4oO//fmn6xuc99xIWml/rGvGIvwcDow+hL47jWh1G5ws
qlyUUM+zb+g0zeQ6tWAAvQZ09yuuB3cqt/ZeZlKAaGvIaeJiRsp5hLjRuIJQVOqc01QDoT1QDhJd
ZxgfSeWGJ0ZFy9bEdKPPBymcjjoImXNgFUMmmOdnHcO57M6BJomA/xEUROHy3Y3PZipGw3GXOFzs
BslNffwyr3RK09vlHGQwMyXknPZVDlsFkpluamUmMNTXEAsJ/+XIz5a8KUiXSetpsi0oxX2ymHhU
mYGXRtMdEzUbojpvYLDaAmyI6/jZdU2YUTRGGsppE57ZFl6xVZPyqFPhUAg4u5OLb0Xgocr4EJyV
IRJ7o3jH/Xw7wYlkdSrq2FgGoftKbHe3HT5FIEN1XAAnp97EKPdYXCG0J/CCZlP/JD7aCzGG8NJ9
fQLDYOmqjAAdeIUKPKuM9Hio/FCkj49ozyOQyfJD5urufzVUg2XE6bz3+CLdiBZyLnT/gdWCfxvg
n1o8KEtLo7yINLFs6+ejUsqu2puAd0L5/MPwB2JOT2Um1HW5H54Xp5P9Hlsp5J5AT6qRNKFSXL/I
Aqh82q2PlZ9yqAdRAFVxJR4F7yjefTdB7CmOWkEpnz+zhpIUcVPXyyz3+QkiSm7TJTYVBWGKpjwv
LQ3d7HeBiIyUGWVp8GEt2kf6PPJ/qjZ9+Y2zMfUvYrUHXUhggG6Dk6cvVmJo2/4hv1jVnCiEWWxh
9h7SwS5OagF7cpYoKzQN6ADjJpAJqImcQecMr0LdcyCU2RTWVB6FUf+dOACcpQ4xbS2af//Ch9vd
x5rvUJGNUYhIXDnXfz1ABPMRh136c3TqsooW8y61do2h6ouH6QmEpnWUNWXLOBMXCfsFFvTX4gch
uoOi1GHWISbzuUaS24vMHdcnVYp3pCFSL8h86IWdXOmrRkpJLoTYzT5t44rVdl/duHuYnodxbVWP
gGH4vuQYej+kghDRfO6D0aPhHC+TDV3+kmmbdajEzymoL5jVCVBYbysUYKp/8TbHqBe1Q88KyykM
MbrJtCKYrrpq3amnOPe7FAig4hIuQxtYOHApZ++T3/lixnVBRRnFxiuQjo9zbhS8tIFQ4WQ0ci70
BX6ac8snHDpBLIXP3qBRxEPoPXFyWLiaWOzziEwe2WegTqQC5uytPXLZqT0e43lg8hIbukQNuPHr
8HgkediIeAV7JX5yLAv4p2AC7IfsaVT+u97S9EOtOsjPLg4lDbCF9yDcTYPXYA49DwpLSq1ZD8hN
H0qxcZs1CgrXeJ5h6sW5PycIPKcO/mNOCzTV+oiTuCv5b2Myh6wtR6+LSV1waI8wkDNCev+lKUBB
IEKplxUwKvK2/aLsA+iDS5DYpgYn8Ah1pn/Fw7vgOnM08sDfOf5P/gqADgB7Nl4/Yd0w2hefLkZl
q4yuEVvRFZpXqv0rb8DT27+tHYyCoqW7ckT+cLZf3MIC0gt61ff/vHx5DDYHnT9Mbmfjh1I4IEwL
dXnfJUTVMvwm2jpl48iq/iRgILUJyiqxpal/T9QSn5t3JbpOLlyOvpnXxonRO7OxrGTSPxImJoui
GuVZmyluknZNlgEdSQ4QQIyoV1+ddTwQQOHK2RYAShtSwpXrhdcsgfqSQ6+oQ5EcizAq0qN2SJNA
C0TSTzoKFkumxQr9E2mkU9ZmHOc1q3MurvMTXHm7wBaaRPFbBQWsRYDYsw3DTYUDmUnjTlsA1tld
ic+wM1lZgtN5DxJCY6g6TxtB9aItlNOjaWVJ17UNQSQBdtRQlwVCm3bUYM8YQYYbtL7KJlw3EFGq
7fJ6WgqkjKQTEA/CQYK6Oob46bGol1hFjk2c65qVJvkP59wHnixc01HPV8l5DZlaXdGljo0YgJVj
OEb/6s6AiYUCXLTr6lh+wVowse0HvVMBQkkmL2wN/bfMp1aOM8ygIN8sxfU3Asso22ddxGZlOqAV
Jsbz2OsZXY+lQ7RCePrhbkq1noYYoXQU5GihOepOAUeafqcg4+X0VYU7kwyHRDspNbKz8+bq1ZMg
mLDG3pzKcXUoQ/gjB+LPR+F6kgSxKyDqu4tR9rJ1z1tcG+tqqVcOM8pF4xRsrlaQ+45UZDHutAwB
PTQfeHinnQAl5kWkPvB5KH5md4HnLZo/j3h0/NNNwjyzx0KmWgQQpTl4oAsh4Zg9CTb1RxLdR0U5
uZ2Qxxs3hY9ms6zozk4uvDlcjeWdSC40cuj56GyilSkcUurjNyrfc7Z/Od7uTLL68Nu0Qg9NNnLr
AghdSp3JLzjT4zhfRwSkwrgvflonxhmMUFUys7/PWIpAcXGiIdbuf7gOT8a0wSFv00Ul2VxGNUIH
jP9EtsZ8IP5cUB3hZFS1a1yLEgewX+oSkQoT2sk83QtMCy/LmYjqSiJCyfi0pite91rXPYFOn46q
Raq00c3selmuK7QgM/M8dP+it6GWX7ai9Z6YbW3zQOjDekSgZgYtGoQHVeFYapGWw0oUjT38L+ta
lC86eEoEd9gS5nWaQ2l2Hcy2ZtFhIVocf5AW1ZxpMA5lNNyJMi48VrpaRxY/NAu/uThJsn+DxxC6
lx+sb6t/hiH2V8ZB4z0zLxWY6t/OpdlMyQf49cDMpGJ89ZqIKcbG1htTjDhK01SR0qleNubppdKC
be6APxP3nnAfEbkbng6+CuXfqsXfEDQInxgJl27WTDrk3SQiRbGAyniBDfh0QveGaoR8pjGOi0CV
Y4vGbSjKTFkHJ98rVrcfjebkZxybLFmcc7APluWM+sf0cIorXVQO4FV7sq3npMF71vg+QF1FwRFE
TX9nyZAkBBFiURIjw61K7gyuNMM909DU1xWmdDGQ7VKCgiSwL9lpRmbY00iED+Mi3z4Aqk52a5S4
21QERinIKMNru2CpwK0BkcMhMVTlNGHx9BXvJXr3SgqQ63LnESoKjQqLIFC1IZ/JPrc6fjN5JV1d
2RnxwzuJKyVfX1B5tHKfYYYaWJKQv2ygJLzc977d5G+ViqpW5jstria6hD0g034clevXAqf2MZkr
DrcTcASnD8xCqNJ+KDErmBszMRk7GOG/BfyGwobuF4NgYCzEj4tbxzxaABdzt0XUo/9G9MqEg7lD
H4xR6HmziAwOI6fbUNXtcD+ZfGPai0EACT0iWTPp84DMIQ6ZIeHbVH1LoPf6KicvoZ85rhmyMcIc
goq5+rxYKE1mvFMNjOPNnmgwgrCZC9TnG8JOLUhnvD8ARZsu9WW17YT42Si4drO5pgU2lFJzGoIl
RKmREkn15zqfWSDO6tcNGnVo/w0gDNBl2xINPEYrIc2wLIPGQnaAoM5yQSlNsTKBefnv1SVy+DFs
lW15+HSqnLDs0XjbcEMvCQnWn7MkEkBln472FefT7iVaOSgHSPjo/Z3Y9/2G6CzrNyVf9TwGgma7
P3UVQDc2g/a/6ljnetotxDNOR3NrzwDqll37H6IeQdYsX6+tXftwTlxGNSszrxzyIlCcLagrHzpm
SYsb2ZzlD2z2CSje/6biBHnbzQ9utiHa0mveecqrHBumrf8dUgak80uoumoACJSQAHyxaZ9M2OCd
hz+t/fIAcEMjhgXKuv+Oaop23UQNLI7onUmXReOCWe4AFUIwiVC3ZU2zFvwEfEDsz8yav0WbHe58
GHfO1MgKmL1/rrCyIrTJeXBxDUIQIv1SFzmuyry/ClrFEKxQpmdqhYVg7sVoSYs8MvM1hwtgs+dO
2dpNEXbbysBL/0S6iWpRBZsNrYz4afmcoVdL6xZ9l3VRU4kpMYIL9RQ6Q0WJID/rjHqO3Zgq2dJZ
53D+E0AHObmxGlpwiCjKiUMKcXn0LSK91L9IxEB/1zHz96MwZZdTnhadx2+6k9jreyyc0WX/bbUQ
zw4fTTsl4HokTVCY/hlMycJsYiJkfIIQ7zFdSFuifnxP61RBtBK7a7hx0Fo9aRVPZjtp3Dp9k8bP
VDi9uE3iXXBC5ftTgBC1VhLj1EyCcW9HvGCy2oesCmUG8E57rf1wucFprZz6bgiF9AYYn6yktwgI
kplMefe+sC/d9fKURs/Hu+qrEEWsLjI4RSzRsK36qAkQ4x0Ril2SEaK2jbxQ+aJFCcZT0QDVJFGK
SciWpRp+FijO8tF2w8eSWR48PC4N5SRz+e2mB4B/ED1SLculVFkCZ/hQjYjMpKZnIqC2Ac5fVKiv
oJPKrTuJKb6XCJVkMh0HK8N9ukKmS30ajQNid+YYjCSAWdXSxDwqhNAgq2RNmNWXsXgAfiNgAmF+
xNHoSh1ndDcCUMyRkfKTKnRmMEyxhIWtnMfirpA5IcmcTKgCzyN3lKV//Mv9RvwKHSVRedOxM3B4
eL4jEd79qTdsRDqmleRncFmJHDMIJaQ7jQRpax9lWPjbscfg//RRA5fXAimvvNzBZthrGJIxjRnV
F+27/dQmvMQ81qLeASPnb6y3OlTF293tEGXxV2XJpifr7NNo4oefby7k+H75pIAgqps9/UuwnwN0
dWrgRg8ugTVG0TNzYR/IF2H3Jpz51WLlWJtWy6mE9owbGChGKKVFIAvlM5VSFVng45jibO5wW8RY
rgrKw7VZUasqHrGik8Tb93QZ/kxd4Rz0YgkYO6yn5XNml0F3JrkvUNvcZRYga/2RkIniXF7tPxdL
cq5lAoi6jE4O/x0ws0IN3dp86eTEbNeqIe0U8Tbi9GTpxQYTmzbO6NiYbu5EI/nJcF+YQOSrjYt2
Ipvlpbpw9SHCSFEvDhef/IvtChmlr5jvZHss6Z8yeAx7UoI+/Gs0ff/tonDxPVJWvIetrA24tIFn
eqIAc/rIhbE0WIONrkL5J6CFR9UZ8OrQThsAJnnJ3TDnaoXcBGbORcl4YGzblJg3U2i/FidvTz6k
ciJ8E+HibhtWMWYVYeMs2RW+CoasqH51om1wj8LttSmLb5vIZkcwquxT3V+pmBwy4H3RSlOJL7Mi
WC/f/17bJJTDDXB3/r+M9eeAPHqa41JT4UyCKi6Lfjr560RLorU62l/m0A0fjkOHuaWL8V6vEFjW
30klefRNQ80NjTDefr+SvOaCcnz+1GHsRxWTxzTr6nIJY7wS/Z77bbMZLXUWbj7INz6amDGnqrzS
EBwCWvGAyaHZykf4S+3V44ZR6OvCsyFxO0XIUW9Jfz5JgsOA2tTSXjnBi4Ow2vv2ME6EEn23EDAf
+0ZmUGbNLMqNVRp89yxEzJUIOM9sCiaO532KXOB7AqDiL6wJCBMT5rddlW60S3J+Grq8tJnnz2YJ
KK/IrPTgeSEECIbHSp8yBTYPq58qz+LC78kGfk5V8sA6cMcgug4nshG4Pk7lNHNmQjdEBJ+Rs6eJ
rQvrdaGXKEDmkrzPfIb3bu0xBOwU6rumtun8seBtTE8OflHaqzAPrqBbpIoMK8ALFY9spDIoTfba
kfMf7kwkTGiUnB+h//gCIenwYKgTRDFTyAo0P8hqVuMiHxmNdJpZQaBkSnxHSeOwGd++y1/6GVct
uMUOn5yF09rCt3uWi545C9WvF83CCl6dTOAw5uQVPTiZyQFLmLLt6Si4ykkzBfrYyLIEJNTkFlul
mHfGJyAaW5bTzGMO8ajxvEGfFa7Ql+kTFIwem4a6Epv4VxyxT3Sd7R/v+mGkH5jPzqMVP+Odu/Wm
tfIZ9zySDPImdUpnLaL+QzLbHQU8RgqETGG5yWt7m0zORrNjzR73W+AqZAEoUe5LOk8TSwcLXRpq
haGq1biUl0gE6UgYVDlGT04LUJ+eVpPdckqBqqNvQl3tyDfPgnYz7BiV1uRcSd/zqNCtdYy8pc+v
6NG7JMZLftSEdsm0XhrvXFFL26WU+XaJNEBS616dfaghyOusCEnMY2onQCIFYbt/7bMGIPzk9c0G
bVUdTqQS+ojt1YnGf3IyfRB+Txvds/WfOOOux8XiZ6XiriN1FAMxBwpIO2mjYFzM5acX0B47rCPf
2FHGSjDy39vqd3umNc+pLzP33ftF+Ah/ay0H/sv8CWmuzg2i1E3Krbgvcmrvu1JSiBwDm/jv5Mln
E6pH1ChJNCn/UMxDizza/KDeOXhTPHtGp6meOvQRvtMn0j59Vy2232Mi8NH/Qj+9NCxvraOFWAtM
Y6v2tFHuNrZgAKnwvlWPQ4YmuPZ8eWQi8ehtbz9ZhoRdR6EUbiHKPTjPyEM3FbdyaI9e7xUE+rtM
RcpmOKs9/Ep4N1gfyYdcdZOsX92G0PBoqSuni35ZYn9S+8TgOQUgclOT2xJq1QEmLCpF5J0IeJ3d
sl21SL6fHvrXAw86C0MSpN3Ljz/SSGvUojqw6W80d9J29WflVBqm3bz00MrL69bYQgUEyY8mGkM5
rhvIveh/tT9iknN66ndkT1KfQhSX5BmA1oklMIP0GJrLi8NgNmm+RXrSy+iZa8+MpcYo2DUaIGWr
6igpYG73DRGWT3YHrKfBiwB9tuon0krwgPrZtyn2S0FbxU63erhhPORn9uYS9mbLdB4ZHXMORZkC
v9i3KGVZFhqQpEADxRD+jZvw14JffuZAfY7UWm2KegsTomF8NHGjp0XOh97jNbzLgvwEzSrlisMb
uiP5V0P36w7W7aSNeExs7djW8kx2KmUUJM2J623cxbazgJpBvnb2m8ZXdnl54o3CmvGlODfJ6kNW
tnBUQDar9kHI9hYgH3jwfGSaV3nn9RgdRq35XlQvSb7tS1KDD/Letg8lY2r/2sm82kai4SyyI/C5
Ns7y/JqkDaFDg0gKP8MSsyaHhdf6ilQglazG6VyAH6a1TOEBOWSGoOSz8AMnTummOrlBoJFayMof
AQTJHmw2h0mncRr+AZx8gHLT7IEZSAcepxpM+5nmq+XK1R94Lyl4yXyxW9BPxWchF1SOI5lVvyXN
WFqTRDv9xd8UXwRrfiWhDX5szQ/ydL7fgclnhlJOah8lN+bRxHtHX12USbkKUS3zL1YHxiDkwU2J
QUNiOHqI7s8Gb/SfDPJbDfU5W94g3nRI2roxxoGKwQYd/l3RINHDefNd9VGnF+r6TNe94AToFBpU
tE4LOn0ku2daM70tamsqFUHrkdPBCTJUM8kkLtx5IfrSoiqkh0LXi4SzA4dOLbojl3j6eTKsIRb/
18O09aRWLfMG4Qi34eKYaGOKf08YaargALf+Yt9jdMw8LcCbKTt94cdkw6oO2r6pCzPJhknHyeMO
YpB07fCrWLWArEK0PjDVJHx9xzysk9w9P9pczRq6nHr8p6GXt4j4xdxGj6dBPRbRGuF25aBCwJ3T
foEe6/AXf6FYli91Oo+NeyOtQ4f1QYfrJ+7+Ng9mkxywexAxgfRNhSNMQdwbMY7f+YrjfMVPsYNn
U9UAp2WZD9+riefbhcQdsZhUYJYDN8R9s5m6ffGTYj8QIb6BTZ5xG20yF5BcSWYHupqTdEePgLUu
MQmu50NbXi+ePagZhwz3Zftvtf5VtTMGJk/Ml2I2NyzrtXDPTcmwA92n4GBW/Trr7tmspqmxh+jF
c7MuSH4npok1nLhsVomX5Hs+e8eH62dE3f5vZi3QNyEt+luAV4wnUO5+p3i/Q0pf1aMhxIT6liDQ
TSozOpCmvTYMYWJD0bcTohQhAuVKyLLbv6zRS2XIis7QjfqYAxNiu3wdPmdrrwX46yFDjJvhNQ5m
Vt28EWHsdujLmA4uy35zbDl8VWAGvTF/XylveQo0cwooCwe6WZaqHvo5zcv0lzISxcrH2h+HC34N
uSolgxfag+WBFi7taO5JIHOHfzbl0K6Ne+Ey9rpzVK2mLb+oLP19tZouEjK3Rhbp8g69TGx0ozLc
k5Pfs8grHp2VRaeOgWD2y13paGJ1RxA3eIeVmHl36/bTw8IIM7eqkbvPKh1X4B9J827ImR5VSKZi
7IQ0KgruEJbRJpU8XVh+i1HqxtGQcBAIPDq45M75muEinmdRgo83b2fQR0eHHqRi07/Uj1kZnvBw
mPigp0rn7tJRu5v4pGzcW5kirc9mse7T5spY4jHrycD5aMDBjRnnBZpiWB3g2AP5i241/AnaJgWy
LecWjj+OMr+XvbsqZDjDPO3MihztVBio2P8yQ7iS5TXHIDs8fBurE2J0X6R2/2t6ARpcqbG64aX6
jotgYDxQbPcsLQEWr676guDvt08AIyRMyrFuy+ueVkQBvdoIZLwleLZSP0wZBOzlXis2qhfsmn/5
h+FS1Bz04mvN2R64hOF5sa8Qstv23pOx7OUMcLepOj3IqwMBYE6O9SJ8l+hLl6vtHukMoxfjf2eV
JyB5Tw3ToL+Ykzwv5tOJzX+3mBGXy3si/qFqjDqtXG2lab2oaY/KWRSaUPlrsQHUhySxCSO6Y8IT
1sTNkMw4vQ0RTKYgwBZyHGyBfps85jgOum2DBOGva+UEEP4XJ9bR4MMUePI0/aixWklKPudgGCFz
wiUgg6kxVs83yys8XOJt/kxF6Kf+HrtcDPACR3v3BIK0Oke1QCSJ8A0m5+6biiWQHCoj/2idgq/5
1eGEhU6lZGYBK3uoZqoyQ7veLgCrieT2AR32HQklQMCX5lb1Fs9hxOmIWCKWSbFLiAhd670rJO59
zJXJJbHzMJjV+NnMFg0rO1SXZBIF5GPZgBk+mHLoHlkY53rnEzFjXuZFi+v72mPPuaBdzUd/rXnY
Pel0eUD3zxiXZjcoHWiz5qW8iZMZvNL8fIOVQ/tqJjK0Osb4UAMPuoqvyHBfrcr5iQcvNljogaJE
IVvZEM/Ygr/haRsxAM16EndZiT7q5TxirBBv7tQXi2ZGZA2P4shkL4S7rezO3yKVZCJHd+fUNPxX
K/OW1hkxf2Djk2BW3evbN3TNnBu+mH41/XAO1pPNwGumZc5Etn/zDbcJq/UT7qlapHfGR/j6tU+2
nCQ8MySUzcqkXL53c+nTB220qySYeZGUCLbisdMluveJjWkVPXznmeFKMSVQaozdXBB2opTe+DFu
UOtfIqsmSIbyZEA5IsC526KA55rcvjzWqcsEDsvU1VwinLMg2ZjdT4fK/+Iuk14lkgyTdC1YqMvh
0lPFK6tgK+oTHZ7zDkpsmOsiRMJteEtRGAet/4iY0Rlo4Bbs4gb/EDI+DXt5g4RTY1ppDT3pPXFM
6yD0jmg8zz9SKjEv1xxrBlKcOCzKZJ1vO4PrRtgVF9INMtV9cKb9W46XZZUfFju84csM4WQfftwJ
XkY7v5hwsty3rSm7FZIM++/regcEFMSyfSMDr/6KC146sNaJnoNbtRxO8kXnj6d1bqnPZAo9LOGq
2xYhF1B2/tgnzvh8nwRL0Fb7c0zII24k4emG/Y6vO/Eq3oMD5YCvPyxPu8lVdFNmhb6WCV7sc5sv
KuCfM/Ukm4WVWTHMVnChlczBrzCwlrJ1Ut08Egrx4A9k7vI42hWqwLBW42sB9FvlqHHE+3zgoieA
/gxkON4mApyowGtCCsdGemVh2F8H/TZhmFDBFVM9ZOZwE9maoNLUghF3vrPEodPEj2v/ieMMyR0a
QbeNCWcnBLm5swaTSxT8kiCa2Y1QbFHyZw/IqkbeWvLLFwY/e8oNFsP2pQ/vXKjHyqNG0oW/pPhn
6D5dYNMiOuCzRiLkOBRniwv+eAboCdFNjdV5MrQKBllBLLIct4LmhMVo6iwCGTUDR34Y7DjS2aZN
evL87O64PclKSa2xcpY3YKyKf7+ry2deXtKWJ+XCXB85szvi9j5xNaMa2esh+R0eDhNxWDN1iMkJ
fe29viR8ofL/eYMJBYBWd1SqxCt2UmbJrRj9bjP2HmyELi2cqRP0MI4gu0zMYKyAD1rCXlA2YEG+
HHIO/KcsRZIUHCMVwi0RP/G1Qi9cLSmhJ88Hcy+Ws6Yf3Ah3+LKiJVk6T066uitxJnPrj+Litvto
SD1pYHb8d0LEmCIUsjJkVvdjDieyMsm/ZITjl70EaT116MEn4LGgaOrIJ0iFzh90IbJHXGi9jI6P
ZN/7r/8q8RzHTOAIoauOmC+D3/yw7Aa+G5ecwVLVZ34ezEkCHliYpP7CrB5LJhOyYj5omrZihhCL
69g/6/ATDS/Cq+SEIVGXysBQdsVWisdfeIl3MrlJtY6+eJbSENB65uh2LuszZ1+W6fJuoiKzw/VC
IV7dlenPphT6A5+7AZtBYzR36IKrUI5DkRGwVUPfejuRz7u6XBFwsEfki9etXcKttIxcNx7kJxi6
38f7hnVyt1aZXO0Ulvs8S6PhJMUjaXUL+yYa79Ll29s6cADDMspuP9xwcgKp4IwPKeQWQSpR6uN/
YuUtNAxps18BamioLKjw6i9Gg4RgFD1d2Z2dxumDOTZp7tElTBRidrh0PeGbOW0DpULM4XlZFvJs
/s/NCELgf9bRUq1NQ2BLDdDeCUIePwBVvyMwrcL7fUIMNgPLis1WwiB7TkdwJNnGNclDdpPsPXfn
3ng44Z2yr/+Bv49YSGny+qi+hoqSIhFZFDjLLZi70aGRHIkcx3EZ5noDNg1DzGCP/EzGnmyd7BUr
5LducCP9V/dsYFjuFBWTHclPRa3VvsUfRM3yPgDdxAbDXHGeXjCGIrpzwQ+yPE/kGkFkhwROYPzi
tAlIQT/Wtuki6ZjIEN8Z9WT1r4KpbOjyWnQ42FMz6ZK9fH9tyUP98XZsE0flJmC3LeIQIHkLIwAv
LKMSNsCD/Bi9rq/Tu51tJ3GLazIM+acGN9VWCSyYlQE1UEuDvmPS/1VTWKbRd/1yVqRYbryatIHI
HHT5sCB7YFrIi3SQFYjvlI8eJUlQUFNEwQcbayEmajT+WKQ8Y3Rcg1AKJnBd+YUnuXwbNzgt3hVY
PUWUI1rNZFIye1PQFCeNGmWIMfjlixpWLnLnSn6eqXeh+cGLRAdi+OSuwpbLUPrerJs5HrKtvZZx
sDp1P2zQW876srQUb4a9qy3qkf8nBiuVwRIe0Uzphd5Y97HMkol0crmKuWoMMADDM1+wew4McCRJ
VL3/mws22StAwTHoQ4qh2G6mXFYZbpzkMjKzihf3Z1c3s0xDNETSutz+HuzIUVQEagnNbiWxhbms
R57IkWUKGF3+EejBEEEGj422u5ClNzLysr650HUttPcMf9b4ToxP9mv2oYjIjGXVEimfp4i9uqqI
Zjq5k8BbMj76/RpWoABEtpi0uGXK3M54o5HJGxNHyLfX2yiIeNJy5a+32myf8+Ar3X0/AcD2r48f
nD+seImJn1epUUxo8p7wPXhzThmSNU25CZyfpfWbgYFmzoOY+LdkUnH+31pTI4LI25W84CqRU2DT
eK7QE3vxBDqV1mhsvFIFikk9jdvR9MQEdKIeWMkOzr/r3PAEtYGCRbAEojPqMBXpUo6g1xV5TFyG
vRTUXSEan5CY+HtiVC6gYgV/gVbf4G+Fj/XpiWlJbLjkrldnrE1HEKAbFc2b9qkFl+eoDsLntA43
wKWJOVJlzlqGToA0ycNJ83U55cQaOSdqjbX7pzCMJ+e1XBABZ2JrRE+ETcHzCHJQBVjzruplmpf9
rQKrttAQD7YOVddPzfchaUrrlSoxOFT9eTs/8hiqa6xxH4iwxza7b0Rnb3EkHvth2c2Frte5d2+k
hPhVLLsC6JPQXzUuPUdaExr3D6v+WfNnBbddISyQHGPQEiuIW4ZAXirdr4TcFDFzPS34hGuj+l8d
3pTOpBMbXQq6RCtPb9uzRb9jdgjeKSWuw72SdjXflFFIR7kXikRaIjIGis2xmhZiGfcxBFI7s1wP
u7zQrl+wC/zD9QxXAzXNjLTvdXDP1G8SXnhEfivHN2sIkldTjlbmzS/lF6N6NO6g85sg+KQ+CUk3
0I8yVfmkYyuCAImJ/UgFEKi7e9XAZyjK/7pQ8WsUzr/HvXLn6DMZVD8aP7ryZayCfcYp5zPBB4dW
hyUxYPJQImfMVc5fm4+wBMpF+zFn9oyThlGt+08TPUrd2TVX2SXb5LgE52fEICSGgMeltb91U1D8
GaWbofhD77OwKIbrspqtBfXBiCSH+FLf31Dy3LFfNJTbsluOMaJB7IBYmQ0lLtOqd/eATTnxcMu+
JeVESsa9eBwxBOI2xtiJ/0aCAR3Inwncm7Hd51yRvC8tWI4TgbrN+AJMZJeCjKM6Z8/4xdWIGKFs
uGETtKB1DDr2ew87mCJoiMUHJhZn2Q+LSTl52NH8nRAnlswjPiSn6bXG/bmjPmoed7oJq0WWJ9v/
1YcbaWuogIsISwY7qq7UnA2HFS1OMbKEL0nBNAqHU1/aYrQFdyQFQHZT7vG4oviQG6E0ie6zQYfR
WXh0vNhIrcn0cx1Ufx87+D78gFcCISPiDttPG4gIov2rfCioCgQGDXD7yKkbPT5ixDRnNNg42b4p
GsVLN65FLe14rShaMs/mi6aXT6fi65N7/CFR4nREUxwQQ+eySTEGUeGmOMNh7N5K6aboO019liN4
tQpHex2k1t2j53VMxvWMniW9Li/WtNuPXmvuYkpmFdXUEolexavvm/APMNxM3hnbpR8dglsp2ELm
M6O1afm+j1icX+zu9w9eGo4Z5lin7V4UmhDCN7vXROXSYG+vZY3OIsN8SrUh4fvqci8zYf37lgg6
Dfa8VgfVfENGp/Y+NrHrslPVRyrMOpnU29bsNFzJ3MCeojHYpcOz97iz1vmyukemQq2xo6qoiZ31
UYUgo4vInC9jH5IrQSt0TbhGAkZDoz8MxrJevowWDFQl/hfAJVlAz19kFfuBH/4RDtAauSXeOD4C
a31ZlCzBAeb+UHVzE2DuH3qTBuVTvjJ1B1h8JsXq6lZlHNywmSjCnOdqpJ5vz0ZzmHbJJAvc/fIH
2YSaBalXtAas/EpafCwHdukCrLgi1V+TkCPPIsClSkhxlhUAFdywQ1CNTYydRJOavRbOP0jL81mG
cZifZgh0t2DK7gnCTzxijwIPA4LcuYJpwwkQK/2XZQH1OP/TLhruUF2eSRvaaLFesKk+ocCBNOXe
tFD8HqNYRiMDm07P9U5eM0xXq9WMeE2br4yzX8YI2M5aZZSD2tPFeRNEJDq/2llyHG8RtGHgK2DS
SV1/us1017ZgcjA+i6pzHt0vMBFSORt9ntpbppnOm4AndHJsd1kAQy1SasT6vKtJdb8WmvmJlAAr
XB3p0W9ED8h+0W25Iz1djHwf4iP/hotPI8berdl8zY/E9Wj3a+zEwtacpfxFpMtS4/N1R2k5465O
MX7D+EmA1LP3Ppl0Esw12QVzYtgXc8HR3uYHqvprmCm/M9Sei+JxlSvn22qR0+08xVp8hoMzirvi
PbSd7Ca/rwJZQv2zv81PHzlVTngjN2+UKQJNGpe1QI6t8GPp0ZY4C2Xh4Jg/QqTN+/bsWsbvhB1U
Jmp8bXyYarxkxHg9brj6oIc38SCt10+CYIP4CPJbVd/W0a6Z8JFLfW8GtXfDfguj516lKR/qrG5M
9vmjIZFYOTkf7oIRwUbUU70RRamEIQoSkHFEpbLk8qShYKTfjPFg4puu1G6EUmhU4QtTQZ7uxapF
xOQLM1RzXCN1f/a3nY5hby0Bi2+R4fshywgvlMgSWGx1j2tYWb5wICzCnCW4twdghoejWi36hKmW
MoOK6qE2iGKy2qmn9i6XJwleMU+0ue0C6ip7ZypSu4Rjx72KmygbfgSfGY6g+HDVpFnkQTCUHBU7
ZohCJr/phggtPOSRxMFzhb1bXD7m+zFAbaa7ltYO2OfBb5RvUzWXj2Pi1zI5QSeDY5C+BjLGoiBr
CLTU/7pPkVzZPkwb5LeWIR5G/qiPqfjKx4JNT1V57SqZA++aC37Z3L/1TIrxZpkMZSUwliAxcfpH
tXQcUfN4cY10hLjlz5dEGGRrM12Kil6IRAESAxy5zp0RFWELa/xY+MDYdyAjAtpFE6QYtejt9hfr
23wrPmeRZp+8UyM3D9JbVvurwwpz3n8qte8ArbBca1NWPVoLq4pLH4yF3+lnB/JdgNMvuDfzqow2
OLdCE4wRNqUJJ5Ahq1XSkMY+PU+WOKwXqQjClFt9KFD4SLFNJqHwOeaHZMwGRZ5o682h4WNTIOl8
5TgxYXPjkcPBghjWbp37IyV4P1/aMmgrGVmABO8KKr1pSoAySWek7gYFqPmXVX5TL44kqI6/C4dy
xUwjzhoaSmQDw7juVCix0h0LNH4y35vk2cK4xODjX7bdzP/pcHJ5KJAf6P6uhH5rnt/bRg5YEGqZ
G3yRv/WcNhIj5V/wjJl7FP518pZd0FRdJ0YUzOAwX4iTYtHpraIzPuptdXBRGpZ8TpzHCHU2qy6g
cHjknk6braEZa2eGk4BC/zimIp4c3NvPwCewn44mj0if+wX0/CRz3K4hLsC87HxeoLf7VPcBhayV
TnrAB6kmDNYE892B8xuG7WiXAwHve9Ne5+2WC20mmrc8a9N9quIHof3DmdQDtBrtjHT9iJxBr7jG
28ijk9VwkxuaWRJXtA31rWAPUpkEwsyZQxjwBwtuqQzf8Hq84DBD1WumLRVwFWMcwASUaof6nZWj
F4lSaxc5KqEWX0cK6a3/tvZpKU0D99ROIBIiwc3HQZTmCQVsjmZ5lS3nP33ewL+lqK8D92HKU6Rm
zsLJD5o0PRxVdwFlZTp2Zs1zgBFmrPDmQS/84SQrx2/NOr5fVSIZKkD3vEJRRE9eexsYR635yFkJ
05JJkQBbzifldNnM/nhn01Hy8lm8VvyYmV74LIpnIZap43XPHj1XMVa5cwUyvFoORNlK3MLNhFzM
mCjVQ2LiidPOq4R8bhIv0byt8h8IfVCXHLP4QPk2KGqJMkXTAc1MqtnNqyPO6wDln7NYiLiN0Fhr
Pqc1P+oe1P54SFare6lHuC98d8nfczIeiDS6heE63HLoC1hbRQVwtbdmiqUDsVgjsIOeCdCgZEE8
gFpaR84frHX8LxEeWK14T+TsE85hyOiMBjI7wdmI6ZaZVuBuXrFXSOM7uuLKJ+l1EDHUFXlai5Qk
7T041ntrsRNGdbXc6LpdZeMxeg2WcevFKHMkOfpgSHyJFgABxyoMeE16d1mWKf6M+vC3cGvceA0G
k0ckpjSVnwO70zz+BvPOxUOCmNeS2EgyqMbgpUGxLfczpJt7Yfs0l3ehlfdBAZOpLFOjGnd/OLlI
dRk3G83CRgnbSmNVuHv4hJtZ/HMlcam5Ib8fBxZYftDUiKZBr+w508YSK7rVSvvmzxUl4FNg17Wm
esrZT5r+btCpvv+yHwmvP9rep8cYR0aCt57eETByVG9zHcI5tL3gmBdCEVtIQGvc3pth8tQllY/J
57mYJt0m76/TWpi6zC70Z8AhdoZPYHRlxe0rSDFaanoOcfiOElYyVtGzQwt5LtumIZp2F4Tu44Xb
jUNXFehSXK98TySe8uhVBvKhatGOxns6RiThR/CIGutD8WamnSAGOr8TlcWeL7Jcgdr42OtoUaxm
RJpgi1jJwmCZD5pbilTKe6XSikD6LicooOrhsCvp69vBEY9QM2r2CZ7+z0zV/GPYqPb8o/J1iuTQ
vLVUcadeycTKD+qM8ARL0QTqaLBUgmVtycMSCSAm16Rn+A9GzZvb0Ge85DpeLtoLFE5QixQ4DK29
gU36H/uF0BGpQczGUFXZcMIzWTYUtJsTqyMVFMYegWhMNJmT5pFjlxpNdEg7k0VX1t2gI2+1KywW
8SRu9gO3rY5zGAbnNshhu2A7BoofTVd1o0P87v8Drw9yyZPF07Szizl9AzEOMNJEY0p4SPizMlqC
yXbxJ7cquBtp32/9OvheeCpk5x+iEHEdt8NMvT3EqcuINUaS007/JjGPFB7o9qZVxdDZsOqoBWMV
WmqMMpgKM/BCcw6Vw4+Yc34J/IG8GPCdSHdtN4LW8FCdFN2Xh2WLbJLyOyPooJweOSWtUL6G8kx+
z5S9t2IbN3lljFRAp9h06kOKMy9bF6dQFVxdgg0T7NUtzSt8LYBi9cwRQhD8XTmruTFNSlc1mMMy
7rvBSUNLaafuMQsgWOgREnNl7pfMBfpYL3uq84GbM4Iup8TgFT1CyLyfN6bceb+8WU5oLY97vCw2
NMIRLeS8ud3Gm8W7D5FSrgnEoKtYRmd2JuLna/FsuzG+S5+Fl4UmQU2vrBJHVhdanhCW8VD8OLNm
k1TwIAGS683fWZRMHQFWIxuvNfqIaQ1OqFwoF8tQOJVod+LODOuh/1n6jjl5steUilBsDtd2lUit
YtLyQnbnYFdLULhX9n2b6AJn2w8OQpToeTJdjH22l3U2kbUqHMwz//+bz6wtDj5d4HoL05HoWW27
a3cnan19ooifiH7b6uOSjvRH9AyaoohJwhNo4Vm6f84WvvRkxxI878tPzOz38dU83qHcbK39hEts
MdgNxNNSrEdrO3L57E3yEPrSUFRlxfY3Ryu8ijsujsgMNWInBIuka1A4f8mLH8TNvs4akjVpoSDv
wXzeOukcvIp0O3V/+0C5E97FStbAPVqP/Hc4kmmRvD1b9Fa1WD4NIwn3E17vs24bqYrvDcbvjLXR
bbQruXf0a+rNl2L3r6asL70F2B6/iX9SOXVGCsER+ruCrQ4lX3qd2kyIlys0SkUlrGcA4HX91YRI
VbWMIFUTC1aaqU4mDdHH506duOelAfhbHjdbl9OU5zOqEfh//tdEz64anEtoO4u/fWbE7TVN58IH
9ndUlFaijViPmUzOyfxlWJZTQSEEwer7bgeyYE65pUOU/T9W/soxs4Adkk1kZ2Pk06eoHWUu1N5y
wP06+e3jG8A3N0YnlkPnVPAZXS3WGyZhjdBev0Rr2L/Px74RwJ3WuSpV5QvsMJjYbP5SXDVzC0kO
I4p1B2/fW3hGVlCfjlK3z5up84D22TAKrlxfJhWAz9qmEcbYfrvNLJ+XIVCglnqB6dY+9WkMLqZJ
+/FLl9zLRoT7ooVf2mR5m5kvTIUaDQmKbwIviA5Zn2t01e8q9b+zCnLPS0qfmfWLjlHnfLivrEfp
Qsbn1AS8u5+giFNcAROkEJagvDvyKUQbUv8LOpAv0XvcQ99eKLN0dYyuxZ+hpeJqBFVolWBqjo1e
6MiMaAiNhMm8iUi3WqRO5IZX6bHpM+GcH2CM9erdSUdnbcl2zQzsZ+m56630a78uSOw8YXVZkBfr
62gdOGvQ13fzpywv40Bvo/kmG6EOxqdwNJI82Qi5IjpTFxp5+kYEr4Dm96djrWOHpPGdBueE4YN0
JS0+c3WIeU2RmAJAx2wa/Fg2/le7fABXgVZY9qnxAWM9unWpsv/ggJ9Y7oOAJxHfZ6J7I/dQF5EK
PiBSWtRcVLlwetmACXAwaZxBL56m0Kp1ayiCCdyQETJFjgKyNXJPHn/tOoitxc34PA6UnfkdPK5L
9sudjlWE0kH8ITAHD8Fe9haMWrv0r28EU9lHd6Tz8rGeSRleBXZQ6HJQc1ZkwfQBfj2KlPP9zcg7
JdgtcSWSpjCnj2OwjbypEHLIfYtSkPOmQLySPuG0i7vzk7zKPp3wVbwMeCtA8Ftd27IRClIRybjq
OVmpva2vPGbDGlFYsmyX/60U3MDVkXgecYDHgsB9t7oPDDoH8PW2bc3sVwvZZMT2EkBp0KbO739o
dS+Bf+8lS5vS523jupBwd5I9kOGVP9kzWaNUtebSeLFXQhfSWT9vxy3qFSNwQFio6sthSd1Ui1FW
irhbOBFHUQLXnurK9NYEo0a1acl5Jq7kzj4djJ5bSnmod7u5SPvFcTAYrC8Xhm2ghj9evf9HZQM1
ctOYBmns7zoDE2GcccUzlygoQyRQ6prBrFmBsa/ygSMGxzZbOuF1UTVnB8WJr390NcA6wbwC1Jc0
97bQimQdmBfK+b/kXlhxInblyG3TccEJ3MJWDFn63lnmut7IyA4s9oAkC/zcmt4ItWNOlsdZ4WrD
UeYY34ORoMYT/G3u8DuOu4j4bMAxR2Cc/TNbNbXup51CsqbOZ3Y4tHjt5uL5ecySb6dpB2LfmtgU
xZn7NtKB8sSS9B+lq6vH6/rpfeaOy5NZacX6HjY4C13OuyYfd7kQfuZn1MNFo6+vRgznzocbaW3K
d2BRs2si7TigXVC7LveDWa/aVILip/TtOjmzyGnsXNWAXZPDVB8qg/WNQo6mrzBoJ+F6MXk1mwlc
w4QlQO7rr6omCZL/pYuF035e863oPBRr8tG7LKqweMMrmFlCXL+WD2duRQJdS0AGxPBliuvJp+Iy
KUUJHKrG8g8Z8F4zWnfikwIYq3Fqzf5f0CN4Q9+o9Q7h28wZXwnfUEn5LirorY5qnB1mdCJKWGb/
kBxJma5QSnKSThA9kyC4fGfRW56ZyvOJPsbrwXA6kbqsvtotRa5snz9ljtv56A1aJpzNoO4Rp4zy
9X6sIcpcKK5b7kbOagL5FMdBVlfqBdCjU0T1QVqSQhoK1rMh+i7VvPF+Udx76rUBHbjh0Fu5U54V
HwWve8C+a9U/SqXqtDR8WK9OncEEriFfoYz5GCognbstMi1GAG6w/0Vx7paq4KVzlTTIMtWqnDNU
VjsNtDWxDCXZDroZh03HnqzQeCAVFz2oHVq6RxQkUenZJkCiuXQQPfTEaNw0ZGqQaPF7jXq368Nw
h2HU95Qvit2ofZ6BkJJCNF/h+diTvZVNiRBIZmFNLTxhdHTcwuCSubWTnG8rEnQo2jnXMBTWGRmf
AbgBP2b5JH7sihd7H/vmJZSIG9ZrXjoDoX/9wVQkBfUxOEXubh4FW5ppirfmDci4A3hcuCinlYHY
YW+45Hfy4y+PlIVheCdevki9Fsa5AQn/56GXAUTJs1h0cX+f6Lq4+XLIU+7p+z6IXAANI9tBg1MW
fCVdfEFyx7KaeiuIvucqASd/qjAJJvlxjm4tTqcgqLZEELqGNXAElgNtpaZKNAjAqtNGpbHBfvRl
VdpFGqmi6KqX3O1oWfHhdLwkpzbyAIh1425OQ4Uws37kNpqa3VxZFHetF01BegCC+K9hhMO9fVPI
Kmc0kKTpXhIdajrV+/rBP13Y/JUMaGF4bLQCWX95PBqdyW/8DgrMIh7+//TyeIjVdf74Y2ukzBU9
/zRBnjhNhsCs1C9YUKOitgCdFbTBJweJMRMIUdc8zKZ2n3d8cIskhmcsn8MDg8dz/p6xfQDLfsjn
gfhjZSf7Ag37th82Si+VFMLlJq/JPigr+0t6A+OGKX0N7CuoxyGpVxPou040YKkRRF3wnd6s/Vek
T43GfBIUEF9CsSnLUmzDK3Ih4kJWH1+QZw49eJOH8+ghUtsegl5brRxDsL5AlLpImrtJu8gG9B3Z
eqYgepmEbcEobCGCQB8DFyI8Du0qusJ10VjigJlIDp9U/5UhFusPFsMFHbbJ37inSqQcnPgixYi4
eg1cGzOym2O87/oMpcuRuxpI3zZ7Usu75ehmSH96LuCGEQshvjTUKFAuLJWu6ChEEiXvt79pkWap
dwrlVXpTBASAA2of7/+ZEVM/ux7t3ni3d+Rw3GFsPIwQYooJpuh6SKgSNvx776a6Jj1/eS+KNQBs
S+MD32gX0i6SoRbEHtEq9rPk1nOf+5wkVIYgDm/rAi+qPIvRTHzAO3fG35gzqupko05Q9rMiF8Cb
TzyBKB43s250nZHYCHzDKbFkEUecaBE7XkyBOnfjgxZDxqToYemUZxwp4jtUC7bgX6DdOkOINmQ7
7shfoiz9yl+QN8y32Z2ZTaKhuQVC54w8swptrJg+Zz9f6JWFU++huUxPu17WkGYSLcpkwfHpkYLa
6TZF2GSBeEiEJKWNK3+AcsB6QI67u6923p1hSYwP1AXhvUG/0OdWcpsBZ6p7Tn0loOWfYKtmZKJk
gzPaJb4sLO13SjG1ck4FZ4+jpcV7vUeAfJJqAeWcl/GluumbgNqC2B+4bUZnFFbNbCZiJhEWllYK
BTFgeNANzlTVzLTyu3O247WF++gSGORaHHX6OhgYPWnSB5UJXMHwzVj7lctDKHD+xVX7JzAJUfQG
HJwJdBRp9A28sv6FkQXNebKKokMYr4CUUd6I1WX6irh0rYMCJqQEPHuu3D+1QzfdDzbNG+SNrQ8d
/5zpntvX3wrccjwlO8g9GIcU3Ph6DsJaTp52eUi2ngbi80VdYyEesdVjjkeiWvlgWTGNq8Lx71ql
be8NuCKrH7oqu4IVplb+6PLQEHxbOR0A/khPAy+LdvpjwER6V63iQ3OG/lJU+L6SjdghwZytu3xw
0MJDYwKHmR9aynf4bQwcTcay1NHmOWFWeldz3I6HKwmUiOkIMECGtk7vwVOpxja2Zh26jLzy5I3q
A+NlRABuMxfBKp6eKhv4A+71LD6EmCTAt84r6I7+3hYxtX4IGgKjqbxlgLwtPsQhlZtBRO19Z9h/
9D/2VKKw2kt/oGkFZmgH83gmOhuWWEO8MA852WS1QBVl9MkdjJ/NPOB8ENBfOsRRdXptCxY08mTn
gdDPZgZKwJJEezxfdV7UcuXs8y6CoW4S6QB+wNjWdl1UWe5X11xCHQrQcwyEXstP+6Bj+MJ5SDNy
OjP5J0rLzMrTGEZmy8DRMHAss0f/bEznLCdJ+2goY8CsCz5mdtAWVyl54N2S7FJOE80qPHt6Q9A8
PFaGb2MHF7iU2YapZyJUUnt8GTeoHEesB0EhWMmJWYb6zLoqWe+6tdyou5NsuE3NdaQTsImU5B5L
QiT6g3cGS3G9+7xsDK2wjqBMnCesL55hIbSVNZJMoztlvIQTWlsON5kuSXH32FHrogxFoYHY2H+V
Hot/hK3+16O8LWQPow8n5p1r1m4KXxfASHTUXdTejrc/AsX40MLZJYUng0MVKGt4uqyZ2nXfqxNY
lnwbENHJN4W5EPAFQtXply4w9FbYVzcZuRe1FmCB6la+a9XNUMLc05V5w/kvyeoEGS0PDWlZZEk8
3zLd7ANJhwVVjrcoqcDMA4SoLsXtOrp5mvDr8NCsx9fyzkLLBzdVHmmKrKiLzqq/oq6gCgfWVfaU
OLnl9B4GUnqw/WTQA9N7ZBF14tZQ5/m+vUvUXPbZBrG21HkXEXM/55IK0OwrR7CN8jtCoWowgBrS
eeS8OtzSrydvLW9XijM3sPa0XD8u291DXNngjSKUAcEUSAUs55d7bX/AIaik2c6R1qZpHs4tGbWk
JbPUNY3/oAoP70LSnS3PF93k7abfexKpVvZG6u5HgN0hbgjDQ9bNn9I0cPHrpJtsd5Evrz7qbjKy
GXXVvmJiRqNCR/uhKupLSTdJA6TscSDocIJBTQUu5l509Zb2KArj8k51VJHPru0Rj6FuN5/kkFpo
MZNxEwyZg1EPjYel1G7GelvlRh3cJygV8EUNwC164ZTERyvXMVUmJi3WX/3DRbMyhkXCinC+Q6pe
38h5dj39YFkdxGqfMeyYU+xBWjo8aAaU5kZaCXcheU+FMb7867PD55MbvibjUEWVGS6CHvfofWE2
A+9zK7IoELIHh2fbT11ylZAVQzwGTRsL+MiL6UnFe47dmZTB6lRFZb3OAUzUjx9tJxgf5R5id89B
XrlKY5Z1eiSVA39jBR/ZPvWgXkBlmZ1DdOu8eJa53EqtjSLwRlEka6Nk44OAH/pfr2i5Tvy9HEwr
5yGnRbM4m9hl8JLIkP98orEnCB5N+yKkCxT8ZYFhksbyB2JkbjEsQ/OLgi/GM9fVDcvh+57mCZY2
kXf2TqPAA7kOglBeZe4Ycs9oDUtfEDFhgVelVsRrplL6OI78x2ik3VS6qMvonnBwjTopk/5tJ8Es
ndR4sdM1PUD81bl58JOs/OlBjggwshQAEW0jJInyRfzAtY+al0OtrExPOEH5mgp3hohaqOExIhDY
rOeQj3UaB9+WdPQuEh8+o1XYWAVOWITHguZuiAAlHnrmBRtWet8WOuihaP2nKsuZgbrMXjV+TYo+
ay+EYlUvDBUuZXV1NpOEsnd2h64HCJhN+OXQIjNlH4rDmPxDukxJms8bU0BoJp3F1m9p7UU/XbJP
OklAyggtQOpN9OXF9nWUcK3sf1edVwOWz9q142i3twfDHOWY4rUftr4gUyA7BZl6z+SgpJDJTHRE
HYFDbZpvMMexOnHkyEHT18iogVUvvrJ5zc/4Xq7yWwGdeBqnkJFiR4ByVuLaitYvDvHc3pH4R18Q
x2esd+ASVDcR1GkcJgwXG9x9gcrJI3bH65UpehiyCcznhgQ2R4UXVNeOXaQeTmqG0rLJFFji7Dgt
MCoY6khMJcbebdIG23yk7QHohulKb9czLnzDW7A9cLLIeD/d6J24dEGst5Qq98O7yU9SOvsALFEu
HxbCWIMTSh9hkwD+sHz3Zdj2oEdxXK0TLNgW/FmcOMNz5avryqCfrIpI+I134EaJOx42dzhXJFyb
oZEwhkSTsbQyjclR4tcwKpp3GYhHcwDF/m4SYNhnpPMfNlthAQTcs4XdISauDduRAbva94gZsKgq
jexzbIIZ13A6J6zO9dttEe+ZMgyb+BlpLsaLETUOn+EZXM2NEJdFnpEfJlX1QW/hlnpROUSibSB/
dp6RxsuDTka795sTKcccLBtm8ccHacWd8XGsj/NMCa7lXA5E0C9/KlnWOo3KFzGMehlDJaBMsgh4
mbenY5ykqkogUudcnIoLECJYMQ/NSPY/MAynb2RiKy9ZmFcU4zfQ4rAf26f+rxgYSHr9fya+5X2C
V6T3/aLR4Hx+jMwqlffPzp4IJSuNHA2iOytTLWT3guHs4Wp4XN15rR5uHgSs8/3Er5Hv7/HG+uK9
P13HXu451AVcOEH69VdhbQdSv9qUM+aYNVDKaFpzgkbW88gxWdLILoq5mFc+nEySlR1NEF7xTvqI
UQ5xC8ahqQpQ/7QtAJWUZ5OzYtyPIUFEVkAA2MvcSknG0gW4+KwWigOkdPBUsxD+G09m9wJhscv+
nPT2VjNmaLr75mK2IpnvOpnMf5ToX5qPkBBrRj2Q1FddbudGz+FkReS2tU9BiNtDXPyrqVD25Vh9
MMpqkFaDW3z7yhnLTXMS3q1tuUKTKZKwrU7tYhmOp2TiVHuPMjJ44QRWqyv02SWpPHjKiHB6xpZg
dNB5xjlhqvjsCQxxEbCVTmQyKbqR4e6ncCQqnuRZWgm0EY9n4z5e+1/1nmqQeSDIKc9VA+HcH7h5
tbprEKpshdVe+Jnto7e0FZ+iH/oZyeQp1mJLGcv81vPqamdRcVTmYwPJYgiz2ft1PANO+S+j6FLF
ADby/KqbIzJqcMHv5nS8MD3ARAszJozVgxx7Qwuny2qeUBB4Xw0VFr2BFKEnhRB+dPBuV9kDzbvr
WEpJ3vVPUNG8nPdystggi6YAwwouBIXdmWjU1RlzFuYmOoIBpefC3IhQwpEnpdJZuJrlCR+P0KNC
sL/Ji5F6VYIJl9j4gFvMV+hmRnPoLAgB+e393FXacfmmUjrGbLZHcKDf4gYBqUSOPnXQdCX1F+pJ
/izDcKaviolKc/nLssOMJmt25j3UQnVU0+VuTpDb2iBz8qLsUifiZYIEIPtaeMFRx8YbQ5WSTwY6
hVnqXIAZIvPzYnOSTfeqkavaiRKb+GCrW9NwU9DI451ttYEJKsSBxDWnZTGjBwXzqQXrz4tFmLdL
CGIjDeXYHE5Mubw1/PKEYQf0TKvOc9RCu7YoIa+oCOvHHIKne7YRxB8+Hi1xOjA74Cbs1z50DeJY
f9uTrZlbboKPmmxUi8lqpjfVV/6y8p7yJcB8cdreSLCoJqbroazwltTq/VwTBqYxgKWnHxu4z6BW
BZd5Pjba39/l42aCus5ixRn2yTGqBDplo6X3QrPn4yY0+X9WJVlU9krhDTCQa3+8GtolxMmU3u2i
2kiDC4tUhT5pdCdgNBZejfN9ffIlbgDhgeIdgeW+tbFzp9Y2UwB/iMt9u/J+knZOdMuYiUoZmpuB
KFxCGAX6qzIUiAQuRYxLAN5SjOXSE5zAA0aSkDqkyjSpn4RCXbbvvjkASF68FvIW8T0b8Mz0flu1
VU6iRjw8nFxRbzFTycYm5a7ofQZnhVLaA7YQpU5aVzmQ6YrVENtK0d/sCCmjGq4GFOrt/eQemLFm
Qqx5o1Zb/9ytu1YNL5T3DeV4rytCOIHzhdBqREm7Ru+W8sVK5v3Jbfeo23NOUOP+DIEAAjbQZJeB
zPfdTTr+arx/KjxOjahzuxY7huS5bxPzSYFPq65af4CIlTdcNgLXr4//AeokegMOtn1baZB026Vp
fhNPnqx9wbZL9TKF0H3FYUQGWCtVtIcVgISE+T4cE2z+QgBLPhc4teSBmr/0Zq3jQAKjEflGnoGT
YTl0kq66MulRrN7ezabPJYBSyJ5qZpLU2/dVzLN3vZUCpkwhXsvdRkd+4AfkhZmvA7gaKDV54z1/
jOrFjfa3Gfc+/3iehORhRbRJcvLUblhmkPmaMzU9fzaSxhM4LC2vd7pJLOKE4RG2OcrUbtJyAHtJ
NdpLpvksZYEd6ESzIeoD8y0d6i9v1ib8cfSRi9qBnqbDM3CS1IazNYdgcj/YxM/3U5eEGxXujUsU
9g1fbFEuGanXTMAUPXyTkM1O58g1hIzz0RXevth1tAz+OXsLyJRo1OMASy7Ou4nGntBG2+nWUVTM
fhVkobCLlVkPpZ1X0m2HGhHHlIkIy8l+plH6+SPuE30ot7PWqlnyrJwGTiQUUYyRNhwIXFYZd71t
x1tIGZCGaLLVqDiXEJKFI2V7DeHOAo6OK2JyWxm+ixRUJMJsBbVIskdXg6vp+fpV3E6AYk5+WvGy
jmHfv5bq/7H55PVVT579SpmwLgDxp3M5AVQTS30sn3j+RX7fOH1hZGY0z7PZ0WofoMGZb3yU9lvL
D2NaN5ravU+imaDkdknJOteeftBvNiLpObRqV8h65mj9RomXSp2GsPMkG0EMpu4q8ufDOQ3U8/5n
yKQMMhmSx/WT4iQp9yTNDbah48rrJtJv5QZ3gQaJX5K1uxV+MIhLFzg0JyeOaVBYurhJv44oQaXX
OTR50M/wyqxaQEfjWNcbpxW946yDmignoYepQQthqNAwUOp7ivtb5+GT19dKMFr+EhqYEvuRFEvJ
lZt0BqfZM9lk6hqjr4UeRu7QKrEoddoTbYf+ZPsqh9VPyNHktK/ShjGY449bcS4/gi/8EWQm3dXE
2HDIPE+6r+gAVFYPDH5OfbZopHH4vp+/fQeBoaH4BHq4h/CArwSmq8N2istDHqe2mSdz6Lmmm6Ci
RLOVGkB9vCQr08laYf+wxkD38ntCij/irAZaqKzHjhLMO7OSqhPzamh7azaNExrXDTg8DVMWgL2F
ezIImF8UCBb669BahBr1IEL4KCYrYvcxLE1S3cb/740leckzKfX3xVJdE5HMTVCuXNPaC1XI8GbP
U2DVYkeXYlDVPshqImVXce1TGXDFzDYCmN9kzPmMJX2cq8nw9He26Z7MxNBC6Ui3o0FlbYtb18ZA
vk3PocTUxZEpvx29is6bbJaK3O3J4yegTiP+zkApWFu0MSrbdZW+C2Jap8sKciIKOswYqibY1t69
G3ikyQ6bzD4LQTfxNWMUULAzgPW2l1blHJ4XAqjf+RDii6MnQZnRpdLygAVFZvjSAtgX9hZCE6hZ
TqsPQ0diDy4T7Vu6q+aTjfbuRNKBrFpvllRQ/5t0TMZbIfJQDp9h7E2IeCs0RP7CbnJi1WtjZi0Y
fBWRvYb0iQ+C98Bdx+Lw7qWCN1kIc2Beyes3kTps+rhFdU4ScUkbsN5DTH8oB4e2AypH8FPwLmKj
mn8qv2FuzV7ka+hS96UX1DvXg1ufgZOT8VBV3qkt4IMOfF1yxh6avkMZaVLd0Ygqjn0z+qIL6K35
nAmw+lXm2rVMG2oZi+AGm91abN4L8hIdtardukExgL6EfxdAqWY4iVIDRhTdQwURlNTAz68u85VO
K42tqdZ71pu3PmBc10VWzQL0FS1ou/VN5kCXQ7YS5JhTiIOuxCOYGj8RHJSh4cJDRaMAphz9qj9T
Jz7TdmR1XyQaP5g+w2RK48690x5GemEDm13RSrHYSMxLDjwrSlHBg+Ca0sXO9l/HEguTc9v03vdk
hi1bff4eHXp/zwx5VdF8GAHTzcbRsosdhd0MOGR8AhWjrDtTkZaZJguxzWfzCmm8fPW8t9NBtB+A
g94a8X8Fnt4wMndhsAJMU7Sf6W3PDrtjZKwgG2uDVPZ/yyAUWCjAGtXHaJeqY190/PODBULZ6aTN
bv70lYJc1i3ky4Ww4UVx3+iwO+7UZSvMPbjkp+xdPTaZBFtvmcaxZ2WnnqJYGCkayt9HGmNhxruV
2D2eviGKl/vdQgeQWywFXsKJOZKr8fuFSA65+4dG3X13Bym2ZUZq2/l9WB8yFjyhReR/GRBtEi3Y
zo9TjD1Q9XMoD0RyHKuttoCk3ziiWLMwurxV2QljMxvGVele4YS9KpaaqaZaaWJhJnr5fYaQJknX
NmdHQNoy3LOO7COdTE64cohIaK7iXLfW3hp0K0MGz/bOZAVU+tB0SprsB0TNOR99dpIpkt15VOwZ
zQ+2SLUGv0t1qboxlp2r3bmhw0xXODp39BSuZsY7RNAkd9W7gDRVFtITGhADl/Zs9HkLxrAa+lqd
FdHLbTQKIJXQ+2zpsWTVfvy0Qj11tzNrr0ibsRkd4b/+W9i3v1pmiD6U5/we47D6c70pfHuWUajw
/0iPpVfKg8/AbW2YzLus4ceiSyE+jvxjFDIAFOchh5BF+s5i7fEUuqwj2ofNSoxmQhiEc1WeKsIR
6WjC1lQektMFSyZp0yRqlrMzbjEtz+JYb2Z3Eq7M2FN+D/hiScobm9SeU9TxTgeOwgvJ+Y1Lh/Us
cdQREYoBgkC1rsh/eVGdDNUZ0xHWLOts+7jxvHCGxgx0cD6AswsERjukBFCApk9og52BV187ehtG
0h/322NkpKfrNJO1n+p3t5g6TW6wY7H4xD62L33xt7wWE2Rmf/OWgExWU5UgPYrglYdDXlC2BsMq
jyjPADimddJxgZe9iJqeatcph9OHBeLSoh5Fu0Hh5lTQ3qlHQ6gkGHx7uoKis3uF4xheL13aGH8D
+2tTJk/O98T2THU9amQ4ctJf/K7+0hZkjzJDd7EPa/Yjma5fWN07yGgAHlZ/OEy7VjvHU0YG4aY1
N5jg7KfyREZmZPBKC6yOe/4FEo2c7KskAid775D+CO6GgJjIjO/aC4+jqEe71Y0rtNWKsBYEeoAu
z0FbOaXfHktuEPTzPzop3SO3lfYa6/zkC9rkK9gHcDOtkGDy9e3kuL4ttC2u4w8r9xmhs+Z+JvVk
b6vb83/Xat9jDLzwwHd36y66vtWpHLjvjutEYNq2XB8ZAiosulBocYQLjhKwQ2xLoWGx6JymFvf8
j/llg3OfM6uaQH//VqvlR44iirDBqbOUrNen0cwI3a082wsIDvDSPp9cqyM7jPAfPN+Z5GMio68c
H54tf+V0mzJDzcuqXNFearkxWQWPDwNDFdME2BXc12PB8U579LsbnCdjHPDAw1DQHSYcmRp3orhb
3YFNFxqTTGUby2eBeqFZc+pB6dy/IjyqFbexe50uYD9BY214TdYYpIRX7Z7ovj+RRQj8UZS/tGO2
XoaTWkTrhPKbrUsdb6QGkNGnu06IskIaVsHz68lVMBg+Fnjhg9ItmZzH8mknYNRF/y2o6Cl9m4+C
m+b5PUDH1ZbyiIPZAKLgng3ZevvS14yOR95REf7EmKY2Nan4CfBqMmRqLUTpZuWh5lxMFsWB+rO7
A1YPjMTEJJmBuq0F2eD6HGnABFTuYsfjivMWIXpMf05hJrDsP+4JTOQ6APAPG5M+0Dx0hGfXQGE8
V+N20fIBtVX2CG4qQpvAWrQ6pV31YlI9ItJ+505zbz7SYW5RaqCWwO4hQvcEQvxEG8Toy5kHorV9
xOkzEkLLRlLYln3y2+wnia7MUAlOVTK97/ezZSPGgptTzYuWieJXGMrc9TeV+ZEBv3C7KaGUB4NC
tBM3fsFyx8VQPmN59crgHcSHoSZH6tfn3TrEezlSiKDYRr1NxQdnmUxN2au5qgWqhGP4aP34KuQG
9RYnCvI8KzdIIapjSKbcsOzQvRPYyhbEjh4Lp80zzON0f21Ltzz3bbFFhWiqCqVk90StgEbkaXOp
mnuFILHvwiCxb/S1iSaPDPFGC4ymDgdQeBu1HLl3d0kM1vFyUO4lPV+2EwCmPjgmthIQ7PgQ2JNt
9cxv+6w3YTxrgQTG0QxCrmpjg8LRKNPvDJxjY+gAThSvK4EYj9mk+jL7DMrxTobOLBOH3nCi8pp9
9h+SzI33KgvKxJ+e+kop48WPDdVkIIJ/gzJ/cg/oQd2hzIBJn+cMMFtzsxt8qVlnMGVHmJuGaPy7
HIEXzpeaRoB4esMB/3QXXeVgWhNTzNw92H0R3d5w0oNXScWFaWAMbLygcg/OnOyLt9kG+boLMzso
htH/mD3v2+ko1WsBZghmafMA6vLeSTgrJfu10DmGOl4HoUJBMPQoD1wfwwuoyqZjmHN7mR0KkKKE
u/mcuYkwaj9LhZwnIKOXRYLK9oZ8MWtLmV9PWPU46y6NJ6xUXOqt3Qz2xndUq2YhkpoNzKlSdU+n
Y25KGGC5MPPuPgTQV0pZxa0OnONKPQB7j6qyf52b40tuDLBF0+q3K65rMNKY/RTJEUH4LiYLnsFz
0FQYVCdjW770zM3R716J5w8m8Voa6m1T82lDrVcvgcTvgbqgMSHe0kVXK3VIYuJsjt1whu5O2Gw2
lmyAsEz24NR3tkquKOygyo6P0NRE8uvaWPl8N5ZTX4LUpkvHeFn2G+0mLu+lcnIV9HU25FtcHNU2
txNwbQtXkm0sfqup+te1pO1CEbQmbwKCTukN0wUgHAWT9T1lU0nlabH0lvD7SY6BEHdOixQLjgUD
YZDpCgylf6w2iJrevTD04m8uWSSQ/4z7mbpwxtmi5XamdglvjJYAgfflzpoaDHixxaJcSDAnJXem
hEqmLFYiNQu+Ugjjh7Vs5x6gJY09ox2z1oUb+Q/VQWLNGaQSyFiFw8XA6YP4cqX2UYUqEzxofSjB
W5IjyK0CYLEjsxDBgndU3nglhY92bGJLQFhxDRiL5X5HD3qfLEso+jCEUcCqZx6ilSxN1lHvLTw8
ES3rBZp+q4x38dh2Kpmn2WOY3XE57lleXBu6kE/wD6R1K4utzfxlZxCk/PP5QO9gefu2N/AExaDR
6DIu9f6DSaaFQm8PZZYMet/6v1OjjxGgAKhFSS9xFYpyXhSU/OmLQQxQ3nAFqnTLDFWXPCWs2mpX
9heljU/1tSZfZtn/uE2iUdou7okutX6xmWrfxZEBWQczKCbWo49RKC1l7Qzh/b3EENsiwHiIaDsf
xoGrTXv7ugLp+35ItdTbb+yGVX8N97DB7PJ/EUQYIKCuHwLLGVa8PUt1bSut/fn6hb0cZOsKzB3b
qyHq1c85OjANnuZ0cx6JHpkQ+vTCC+NIWqvZsTAT2pIgfD50xs3eQ76RBL+4KHNM8te9JSetCk1D
0crVCzCqQeuMmcm8v1CwzZosI/EhB9ypqollHtuxqMF7C7Y5au1Wo2uk5AK3ZP7M9mSx6GImcGji
fUasCFJVU296rm3S4pO86XXGWqBmpu/mu+KclHYuYmLunsK3E7uBZE1QytcZ/hIbeowIOZrXOaRb
FBLetBTfX2WS1Vr8wyZ9SxhxjhiOt+2ACeDr5QnEF3OkPPpdgE2y5FeIFGNFrCeDIshCogOpcIU6
gIQuqC7609f7Cq53/qxmNOcH4DypyqfBV/B1byvkTinvF+uM5UEDbdmX+argTfVsuByiKKajnaXy
MS2zFBkDFbGl0RrdZnOU3ZVN/5dRbiKQ1STRT6MR1hUOWl5Z1tV+Tkdbr630CUiYmGpJsW/2CyW9
9/tWwdmUF29wtS43gmSUqFtTN7o46mkaJQQHNCLg6dD3Z01GyltpKy5zZQf/p1pRbZlb5sR/zmFp
ZBo9PX3qbL/ZDbHVSkpseg3lKvRWjmN8a/+AmxB13FWX/kJYv7cUIQk9W/Vea/ChE5S5VtHcYMHt
F3BqZkx2i3Ob5IsQnXXlOCOFN9sP7l0gizkc3ypBsfkOH9gmuTAVaOOZJXqQY1obayFmGuW4RXru
bCDOpicVop0q+Eax52moyDjux6jT7AYKIAGIa54eWaEYF9+TOWd/vY3EnJnW43jDXcbOYhFsvZML
kIMBETbVUzINV287Sm0eUUhE8hNZZ020PRHvKnyS2uFmjlQojtuh6rYZM0qQmzV5p6O+djhTYzLK
Fp+FMcPpCza/2/JK82yixAkHHIS5B6JQq3Gio+apjjiB0i0WtKi4FwnsRELpZPY9ejhlL42wvWQy
5bzw8rX1lSte2UU1Lbde+dl5cU/AO9DqokI0cLKWeQhVSQYD123akvjBKbKgdPAS8tnR+G2m4nhz
f/T0PQ4pI59G/gM4On+L/x3WcmuagmnNd3zOpe946sFrNTuJ0+iXsSW6UIt+ryc0o5/SrUnGqNF9
DMeirzTh+vVv0Xison2aAvPxXtp5Cd02mr8FkDLDhZmm+585+cjhRDE2EUA+EGLnLUTTod87x9J5
98ZpOrrOZSsTeH9iH53gZ5FyxdQ55CHjhvqZnN4ZXVy/ilxLkEPYZi/jETzNEdVEIHKKfBMPhZdW
w7g8kO5Q6lf8E9/uLnXXhcGlptBu1wAi+Yloig9gEd4rR0e4NPgWzWpvaB6u456rWWSDvsK/F/c/
DIwrR9PUKpxFcR82GjsyEB4dYNfagwUbh9cBLlAA0eTbcTD8xDEdlgRN/UhIsU0R/LW2B7FatTOI
pU211YxB9DLkDM1nRsE13JTZliHGHOd/UskCa19djO09Q6+LLeYefi9jM+ukzQg1PuYBcBS4zkvK
jb0nZHrLfg8DxPGbU1ZE9Tvmh6nTvBNfx9Ytr/DJv7/ut/NRv+O8fj/GJLWhMEJp8ys7RWS+TeQz
FvIBd/yNU7XVvpLn8G5dQ+E6Y1uV0mJa8LN8tNLrPHBG8WfWwl1LgiAbuvMcReewr+FGGiR9QReD
wTPPCL1sOWdPX8XwWWERmTj4KkvfWz/+VckpmSU19NRmQ9rALGmx6GE5NUwggbm1hkF47VdE2fpB
eojmGNXjdiqlyV6RT/dWDEcAWtKO8JkioaV8jr32voHko783nnMXDTCu30olSr3T95/Yhd3lndru
AjFtBFh7VaTQXMYMRVAOrmVb0yWVPIWuvqYz12X4dRl4M8WYnYg7h+y7plL7+mNPh791Puq3HnuW
aIduZCfljMjUjFo++niKcWOxD9DSVnRczEhQ35wXt44EmEWF4O4jT1vGqccIzP/HTKLjAmv6I/ZG
LTtXG0PFVLNUkKJ+Y2TaJjVY39n87nfZDN7LG583Ynyrlp5BRdTwe7RTAjE0hzSo2thm6qgBPBl4
uDerxq+IxD96k/OYnpVw7Xu75HbmLLoGFGN95hq0CutYjwbTd3ovUpbViq4yEPcBetjjRl/H9rKZ
ibzRyJLq8jP3P1leck07bC/myCVFiNC/9He66X4Et3ERurNXWdYzUX0qjeFBVTp5N38rIjA99Vg8
hOdSnsKLQg3w3ZCpkHcac+XdUZtEM4vOKHCMAZJyxuOhx66uV/Txy734+O39A43UUfX8xjgJJpfC
Jn7dphnzLFB1521weqBWVIxFRKyVhiUwgo858Pe57SBGZLIEeSzszZwA/YasTa05+sSrUqXJjcXl
1lZjekVJaqXyCUVRdAo4VrQQ1QfgeG7+hHTs+t4s5LWnFNqC7eLC/jOBWTNzhROuaS3pJM34+7l4
2GthSJk61qr7lZQRzN/+4hm93j60ymX+ovJTNr83zljfs13/QrPseocNObIOqzAuadzSQjMDcb1w
U1mSkN5EzP67rouXUDeil8eyOpt/RJnc9kAMBg9NmhBXjtZyYaMSA4/FzShM57N60oX1HbhwxynT
sbba/CjP+fqufaOzzUvr6Ff5CGG/ijaTQs7FowhaoHd6cX7vUeD6YCTqDnGY6nPfPjoKusb3swXR
3hL82k3Jiws0BV/EL0nX9hE828xeTSuJa3J70h5sbZR9hBA9kWQ5jahN/1RM1WQokTm2iT329fX6
NgQ/FMHBcHGNiz3STnyTX4pfVYb4lyyXhricec1C4ecupekBdP/xJT4MIyoDvz67LGXZ3piFLd+9
wgXYahmSEYnOHT2tkEg+2Jry26deRg86C9hYex/WtWzQrAyf0/EBI5hE9LCYGLzUBgFCAB9PkBXJ
/hIRCRA6Tverxty14sww/LfIqMIA++kwHP+9FgF6uYrYrYv8NNKRcQ/UdW9HpKmbuMBl4UtDStUY
IUpgXL9/IaIfoplxXQdEzihJ2kksYW45LC6DulddjMsafXfHY0Mq3i/a/Fjvv6vl7z/R2T+8BAF7
hLab4jYJRncIkwtlLcENcg44c2zOc0+SKl6Rik7loipNntJNtrc9DtUaATbPmScmdpAbdmROKnox
VrrQa7dSbJoCQwPv0z4geIc4hPurf9XVMPks7MC3TW6hX3vq+3r2Jz+lPCQxZD5KXX90tInRUvrg
i3KBl6i//ldfQXAmYTJsNOec0ub1Kcr9iHYlonn4nX1qaWDgl7niDFJhOTkF4TR+I8Owky8f/osl
f01hHyeDwGoltnoxz7o+Xw+fos8ZbXOMPmSmppTbVAzzbdXuOIJZMNY9Xt+M5dry5NTFqjq2OqOU
tKdfBQvlQVIo9Yqf3YOhJJmedyfJ3Az+q++209e0PV9iWA3nDnTjKGp3Aj/sIt5JszcypJY61VhM
aGkr7xddCgLwr3kluuELSIB3Pcdtgx3o0y8EslTsGVyKbwcDowCTxF7fRRs4xY4/JfyzWSHbZ3CP
P70n0zQUraFi2tkeSk8LKx8QFmzYppzhMHmwSIQODq3cCDlDDeuLEHGGnfZ279/21WEX0sIkcwUA
a2myG04IlbrHxgz5T1N9iL86n2ns0a82O44gNA/QniQf07yRZThcN9t9a8rwVAJKaAgTJFfR1HbK
5zxfA+XJNlTaa9B63hDek1mnX9QPdXRLvvelD3wq7oPzLlYtuDJlEWAi0eUcTJK5kTGOKPI329WD
wz5CKYXsNLCxy2e4FVL1BbvIto9k/g9NE5oNx1ASeOYOrGY98W3Oby1eGRi3M0xLdXqFHbDhdhfG
CecPHOWkvQs91EqU2IPWGHqXr5E1Djbn0m5Po044GGuGl+uFWqlr2c8dwS97neLXrH2/VWc440v4
JXpsRlDn/JD15KsrnXqjzV7sotmNTBampbrklneMIw4oANWkcriDg9ZD50aXW+PSa0qTjMzRg56s
OWn1zvP+K/r5zSpAEpHE2dmJ8shRA9/BbFXIFcjCw0Hs7iSnb5n0RgXNIifv/wd0InVS8Vzkfnq5
PJb8vfuBy0EWLsjnmQkkbd3DdhvzRFnOusGw+wXR/bj5qJo5yDnwA2FRTV4EU7kyGudELZ0KurNp
puxavOo2N6HRh2eEublzLEfXZsH3zNrgU4ThVD1ig/NRHCeANDeNYj1KXVVC/Nw3ydkPGd4bwfIJ
UQsHCFNJmCh41mNz9iRL5ec9dOOi0otIRlKJ35t1wOf6tdeyROpT1nZJXBkNYlp0XRuLqnyFNp1E
1+G0XJ1hHBHYlF/Ax2wzZTirysTLGwQjiAAbD77dR6/gtz85OV+WSFVPBNhfsTDCYkRxYEuEAY0c
etG/cktpc0DuABM1WlEZBidBv1yhbdN1PmyqN0xRwEyZujZTaHOxqcT2OIwSmnv7Hbz+Dx7U5qH5
xeG7fCmS3/U/etjv+vg0odM8KfTBN4JANJEkmzXaF2exWn37zDFsF0+1axj0dZqBGCltEwzZ0/Kw
RW5WZGxerA9g1tGVa+7H3b5z0ozPDk1ufoWiu4qcNxpnuXd4VJ+fW18Reg0JjBao8Xbun7ivJBQG
Q9iCM3N8mrics6T482xJ8qvRhOv7qM+Bnvb2g7mZ557X7UJei2PZj52O8aVlykFAMyuB0/oSUPwB
j6VrtQKe6VZ6U3j7BoDST7GVA2kzeWmnNa5D1/frozvl9aWrbJ3mUuZUJOKwV9UFZrbptZ+Tv0kP
+nYqtJCrp8P41cmTDCw5E5/ZHAxfB06Nv5MrkhJ/G2EolTuJeza8Rk6AhOeARNJJz+5BDc1R4rUf
xyirbl+xaIYNbBS5LxjHnVL+3p2YrTy5WAh/bWPWaBOSDDWIMzz8v+GpL9FeR7mOKcIM0WcY6vbA
rjt29XuInQEA/CD3ub5JcZ64xE3MolgwZFkzlNuMRm5ohehC3iWCHkOcnLp/sIebYL/hYa7k2ddc
sLstY2hShjmF3bzxcL3a/NnEiHWe/ED0URt4g6MTqEeQYOjWXfwilY4EoLxMCAvrWgnG4GfDSR/S
1wO1pLngHol+PYcf1OPpN2/HHatiAHth4DriihYfk0h6lBZvufNZc3dXI8CgydF/6z5d1FUOYuoc
PGGXruiFf5yCeG1CV/imkRSMtXYw5ZshoHwzkYcmEWunR6JZX4P4pv7hLrmhVHKxBJt16nP8dHC/
C80Oy3dN1AuD6/ZdFl5qpTsFFfQMSN+7VYJ09jXpJ7Pyaw7oHFp0OY+/okMc5S29ac9N7phSI9Zp
WRIa6HSMWE59GkpkXsWfR86YU3RuC62dQiRYGoFUXFhsiIiu6hUVtKcYgeGedUPypW2cCD5pUV7A
WJtfWuodVQoOGk9WNn//OaENXZh5PQyH8i9GlZHEDYFFLOn7g2Ht9oJanhf1acb2UPo1teS9/wXf
KWiigfnHuhFMpqgjR3tB4EdObBppp0KQ4VBhV/lJ5CAk5NX2ft6eCuVVJLBJ/GuWTCDrPcnHGuR0
beMJkav8rKsnQ+KHO6PtPv53I8DDnXCsWfFi1ng3ZbxbKOPEeiZYx+ow6VA7nXDAfj55KpYDRt72
QGCBEBknG3se8pxnZuZk8SisuMaealz5wa6OW73U2VuTikC6FS54lzzKQiJRRc628zu1nKi9bmv1
Ah+9HhTNJ3G0+1gR2Gsu4+G8lmsGPnuWtHuHN7TWlcz3chphIwZBOhEuIDbSlX8zJ7dZHEFlDQeE
jpMwFdJw29HT5R4WvzI24ycwfyg5HOVELTrjddFl2tRddEZ4qHBN0ICRXf7kSLA18pSa+lBYh4g1
+c+qpaCrU3A4NX0T6CvCU2dCF3C+69/uFHgEXSVRvCP0ufMsV+hjid40NTprtVOcIniQ8GYhF9ys
w4/H6LjrbPTRm25BZCQr7LHwll6CFoQsPeCtntKT9qqLqh/b6Yi7h6W9pgCbnh7O09rITRnvA3yA
9//KHlAOskiDHWTHWzNluVGkTYI0R52pEwVmfP0iQVCWUwDtD5F+UzJL6aoU6VOllwFzdphRVdge
rTITHjLhFbchA31PrN9fxFfvwhG0t2ew6YvpdbtgqaLBwrWbyIWKS+Pk4mUgjepMrac7K2esj4Rh
Lvh6AoQGxa+Ox7Gyu1edhxq19qm/AxkV1dDi5xgA1fkwS4lULh5I2jdWcI7avN0KlnrZVu2ghUbw
QLHq+3BvSwB1ebK2UggH0VobAzppF6hQL4DCYL0KbVVjPZxGkuvtB1cLAlnmLh1FHbEEVymszMk1
MGCWLKwcAfgg+Q9TixDjOXGjoTEa40MHYoJwwY6o4xgkXQhZ46rSRFJ5QOaFQQs6b+YHwSo/iqzT
iulk1pteYGU10W1ejLYpXxhCFav5yWckxf3S1OzURiubz/5xc66D207M09siJcpcaiTR3HUyso4O
ws3gyjvibYLHyk/vQ8uQMKs2G8eERCmqjII6rts14IuGAf6SINleiCORAq5LAjU4qPolOmVBjkDS
nfqTRv2ythf3PEvLydkEECs2V2yLWDzbBy+p5E0OuxGS7T/sf9rn5Te/P5UNhERvXpO4Z/DixoZH
Wzp7HtcnsR29s2/ysvWIf+553b2aLZuhunG9aIUmTnkOVD4pe4ZAO2IsOh8RvNqpGL3Hn2TIU7Nu
eXSrIbDAyLstsfzE5Q5c1GzenV2kAkUyeMIAZoVxXteffg7dCrw16ifF1nyB0jWptxU0qj/ZaQTW
HIeFRaDmZyjXXbGdZZlrK+SUDuYBBejH5A2aC/Gd8myCvW0uyeAcJHkkwvBbvBLcUQRqnVYi0RX3
Kb8Ylvi1ceac8E/HmeGmZ7QXc5b8BzIifJH0dXoJXxGCEFZPPsM7bGShKKQOtabE4Eu9YI63p8Yu
O6vGlTSizFUW4gsr66tETkh0+/PvTDrTnsU1MK5IC/PNRknjr5ND4cJEfoyyKzOuk6Q/uJb9msNj
R8QpP41/hhOvQ5Q57qdWCIvAh5NnpX5ZGQvm8zaBQVNFr1InDZSdjXaYwA/CLvk01ofY05DCDIUW
c32ov+O+9qKGrF+iVEV4RiIonK1rFerAN4hJgcOCYOwE8m9v0m84LtJYwjx1ZHgo+m2K+awCZsUU
7H5axW8q+z18vlDSgicxsnasf99BftENj2d3cafrjirfFffLCNie+HOb9gHSCu+MbLHXJc/QZ57g
P9++aviTb00RSUbgdQZXgFmZwea2wbbICkVBZEsHtRVrRDEEIXz3rP1PfXDIef4XZAHIk1HAo83S
G7osUcWcvctKZO7aNz7/XshxZzb/r76a6/jbs4MftaGh3m3kjTFR0woEJsKiO0vat23kdsJsJqiK
CtpMxkqKucEtWsxUb5YbUyecdRAT5dhPg3N1bnhiTy27GBO/6SD6VD4KYUi17i7Or6wiyCgeGMF9
ulQ6eBJek16IyF8e6K4YV7SsfC09wXNZ8lEMSR6xoLJw1Qaif2g67BWu2jMbVVWzDU9qXF5+Zg7u
tc+jFWMX++XqrwwEC41cTkYOvS8qv1tig5q+o3RnkZQ8hZ0wxgyhWFY1jPogMalHOhOdY9+CchlI
GcRwsK9dg6hU7I6BibK3npIdiXjASZCP+i6qy8O/7tMWIHGoxIi8BU/w9AaeIcgPPnOfoR1+0Vf7
TE2aHUd8JLXR/PIHEzutumfcB2MxfzplnTiEAc+kbvlbURQ6P5G5nwD15SgGBnNNw4OKzgE+CsrU
MJmBGR4HDKZJjbANerNuznHqCdx4Z4z1yfihhqqC2b8UpzACb1WTlMZ6YlTcx4+Ll01GREvP/sGS
dD/9keEnV5VzWuwrU8vbQ1vgwy+h8tYxx8zXtjrJlVlcDONfkoMdKmduhZGVYxf9pRWzohH2KMXw
s9j0vf09B3k3pYrzovvcJ6qEGWMzwQpmHGuyMfuGWEaMN9HN+Qzow60RuPqzg8v7iLbhiOBbzk8v
Hw9nw9tSZ93ooucoGFzfDAMpcmUoRnexRFho2lnNro1OxgBs5tQofMyouYhuvRDZ1IQhoZ8YZwKr
b6F+GtFumwT3Jw6MQZo8QTszNV//WQgn+VPWsVrFDDQBzAv5MTdwHxse7itHySX9f9p9mZ62Z5tH
gix1A6g4b2aQ4GHa7FFgCFRJJKu0gX9/35pMXtU62bPPMjYvnqFyZTi23eaut3i9Um6LTUjRocrf
UtnHv3QDF/bcHiQ9MG0vEGRYMQ+csDgHJeFgKS//htHWa4AJAk/nF2j+lZ683je/+LDJJIvHobXc
BY+3W9GBsfAcyS6Ep/0IjwqLw2vGTNaW3czqFNRm9pz87O6i7IdI/BI2w41e2dNnrLxpqZuh/Yqb
/1Z811y/joT6IzSDajpFVs8Eg2tgg047A6oBWEiA6Afo4M/uHyKrPgijlgn/OkaLNAif4TMlTn18
A4HiFGYn0l3l1GtlF1B82KrhzqehlfKjxkX6xdSOD8gXVsWxkZrewLgz9C54Eh7sktQpelWWSC/Z
Gpx3A85wnxfMil/+AcIFDu6++iwxLhOqu96gLGkO9VG9DmUrH2wx+PXa1oy5x8Gn10F6Q5nZFz5F
FsjShIwkskb7WHAqLHUCNVv0s0FedWodjmKilPuISBEX60A/i2gzgcIt57G4ChmKywmdziwRQgYa
5hnAkDa7E4fxOY0OGFpPlBqGyLJny6S2xKnoKW93JqlnEwdz41OaD1obW7ir06WO1wvet5/W3AjW
tZPGTng3KBj13QL9PZMARm17EXIUYz+TYP7t6dBFOuLdYEFBQxMAkwx6gq3J3gdjWjCX9bLJKemi
osStk3etSFES8+CVNPrU2PdLGTLwDY87B8jicAPqcW1Ums2MRCNCtu9ysVSVMplKFQikwg4WAh7m
d/sE6ju4srTrOy2h7/PCFUH+SA005yY5e7KWI7dfnY3ViLTSzCPKSvvL8n5Iac7DwDh1vOpK1w0k
lc9x0EAUul3fQqFFy7j+WJWDDfu68TEodjSHfih45DkMkgwJY/FSwhU7WKcwoTY0Azgmqed5UyDi
ZWSqlnDXyCuWfIFpNoF6YNlWSGh3P7/WF8n7hjuRRZLtzTNh7m2U2WO/39BLZZDXVNYO5laA1QdT
x1I1LkRDMa+Hum/aOO3bxGrsaFB+3u6PJEMlgm+Q7nT1tlJK3gnSggFfBsOAnODdO1j+KEb8q9Qq
UCTSyLz+oZyr/GrhNwrALU7zM2A4rkG0o/muoHL2RoW0fjbHvzKs8hfDXebXem8XOzWbbFR/+kCd
Q63msY5r/IF9n7pXY9WYldrAbse+zqrxGKtthg0CgKxmSWGz1QVm2cxog5hR4RxTBvcGk5STFy/L
wpO6lsJWOjGxdgq1tlSu9K36YFHQ3RhnCLA2q4ghECD4zn2OOlkCdDKdF0ANaTP6OBnPAj10Lwoi
1e9Z5HSPkTUbxhTLgOpbqCkT2BR9SGbfsrnFxvk+hcwU9x26cV0VJBRvdhtv570HosubQXAiSWBr
CYuArPE51IZNLvo6VLCM26nAwYgWfZ5gkXLiFT93BIY4gQsPsd19NM7PvrkU+lk7BEt+1T4nv78D
omeig1HOb2T5eE3VvuLuY/FXkJGte6cF1gTntY+NgGm0roOyUK/+h7IqTa7X44/0sYB6tMXjETZ6
i4iqaN4UBOh7JatlKbOxIlJHqbIWGd1qE8EABTg1WB+x6jODtZ4C4rMiI/Twt7OCkoUN5fVPiwgv
ER2HsNM4x2oe2G8IsuKStD21EWZeEh0z7ayNySwxeG9/dF1BRPLpeijaCBzm6pTeQ/M/SfALigls
SSSd3QruYUc8ji0CkBLN2BxH2MsR4aT1RB4PUW7xVM5Dsm4rfBXtNhsge56+IzUOpFs51TM44nMO
LCia0X2MwaFhzy4YHf++2297Kda4ySSCZiKPHT0ckG67puKDdPb0vVvKuCjLJhh+7L3s2hDDpzjr
hJSVdhDNszvEBO9h1YPdAKNrvvH7hvjW7LQg3kWqzSr8WflkqS2e7MxFbI4p39hgg72fokIVrZEH
OfYGoZoyeuUX8gyaWwXMBqnHAJcbJ7CnADcRhC3RIg9QXmzrHjWcFEZ8vEt+ulb5/GtQHxcz2N2n
nvI9ixzNn5Mio08fa00e8PuUawkPWOXjHfF0/w84FPWlGsA42zzvCjN9dDfYglvUIPnuwAvIR+bY
O2vP1hwaOSohI2oNCRkbq5GZgxMSkvVJyJ58L8fQEPkDBs9rAguBGhGp7yLxP7KmI1qsFgn9L025
y4WdE2WKJQM+gFIN7tsXJ2gK5irQ681FxYgbSfz1WIiJRMlIKoESadfyT1eDdNjFhCLDUV7fvtQx
SevurwwY6DElZWZv/QkDnuz8PfNmamaDbSWll06bYgi+sI8UzL2ZuiSxYBQY9wr4mqlgp7CD+iv1
aRlL4qKs8bu9so25lFSH2jQiw9ahghI1QKsOcMlMtosXafWBYwriIf8LA2Kwvw2z4njI5RgbFJ1B
geNBZZSfcYHVYTYI2YlF8vVGnVAc/UGwQmIrBarW84HzeHAd2ioLLSd4HNJ7JNg5iMcE82u1fsle
nCfuz45pbVJlszKCLo65IEDY4VxrvLtgfpNggwf6ilCHZbIUAVkc/ui82U+d1N87mOQhdeupx2/H
XHku+Pzbh+EIwO4wKFga2I0FhNVprSJXXs55m1+qv3MkiWnAeuOOIJpncRAXnoTRpGQDIegMUKjC
DJUiJE9libkDS/62IDKXic/JpVB4CuGnSaKZ5lQaleQMXDCDSdyK1MRFymdeza+OSyrZLvgES0z7
ms8CLb6Y7VOlKdsUMb7pjQwJUB1eDlbWxRfvn/MRRTcSl78AxLDS35r1qDGGw+LYQu/bAKze3yUT
zbMbuT+YyXyGCcBlAv9i0+LxKUfXaqGYZ35cu0qpaK4uiIy/G9fiSCElEC7GEeu27luNY8rMnrkB
W+0QbYa2YqUvo4dqPUL4D20oZI9V7D1kJL22As7j77M0Iq9W6xMCxh3HlNlHeyCZdC1U3iSfa0Xk
kQKpC0jqQVv6Bu3OyEGzvingql9inAyqrwK8mNJYFvHvUK57rV5PgkBtdRJ6E8L5LHnkOQZ7kuab
jSs+6nERbNwhEgIF/EIhonsF4+xWjSmWttJMeoF+UHD4tQ1QiUDIgzpaB32uYq7/w2fd6l6gWfZ4
FzETtQmFbGRrEzeUqy+DGhNUFaGVPOFDQbF2pNeID4zdDTfr8Fua2WTEkV3ssFs85IC7JbfEI3gk
x+evYkvyDR1EgU1d7VYk0jg6U29+3TmCW8OlHhSb2ENpURq9bTEsCGRtscTjUpIawfbuODtQExTw
051VdwgMb50zdWflG0TE8mmmjqJLg7t0HDwTLdDoQpp3FruEivTdvbkfj5fchdkpMwbhqXxYDbxl
5D5yb/rpNdFdvnHmPGcoYbQksdbl/Ufi2juRmnyV+ERYh7GV1XG2stpQX4WRCRg84D0RRNtfxfvA
SZOtJNSy3aJI8WVmRu84ovkuyq0A9Kv5T41rcnAgrO3feLeKiZ87Ikt+OIcrUe1xxNptop8xy6PG
GGnxTlO5SZzwGDs89SsY8QEui29MpvsyXEwBQMGQ5CATPNhAOZXArNQy/i9pRS0V+5e3iHmqQ2Rv
gVS4wnpakzHIQhXwIHbHWetv4IChtpHCj4ynQd1PZ/bZMI6xXjRSvOZp3eLGqxIwU97Tpot0+As8
sA+Y+BqDnWUu+tpN4fmNIC2qFoaG7MOHpQLJCor70HyNUKzgUB3waiEK4IY2BYpec64ks3B/osj7
fz2123G+mAWmBZ7KjAIb3TR/kx9rNe+rX+XxE2mbrMWAR+m18NHe3RGmQLFarL9iaDYSQrwekC5U
2lXieOyTW4febBux+pMAkqy0QZOnB+yIaDgneMRb7XXwSNEUtox80ix5d4gbm6iUUGsGs59Fx8Z3
ArwfJVPJUC1VCOteUEwvW8X04Ci1okDOn5znK8wbkaSmRcS6BLJBpmopCSpDbcSlETgF8PxFYSlH
/7ZPIGFY4aJkNYhlLBDWvCezV7vS+42AG0cZK+nySFCx17TSR2HFQ+NPm3dHwKn+m52oOXWWPEz2
0NOZXh0NmstcP85AquC+vuiv+FqZSbbfOcn01yRWxVv6wKUo4NbatQ8dtohLvdrXCueWLlA5LCzS
KlxMyRui9y4PYmFti3+gKxk5LYo8N58RqeAFAlXCDtAWP+BpGHOsFnIHEOL264G49QUpp9bLksyZ
USnXRXecRRo9Nrrr3d5hnYlRnc7iYFnwIQHigviyZQGbAEKDNXb+7I9ld35y9/IY27bFxu7v86et
/mZce79lWNyA1Q1xFp3xbxN7yHUNxl3KRK5aurkBx1DoAXGykTzjeQx++zBnDhkQ0Z9W3dz8TmTr
+ajXR78EW6M5JnaVZi7QYu2vVy9w7SrZ0ez/iuAVffiHdVZpcf8iKoysQftI+vXqfFAF+9ciCVxU
ykKLrGYCV37hmbU0U++2WWqt9IprUBXQOAxtkqtFqjiRkUmRS9o+XypLB0CHUhOBuz1SfLsBB2kY
7QpymyghHksZ3ek10ChEZImL9CJ+UzBVbvotEItDe8Ki/+wL5rK8f06gp3ihoNbVEPjirR292tT8
8OfE22gmLHc4eGFEuts90KQtFa8M/Zq1RnApOiMqUNY6CnF+dEDxr6uwHIyGVLflVeU5UqP+FMwI
TTQCzMAIPm/QHJy4dutEPMVShMl6PDgPSPTbkhIyNtUo+09R0LSYEJAp2JcjkIaqshgOxxqlfwUP
0mjl6XVICzS1E4+r1p/F2ibVSyGHtePFq4x1uOEYJpDbv705xN5/VeLZQINK7nk0+gGt9EKy3q+9
zfqBSn1Q7fV4PUw5RtyxJ2fs0MGKNd/Rn5rDk6IhY/sv93t59G4v4fras/TGIeLRuuGI5DRSMhxh
rdPIQro1KB+Q1+iz/1kTmxJplNePvz2UP4sDdH8H7XfPrDa+yqC+tOi/+AhWyl5tgy0BSHN6m44v
8YAfoLvgsBzHlOo84bFwWrD6QtRcQBwWNmWoTZfSayT0GUb85fuJd6RnS/TXTVhkWyfoaXbqVUDv
p/BBqvWlBb2DpGfnyaKhwybj31Hy7yGyWTQki6GMj2fXvxINpaOsOl2ixXoaLVxgY3jjh/RMuWmK
Exn160brD4rBHVO9Han76xDLv8yGPVj4FymC8V+OkCh0QOI3ziwe0DZnhq+QKzQzzib9wiGCdgOe
gUdaPEZJtaV/gEeg96WgvP7jW1a1Q5xD1so+cWJgIN7kDKRDRwT/cJYCOv15YRJw30eQq20DL2LL
3Pqe3tAld4vJtHto92kONSEHEW6YzZT+v1eEBNbWf/MsFM5VzXloSnk7mfil1hz6LrXKRui6tVwr
8TXxocEHBl6tG3GiHsCsol62BtXAUufOYyYnXEZHMqfaC0ShF9CxWgGYDuqMqs+HjBoaCYCLR9Ws
oaxxq12gUf28PGv+brIOrUljBTr7EcZ0jwFULRXrNY0q/uoS95G8MTIQM0TWBiSGhQjg1L1sNZu2
pIaBonBRIPgaU8qy/eTXjqQR9cutFiOfQQuvrwnq5c+tjkDKvpcysMJVcihd0Ld/SQZAQyhGX7rS
/vkZz6bcPB4+pUijvsF/r9MGQABmKZqBGYgcvbHTG4vu4JQVZpEjOlXoPj7yQZtCD4BBluz25bHc
I7dr62oPDRz7bwzcPaGSbTlvVhhKuicSxl4uuCI2LRWSC8zUCwsilu60KahSYdwQV7YcYJI4UmxF
W19XVunvWXPOJYeolJ+mkkf/cMTM3rGpOc4mgnCgiLLe7EN3cBfc8z1Is+Wc8BCyqdk8FPMnQScn
IN8z8YPQYYj/IBpxwnEcSfOclIzHO75Ko9kPvddpAk+Gw5etSgF0cgvqpoimiYLvMJ4yUmtQuZJA
Y+miw0lp4k7W6rW8BB8g6Qc1+e0mrE6oNqTNgaBgeoEdZj4O6NOoVzFPeed2d/7j3w3MTtNKni9K
aWuodDDhSw0oR5DeQr/jZTaUaOCoZv/y2Pw9IaOqKlf4aIpAVveRyvthB7MXMf7LI5ERVA0dhb8Q
Zfa63wyqZccMRumBnVsSc4NaOCqN96/T6Lg3pMvfC+fBZnRLZ5kp2BN3majhtRrChmbtz8c7x3fo
xJ07GJg9usTmLj45c8M2HaEyfvjHjRA1cF+xWThcM+AKyC/oTKCqo+5fQqsKPtMlbh05dODLuvY5
5a0KSuTvNwgjFwMEfYPMaEh2EoI/ICwQwhYMZeQyT/6hdhodZPvtGsKjiolUPY8BjN2H3NRA0UwD
5OruM0HzjIVeqMUhPDE+pKCyTsnkX7XZNWUdTbl7NwVsxaUYzdLTUzKTt52H3iu8dOhI/DsOVWma
rVyUZlClO7cUcA0b3X4SYDZDM0RfcEMhSMzWrqqET5aa5DXl6+LGPy5qEZNIcgegks6hVJFWZtks
yH9AqTy4vy4XSeQ0wJ+z50+cPTyv4lGpfiGJ1b449hwb+tu8Hiqh4aqmlmesLcyC5nJ93K+UNMfE
iqafV2VFRbpQNCqEYbNv/AD+ujuKMv1uq+tj73wd9OrPBZ02ptAw4ZYIqqzp0Wjd9wmh+CIzzFqV
PRANfSQR/Gs3LQ1kmnpjMJPDcVqJZtnagKjUvFcfgouP/KXix9DvQF3Nt0YPJdwUYbcR4qOgRnWP
xTD81lvpEUQTfkhssXkMgfV40qnoZZ8IgX6lPetuIUeOXSNNSJdoabintIAdZzfqt2rPNMHAaPNy
DlWZJivr/61sXRD5bT23NPF5xqmSAn5fqXxYWDehKDded2eGlhy+vzYUG4zAnHVJDRDw4Dh5gfAk
U0oVRGSDpDqg7cV7bRHEjqavn4WJHaQYvEnnd6F/Wf5goEriTuXCF/SM7BkDfU6Ra8Vdg//MyR3o
9loTSst5D6IL4qdB0ZLcWHlkXTLE7EB6Q2fj/wvcsdBWAGD1W/A4uhZd3a3ljUq9cjCgzDW4i5yv
0XJyGGXSi3joB+vE/1fP/NDDsR8YVLITlqgeBJAiEgO9BZQfD4zG7ikvepcqxpz1tjxhWfqrFuhg
2ljRYwRB3ZjweF5b4R+UdrxUq+ZIvExZK/oG2A7BXUH/SnKHCC2HnGLtiGjxwAOfeeWAShEu1F7n
p2nN2tnby+7V06z5g9LAOknAKjDZPbbU9BGvjDPbH4HwdwWip2c0a23UUnKOzqNYMtx6M0UluyDh
y3vWlOkIFBkICcNLgcyXHATdPH+XkiS9SwBs/PjteTFIFPqf0FZSvhnPNTbxH1XCX/+/3Tth2X+m
LVaGr+AYdd9/aMha9QtJlBgjQcHpNMvJeaIJtVImuo9ceeorpAc64+e47fqXp1EDjh+k8u3p8S2f
G+Wyb+mtcxiJAyzmmeFI/13e57pVWf4J5bjp7b5j107hlQQpfrGA79WKr4Bn9rhuC7mR/3Bh/ME+
XKnEYHHP00uWdq+3YopJsf+p8HYhR4O2c3uNL5gDDPfC8gt6MDXGpb36PEWqB/fV54fELrA1ezrx
f0CWnRAL21cbkTE6qqEdbPF6waGMV2HR062g8n9FPdxGuPcw2wTa5xbvY+L96UtDT5w2Bit1dpZa
7Kh87dO6ty4x2fLyGqYFvJFYaSJtbGKA8xp0jkll7VlODTKxjZjsCS51w9JfUxylnBbQirGOfrxb
B+VeSn5QCCgzm5GdtoEcu9BJ326sCGV+nMDm94NQ0pI4kDcGRPgMMydYZ3h16n5wEoNRaDXGS2ah
536iOMTFSDeUEs8xhozu0SQh8dgMC+pvKcd3KYtRLjHE8BUzZ8yCNKwQMkmhl/EWkZchbnJt/xdi
fP1A3s88oPDg4Q7x1CVIl816bd+JbTbJAVIVQcZ+mgX0xsBXxC8ErBoCEUG34IMArMGOxAmD9KFC
jUGwLHFNeh5CZnfSF+KOPRi9j9ej4OzxL8KVsSFMxOluKhi/1aVtmqgWnyp8q4CiGzVe8p4RLZGc
f2n2UYAJuaGsR+MYqSKKezS80kNdZe3yov6vXWy38a1A1D0xhPCUfa4RdwIIPEKim+9YmtyiJsIR
WFqmo5gBv+oxc7DMoxmZh0U0hlzd921isUj81S339LKqPaPEco7snRf0ox+AHPS1g5Hmhk6AAUFX
9F8wwNwMIxd23IATgsdM85cgL/GNfF8anEIAbk/7ZHsr7Y1AasTRxtONfyab5HRCkq2Btp0DxyGU
IFOHiiP+lQ2fUcM4gsnomby/pjanH4pVkMPtP6/rDvlru2026hDxad9hMgju0ywEk6Uba0+HkhKY
iDZS1TJI/uCl46hSDCrF1nT62/kqlyUKRJOIgf6ow+9Eiks5DCL/cYHitFaS+HhuJ3uBsU5uYGdV
d04h59tecPzimHvQzBfs6KPdw/kKs5FhkRxA1kG/MV/a8u9x9VMVUAiegmpWE0Sqtq3gujZNKor0
tpFtEw3TndStaSY6zEQi0pvwihmgClj28pYhr9fNvwJjwJydCF4KvUAqklu3Jt/MwayQPa757bhy
EM4/luWrL0tnb3GHjCTJrR9agXpkdwrwglB3pZ8TuuuqM5LgVn/zMEe1fJNwDhI19Il6FaPDVie3
dYfTmmMfSIYjIT9ca6Hjomf3ETsw+SidzuK/1i1OBkfmmQSMxBvf4X9iO7D/TZKdl+OOm/owAkd7
awRG1dC2DSMgr+wqhjTPUOJbM5o46R1foyIM4v9W8f2pXRYiZ1kmTYuCLQOmv1ppZxElqJkMvcNJ
uhWXq7XUTo1EvUcqlt0cUC4eJobMCzSF8dSTAoTbs1D93oqu24nRyUdU5/FCrUFcEeG37qRSuQdy
toIcewCo6pI9LwiiAOSvqz/+tIoNHcHQsVLQR3geHjqfD3Ob9sbJGSxc2w2ua5dYIAWAuuSIknNf
gUFUxWMNZgNok3RCL/5mkyhNnlrdFSvh6Mt0xRucYpAQpMGgRyFWiEOpvuPsf97LbHr0tRfn+d87
Vax57TN8xCRkWtHakjiumBZz8Ec0H4deMARuQNpPrONChvljz52Ebnn1X6AXo+z23x8acv19eP8B
i8IqVypiAroXK3id1K7DNsYGG2yHDZab/AgkNbL4uy7qkXlIkeJ2oREvHwZdP0e2+Duuh7Y/Rold
cNgdzqHH59G5LVylONibc5Oe2WzTV9XI+vR5XpRUl0PijZWXvw5HK4EpWOLDlGL51MCfAr6D9OUY
hL52G/Fhm7PwWnFa36QB4MQqw4OYlbTJ0VyC/gN8v+pLildrAvJ7Y4gKYQStU4m93pv84d4Eni39
sRprV7j/nvUsWLf/PWqExdiMpS8HGvZFU2r1STl26026fOsYUG3AJ9uHWymmP2bZw1MvudjJjhuY
2a3R7WRd9agFqPodCs6RHDXSO04NpEjEh7CoB3OfxYPEYnqLisuqnBF06WVg7Z/cRDKUuN/jHWwt
nT9S88OtQXiOU+IHU7Qz1PgjpbGZIN3PyuDfGHMuRaOKDaxp9gNiyEMRoREk2wPuWzIwT29Zx0Ba
EKbmJ5B3JQrVuEAFYkmArNOGMzEsHgse8SddkSyMf8wU2fCZ/iJzIwRjlcowQ2yL3K4p9MggtXeZ
bY3m3kDnzd/slomTG3+54aegfx35/AN7/SjLWyLNjFvthd2wTV2F9n8jqQoXtIp6k9j6Wt4hUWx3
kKYorfrT2wiNDa8oK1ngW9Yl0mjp4IZ60ZMYyEFcyuMPrg6nRVPHLYJnLYpXwXLCnXY0oHYv747F
XFMdTADyHe5EKmxzW9/lXB7I8yBDs1ygA/W4NMj3TsmJasVqBXgBPO727o7/R3VdmG0mR8TZkNVf
y73s0gkC/AXrR8YUI7bAD7dvL9qRcqYkFQv4/aY4yMl0gNiH8lgwbz2+jI6b4qd3blR6v4qPdZfv
Rl0Lr58pzYwtnnqmyV513uRKIQuaRANK2WoPzPiAmhIcy12m56R3mydAyvkFAk+DRlC3nX7PkteU
gA+QwVf+Dk05Fj+oGfQNRMCXWmOVeJ6Z/7xRSs/57dqq0vXT713MVuNvHVjTsp60A/IVjnQ0QzF/
qRRIRBmGhos+MiFfydAqhl2afiCsHrrbUy+n4iZ1xs3lzDJDMN95I2VBGvwOwnbipXAfAdXwrpzu
ggu4IhRAY7Ib/cRwta1prcQbZTj5q79p+5g5sirsshEeo1rs4AdD+D4n0V8oL/u89s7DLqkCCDHv
cXC9anDondiXndxZqsvtAuwYrIXaGGREjIupuR9cNbH5auOgXKhJdtgDthts1oLc1HydzF/GqtVt
uUv7+cQ37AupsQXyTDOHna42aLaYzRpW20kcaN8D0wnMk+f/kfPBHKJbTnnIwUCFejs3V5rSHcmI
uerwdL68/gFtGzfG/3395zFLSi2x1IxjtmT7zrEsphkV4U0CjQ/kkwsiqbxnfJNWYZLQUMDNwJky
0Z5AzbG6Wo54j4dTvujOHI55zG7HlKVRhIvzt9YcGZxW7MJ+UMdjXvsAO/5drie6atEmTWJPwZPM
QT/Ii8T+XcxHzcNGk9Kr7RWbQH+jcHfekiAefSj9CxkU/edTH0uUqZFYiXP4x8/4lU6koAzOYEoq
frmWtUEXTj9RyozwVoiFszsxjBi8HPqJdz/HnVW/v8ZE2SQ6FvNdx8y9IrwhYcCLMtXALFvWyfTh
WIqV88aydwo9M+bMzyaeVjPnpTy1JBV1LBLCK9E2CtQ63b5arU2++NbiHRfcXHlvLrRjV+u4PAWd
lFb1S22xGkVngn16dDHWaC+ao/a+9Qph7CY5UNeQN+gh35ZqlnmQ+mHcstsj+aE4qLJQnbIdunxB
WRe/t3aVqQLeGM5LtWhuI5jcY0Pl1iXYdR6c6MKpYZ1HMHE+wUAeqCaZYpFR6wCqbJNjHrYRe6m/
6CGUWahXzx0YbFFxTmdB3akq6R0bGw9SgzWY12mcWCcEHtNKr7KQpIqsz800s9n7mWaakrPG73YO
apZz6Hrp/U9Fitk4F40LL05EBGHtafP7rISq3AifychrF+x5XyvBzP/7j4efNiyJZGslQRGx+C4y
wSUp7Ld1C6/ntFNpjo1+UNhNFdwv3xIz0uW84UxWVvu9pVORtSxQkn4ozKl2QjZVs+UqcgPTGEc0
IxoHB0v+n3zaS/nSGuFIQz5O4KIZJHf3VXgSsSfOTiOCbGdx3vgbpEQ5JrxasLfldXwOKRrPv/ni
XmrlupWB6b+VhfxGz5pTIGlqNGOOzFPUW08b7F8EXk6IAYKCG+y+WBu8pKlRQz9MAspbcVGJ2125
p3lwe3Zp4anRn7sj6y0EPA+sH1cOVP1fsuGlG6H9IOMTkxoL3ZSg4D+ncsRjx9XiETOJPA/FRkaE
nzKz3SDvwbudYdEZ0NGlCfo16lHyBzAwkPWjHEwW084ivmWrN+o7vr7NMGHqNHSdgPRmr0HgkyfO
+QzvBSxie6yBjofbeTJfQy32LCFYP0WAeJPXMEcQiOrUYb5mY90wYhHAAqehY1/90+g/N3mpVuTJ
PN3bwJcrH1i5rKpFJy2dGelOBlOwjArnEZCksiIZ0dhBMAo4Gvrv0045/3tbd8NHeALQSz6+kzRS
TnSzqjQrzUX6it/VOvW7MwWrOEp31WGEiB+j5cJh1S8n52Vz+QDlA2wF0PdwnVS37sA3gzHaaVxa
S8Pg3UGBNNvIyZzjjmRg38BhA3FqN0xDkwQ+mw0Zf+XUxITX2ZbWV9B9jnIfTO8lzMY43mwzAYtU
CkDg4oDpfzCFh+lxc4GAWJLO+btqotkaHdxbhdI70j9rtiNwFxYp7x2qc+gA+vZWXZjE/T7hhzDm
M5f4L5Qn/pTUszeZgxNgDjv3zukhbpvy98k5vpKL2UYB5MUCZEVRfXp6qTYllUFoAbsCSBXO2ivl
Bw3lmH2iVAwZnPptkInp3xhEVeg1MSSxBIZPYD+2LOh0zkuHu/of63uvjaNI+WQaNqpK7WdB/8I+
zWR9/bytG4zCMcqU5s0EaOxrPWXuIkiQQfMVqRarRp/FKRkhX68sPOdNe04YoPNU3FSf0gT0dl4L
LwNts1iV9YZ5bWtRca3G1tx5+/MhEXQqP4XtSdJ0s7Yhiel+CrmkS4Hi71ROd6DIkOJnXACU/xs5
2+ZgID8ZqBiVS0qAaOm3xKKcO8VhGAvpMJ50iJe5DQSXHrMSCol9MAlFfWKKfvr681KLDoSYyrft
vLPL31cNZudRnD4lDqCE5IPMK1JC79MnXK3l70vR1AwUvU9OG2LLsnBjkNAdeaCQhgBaUH+0oWS2
CmKqjiRv66eYEk2+fq8bENWZswt7Yte9MA0rWrYSUH9CfCHFozNILpEAEqZFul0qm4/FppAxiFsM
l/AqZoMdishzisVz0hjR03Vq2m6V+RJ0Z/+nA3XPyl4s+5WCrqurbv0b2/KxvBJLvb5o1HolxTtL
fSEQ/+3qNQ5BwKfM3JnpD4Fcz72xl6/xRtjIF9b55GzNe8dmEOtYBi6xOugWsU4EoQ3jynZL/l19
454YqvhXsdnuR3hFHqVnSWgLlcFD7WEWNLZT+PQwZF+252TT134NJs1zWnPxTyaxLQlj9oe9++PV
8nHNiTxAtBB1Uhp39xpzntQjoc1JKoX7O87y1WdDmXQvcQQfmWfsCOeAwM/aduMO5uFT1MopPYvD
OQ/+5ek598jC2MYXLcHbXOV+3fCybDSxWXy0LVCvFf5eHo8ZQmazG6QglLrO4hPTH7pJGnLgMB5z
pRB3mN3D+FJCxYO9lqF0QWInBcE1qdpjnyFR/gA0259/4szRGddLBpekIY0UCiXqaTo+aYv1jP2w
JeuwVTvdNfj8DMQpset+MFYFfrrEDRNdhPU8XBCh469rHmQQu+3suA6LQqVkwl8afpUmtuV+jiaQ
xnKQuCgxt6Cj9y2v8RFf5BM0h/T0ZTZZiTsR2t/Rz1SWN80Tjz5PE9t8MX0rECdMdQiQ+LbGpGcq
mvyHChg2u4sqYNXaRnE1CFoHoOR9yBLeZ8KdnNWFGezx0ubAcSslN7t74/J6VmCpie2f4iFA19ty
Km2oL7Vc04Rk4c3wYCVCjYaBguz5+EiojwCBvasmsoG37kwd1ETSVZXP3ksbpA7u5LFz+T2HqNbZ
f8P/LAdge0ycn8DABx20Tfj14Rcm3EoMn5x0yjUCq34Cls/L98b1Rdb4nZapF++FrqPo1ZA+xfjL
BdI0eGZBG14hPhbs8px6lCD/vOIkqOpiq2vqLtOVbtmd4KUk6mas0dXmJLjSGGhsxmkBvBvU12HM
rqBGGZPK1z+cRqsQ6NBu+hxzowL9OhW+VMlP4z+UByy79DFaG37z1fnkIBlk4ldDbNU9xMBokveL
H2TdSwkI2S/Cdyks0xKVauVI8cApTMEQWKtE27qyUNCIYBhrf2HYYCtWirOsMoBJ3zuv0m97NAiC
CEOBa/BQGZs1ugfeMlh9pOmkEinnaYeBKQuQG3dSB7OFYZfsd1AuKrxEby+mNotISXLF7Pl165YB
2RmbOX6sXXGF0D149DiQo/5mt3vBL67tEkEhz+gvPe+k9+SIGfgXTWX46C+VZtE04ucNGciz+GMT
njsGnOwT5kYi16HiiqCKmRDeskE03gnm2SMdvpUx+20+EEcbdoF7yLzrog6vn+WmqEUVpJQzZhFo
G4gLELIYHj1BIYlRGbno6pQcj85VLI5XE6KuOSBfmIMJBenKxxCskq0kZo7ICaEPuiNF9EPSgyui
Wcvtya/qqPYcpDTJVvT8IaAW9l82G7SzeyC4Phh/qLFYOD8JemG/4R8mnZQCA5sUOrjgjRk/K0iu
eZBBtT1zGFXXXRGOs+Q9b60rOXlqwu0GeMFUh4Hz3h51T+ht36xG8AybH+/756D2CbvQiYHlh8HW
DsHNfnQJgcELBxIzpNu+8BDh2zd/8War5uHo/+9khPoXSyWpazq0vZx8K+SYspKOuG9UO3Ae44Nk
T//9cgUA6CXlOnNcuZ5SJxAN0uT4Qph7RcxsJkBmUz4d2SOKJqA+vzsjxc1jJvaOac9Mtgq0KLAo
jOS1tzg9+yFikjpXBUQjnvJ5Gprjq1UVEbXgbkINmNYC4jJg4Efzat684bqZBBiLvXNxc5osSusB
QGtwvwYsM7nMDFp1HC1rwavNLt7nDQ/IZ0p64DAUqnNHNgVONQyVdF6X4u12bBo8orMS9ycublvU
I0zYUM/MnGssKh1Jo/MKRd7rBMJJ6sN1rn2YLlOSJ+ENdXX5efiZFuLlG+8TsC1zunoSal2LSLNR
5sD0Tblv3ngp3L4+hMFAjOSd0/sRCz3is3LtBJCqlGR6OFM9ozCGo+/8/BTikechKvLGdSXP2odf
kB3BAZLWUkIUy52uTNR7OWnvoP9+UgrFt4Ps5ApclJr6+pnSl04TPhsHQSxBiQpGvcTAXvpSO/jQ
KnrwQ9LKHc2Y3o+D6J+M0qvpTkkhcBgSZSzVNMR6V6hImXIO4bZGAqTGn7dALRhxOrUmw21BwZKy
c7Hfvqcx+LI9agBrvCeSwz8bwd3Cxpeudm1tJ/EyAl5B7Ef4FJXt/zqbxr2qglyJQT/HqoG5vjIl
DOlEiSm/f0B6NCW479Pl5HPzaaR7HxZcJ/PcMxsidTOoWOZR10gGkKOmN/dvh8cL/cnMbYqDLRkd
VwHPgt4PLajv29tx/xpFKYNBWhwBz9kNYSps9gWiVxlKT+CT6rW/cY6eL68XtLf1vvJKUaVkas2E
ebZpmrrcwMfk7YSQW84aRnPlZVOxgGqVzLWOBVvNN4jLAXchiYpFZrWerdhLwzgyZBRMjq88VgGR
pTW/FUZFlNM0fC0rZ3qjKtbOV81g2gpn/qMvAhZYUxMfi3TOtqDDUSKqjmxO98fB1mP4oxRvloQL
Ks0FJotrLdugMDphyX484tQE6H3bTkeTUSYc1rsdvWbKinq16Ddhqyy7lLg6XTSNBb2Y8YAGLG1p
r20nbMCfldidF+mIAQmL+/GYi7GdI9+DldRycsdTLyngSarNDuygrFQQZcil1pHBvG2vDFzKNIS7
GBAEZpS6+YDLpQy+0yJyy/hRpmvLQkM7NvxRyvHqsBf4Ucw4o2gC+oEfWWjpuARWvHce/qQsEj/2
O4gLY738C0Ml4zXTcF4G4vjrUa9oybh+aON7OXoe24BD97CWUKymmyoQ7DGGiOtTNAz7RUjijqxd
Bq8FZDd1ui3jWoZ3JqZoHQfKwAFyF/fsxYrLXMP2n2tHbJuzegzE4W1borOWnQxAl3zek78FCD6c
wwQ2yf+wkrChqvXjW6x/JnXXUUn5IULpoUnznDA6GBJ1D+G2yqaS2AM3ASkeQpH4M4Cqk8yYBVYQ
JlVyEbAZ+qT7UO1G3r6Di8NWudgci6vqaaja13SazXFgs7uVH2MruqPbWvX0PXWfUGKgcv4DdY9e
yxSPz+tGxqWWveiBWFZhszITL3xWO9Da6hJhdIinSUWRQ0RLXSctkHsZCcce+jeqSw9c+icGSHJZ
iCgiT8psjVu/XhUSMNt5OyyetlmNurSe8uvYFjoYukbl/mR57r/yD/cZr1vvfiO+y8hkXchKHQJY
3XRq51qjZ3JGeSmB4O23e1BGREII4fdUijSk9ozFSQWYXMd3z5/fMhl1icg5kom+AxcCkH5UDScJ
ZGJtyZ9CFenw7nz2HGtLEsodFyGuHGSbEyW1i+nHrFfjrojwNx1Wkyxge5RIAFxEhvQMop14Ikqq
ZD4u5WOrhlt1FFp3fYfjqRFsorBvo7pPc6GnpyFZ8VpHihmdGEAUKKDG3lvuzJKEdbAPGehTp9fM
X5pvVpGd39YGRg5P26jUo1QxoFCkrR2xARwmmWRcnbcmF69t40H0b/gKiESoG4k/SRqiC2byEEJI
b95+MRYdIyabNOyvkD843ErKCT/LmYZPTsZ28Ne4ak5GYUcy80h9RUvmI7fNjyEViduYumMorKaM
tR28HllTPAimwbxlJGGwqZZKKLeaeFFJ53yGGBhZQXfqInlJq901XM2UbsN2dsV5opZhAVKNyH4C
J4XPZEAoX022KT32t9kCDcbIAkSqMBgOgwaEJGPZDSL2oDbuz6r0W/3ZVjZfQvMeSSUj+o+KaI7T
gTM3oi7+pzeJshpHn2JGtkaFiy73y2bjmsXwTYE9pNMhQghf4Htqd8fV92Kiay3Pvhofay1ezcYJ
Z1ud0dG57/qCJn7pQr2C03ZH1hGB/NQTR2qemq2ARqO9iwe/iqLmdtXxTtEpqGqek760lbzscMQR
7+NI9LqG8maBXLb9JFhwmZ3w+1Lg2s/Acx+x8nNJpYkrEFQoBmnFkyRiPDlNvYO8T1bb6DmqxCGn
25rJGm5wDoNxMzqSXQkV79lKSRg/uTtf7u7NcfJqoDQeGGKhqbYNrK4vWyWo+JCNtMJl1+St9J5P
NB3JdRMJaM9FdkoyWRUBMHHjK6x8yVr7+E8i1Cij9nf4JvGy3Rz6lgStT38aVyzn8llVZy7JqxoU
+j/kBkY2tnA63F45K1NPDu6i8rrkhi4xe8mYh2NOEyEwzLu9A5GRflTV8yfo9Dk7T595fHLjicNl
Hh8ypkXA2saB096SIuZosV+Lio3ihrfBvZqHX4vyAK5VnvUlQn+4lGl6s6Oj50Nh1Al6FveJZPGT
OeIKy09WLX/Tir5mfK8i3wq+WOf4J3EOHR93oVD0ExGf/u5+7RlQtTIGTHcJSjn122+Qy63Zp1ge
hCex9opQsw6+C/Esggl6HQbn0DV2FcetjXUkDbtTVot5tpCC5SzokrNlZXcrWQHLDtxKYrCP/Fq5
oyjGihvZ7HrglrzwT6igNQdK60zEJ4IrCR5OKHkCPETTFNgLErFUJK6/AqA7ji34eJ+CkpuIrIgz
IEUENC/HSBteCgpkwTM2bB3pq0Tl1Qkno66m9Z/8LcM9hdAIeZl3kuurXrXp6UpmunglQ8ad4dB/
aT1g+mx3tMQ8a6dx05RH1OnbOpDf9sz0yF3oWL6LrjwrvlniJl8E3QIJbzuDlR8C8HeLk2SId2Pm
u5LlYqU5tb89nvbo+2ffJGkQAuhCaiI36T5WOpuYnzeZjjt7oG/HFxkQKzmqzrrD7x48Mk8W6/30
vtw1ZcyEFfQszKB8MoHb7ogjUgjcCKklry1HetbkY7QO1KKRpDjUQ3w/ljHLkxakPkHSgvsdJPab
XHkQgFpLdgE9nwpDCduqSlZTdzP34MxNkDXYujECR3Y5jZBEUe+/inJiW2AiujDE1o1VwfkPVn9n
4XnyEJWO4YRB8seifYiq5jXyPfnV2E5d8ldVqxKWcurpovNpvL3J+tEc5X5wK0H84/rxL6evHALc
/jzL6tNLrpOgQ2txBXfpn2mTD79GmqOQwqhuU0eTjpnbBmllbMK6knNs5anzBqb12QCs7cggxhcu
ouwVisIkhFeqiSW5c6fWR7/hdenLoiidSHlZhVE2IgvNvk5A0Hld7mPUOYeHYbVPOIWoew8YEJRU
e4iJCPFXZA/B1r0AuX+SSo4m6Kmf4+7UDGs4VNagDyZTMYvVZzrPIyOTmC/QDpq3dIerVLP+3VvU
B3+8DjcZziKkmy+sa9Vc++Xbr+GDx7mmoc4B2XAQvlw109DV9HgRqGVa/dCei/6c1wZhFes0RRAw
TveUZCGgYTNo8JYnf3rd3NP3Jy76ZN57Q227/sAmmS+ddNWnc2/YIBMoRoKsppZlkil4QhEjafPB
FcIF/R5maOunqPjz+VoSW9KYkYDzmq7xJo+G8QMTRCmBQHNdFkQZwh6dDe+mkKw7nwu1PtkCtPEO
9U0bqUWIzgDCDtPzfMZYoHO4agNX3Dh3xLGceK5H4aR/ASLZVhHYGRkbl0tvYDVD+AXgRnHnbAEx
cvXq7ETg4qpR/9XZpu/5h1BicHpgtFskSniW/NC7aaOeDnZC0utVfpQ7YM5llC2t7Z41lze7sHpk
DOqyelYXUTeyFv6hmappf/i8wMltU6/3LZKtWgLZqa7RBRrZia1igIQ08FnbxBw9+bT1INJwqk13
Q0844XIrGfHkj7BAxn9KdFc+/xr+/SgVlqeqfORGcS/WxhYSxO53n565BOEMzFqJ6WuUOOdxrJ96
P+iCJ8gcAL4Ki+Uadm+YmYTAQEoTm/BYLTBRn/PvN0RMD9u//6+uuh7+ro+dlTErlrnITrLZvS8R
A4Pi45SA64O/RcLDcb3Xu1B+MnjlzkkJzLPEC2JCH5pUwyiCwOZNgx/A7FagELunlWYsc5IIbED7
CobSgr5Tlkycq3Wl5wH8n/jmwUoNCOsJCmLFH2pdjxwx4rqk+eFKpYD/CgwTVyUfRtlWgxvIo1Kb
yrLCt0t5acvomMDknPVVuGPuOusMOh9Yz+w9aJfQW42PBnQI53h/Co9MN+qP+RbKcjxFljYzOcNd
ZZGqZpiBaWrjr6MPw1FFLsGcXSvxzlrlXMehGDNvlJiekDi15r9kOQWWIWy/t1IkC7H+9572Wfs9
TuxFMq4IZjTdf6FlqjN/9zC3EeMMF1BybeZ038xFW+UiwrEkpnFZ13f0zyg+bJ+bBr4X9Javrn2D
8gsT/IGc9IskQUvtLHd9WRa3cGTQrKGJG+RnVtIDEPcsYgHsnl2JlXZanV+kJ1TEeQ9JjIywRfkA
8uHiTM9gZiBcGiuZX686d+LEmUq77fZvy6sr9LTEaedQvq2pMNMA98h8Dr7gPJ1snJinehz5w0A+
XOQuJ6iCQ15h88EgXrAmEbOIFveLNHGtvzEme7OlK/Ohf4YxXw8LF0HimMvPjFQ4018zQU5+sboU
RwMjaagB3LF+QXm4EIW/xYmW74UekTTa9Ww4inUbmn9NShfclOZkjBfaFWLuIM0/fhUTHwGp5FIK
ApdC3seKmQCuLQ/Bx/5mrmCw/YwkT2zUuQmTo4VfbAnhefw694vuB7igKon787hYDzMe4BkT6IHn
fBx+fFaIE4SFgzM+ZtP9RKUcqEmrYlca7h8ngdbb67OqZ/MA5QdXvQDOb1/kRlmjSj3Xt7gjID68
AMIbS84dL7flAxA93il/rf8sSHPdzJ8a8eIPf2N7F3L/hKcpAMfrp7SuNYfL8sPvQFJ3FpG3wvpU
vh1dGgNnhExrE4qeD3d+yv9zYUSgLYPNmM4Xv/gVjMbkKU+IiRtAf0ZEAMLo1vI8O9hU6UyJ/PeP
CC49RcoBpNO1rQHLclta0TB519ymwnobbR0ve3HZQObOsERN2ZuDNyHZBlgLH7O8YcO6eiqGJJMJ
sd6X7NBaUQf6FtZckvlZYn9JMfWwubTTgykY/stF+ouqs5c/yWcGESBrXIfQnpZ17qV9cV074hNQ
naGV8r5AWWq/KFOyKUEypiCb1aD3l8f35Y5bwdKuEog3k3TYtMkRRnrlFbRFLKe+AlctLHMmfT35
HemNTw6ZY99dnr0dQ4fikaUV9QRxHHWhaAUZ6w3amBmvohIuuj2ps/g3nmpNtRkW13teDp+0fVYx
tnD3dwVSPfVa3NqDeFKZgOYPzR2qX5c1itUBuysHJ4uU2XKOScse301fB1S1sNa3Tzu2QE49vPSi
ggk/4zcGfi9SV1il5+zciBtkjg5PtRtk52htOUtREIrs1YTd2wCiQlJPZ24Ve2YsY4MxGTcG9Gg6
kb6f4kxwFFt3y5owOGk7/IGC7Ctj5scMjE0K6o2SNRRHbxucxsDBPWbOP6oHyzLmfD56C2ofBbie
c+ZGU0fVFfIKpdri8vgmzHUS6JBd3/ZftSALkNBb84w0cGUottGCHyQoU/0uRRga88dSw8dlf7XI
crKIn5xiaPoha7wvhmGrQfhHZVX8qB9Nz6Y3ZfsagWWO81fXAP9ay5IWMUCGk4E+LGIvxsG5b0tS
QPeoYA4k25SEIN+q8gFceeQZLX9WOfmqVkYd0oFda4CjWihg+Rq/c1ZmRP0w940smpafDI4wHr+c
0rU5sPSZ81X8wTi9tP62wi+yD/FXzzLr2geTYjHXYCCZcofN6AQtougu5OxEsCmI8lG1Ye65sbvj
35fiHjTxhaoZ8B+ORQMr6cvV5ntNw7p0mNEYt0nSASpK7MqBTuw4tG2B/xZgERrLwin/vkYBmt5K
DHrtbqOESUeyC6F1iMu7Y1E9BjTYPCAibYA1MNnDim+cwSsK/oW4Fpud0+DpvA+KdGovn8p5efpM
dqW6e3fqamSjh1lp8dXBJ420f7JOYZTAgo/fOf1brRAq5Wr+/D7Z+yW2eiB2RmJP/02rk074H65R
kHHqRr1yNUWhXLpF8gtRc9kjc8/WfgQ+/rRMv+OJ5EJAQxXT13ERzs3SagkgWAhDVJKc/n9QxHaC
2GBeypmVON/KdU+NZ+cXyGzDAqROnFUw8qaytACe86mLYoAt0gTn+0g1vtwRWwmckgVENksBdUFL
kA9GjBciyhSYsiPdppdljz7+htEkcjiWEWYfe+mGGWCmWRY0ZXBV194Txwhp8z6TbPk5LQ4+LpUH
TvNrqMgWW15bWtsWgMESCCj/Cnmy6SEXp4UoyR4gIvGpAEchBSbLbPSVFEXS3AxPeFeykM7/AfGR
s8BNjO0OALISFvM68J6PIsixqLEGIHXg4CRPuskg780N6z3p+BnNlIIQQDAUuoSsnKN99AYxw/p+
TnV8OdZUVANiRZf75LKtN/Rfz1AamBotFB3koBj21mdRMBTD7tby3aj4uCtbFkXIDZKjf+idTF/8
ZvA3F2fSAEBrdtODQ//X4UNxC5eR5IY2xaA9BXAHbwunFBtnEW8if/uIPUxwVCuMIkUNq9csPm3x
uw59oG3ccmba/tK2nlkCeNkFAIIdM6WHhjFBIFhJIzqXpn9u36VvvQmX4nikzzgspu+JNpTKKvNq
xDlHc5G3W2bz64cXlVYs8AkEDelRTa8cIIM5Id/iZqYe5j+McxsQDZml0II+w29meM4sqq2nu2h5
M5so6xuy5b1GLtHI07ILi9zcb7ulh4mtLyjvQj+tAp9zri2s9dSaOgFEYQMgTlxvztRNgwYCaXT0
DYeYKU6QNX99XwlMvRoyZJpJOnfjqaMI6drwcScMxJj+PMgr9P+rDTipKf2jLhsaRJecJxbnJEjs
uPf/IoM7arMMkybLmdbeeTxzz3ta7B75j/Lsk9zEYf3dfKBZq2EnuElI+C++j9bo6OZzlMqEn2u/
sO+uP2GRy0RcsOVkG14ZBWPQ0Ma75xX5Oz8Pa2zRP4x4Ivob1hng1qQ59zgNT53lnZ1uO9F5JFLF
21hIfrThP3ubakz+eablumBc0rP/1ZZDltDqwVBA9Us7jFn9DIldfZmojjvCkrrPAHYhQOUosXHJ
eyxSYetW+BRh3/O6FYob+vvsYcXAuGHWsDKP1CSq+jlqgBkBvIZQOXZplq1cyah+0n1Gr+1zryUf
LRXBd/gcn9Vm1qOSSxpyOcLuDjIMmryauluFkyVJsuwYmRQhXsSxgLuzgxWZXhiKATFMtCJP+iHX
49E/kBan7ALNVL7NW2CR3Zm9mxMBZVjbbBeSyhtSsqvDEOmGKo0Ri83lzj3cd21kUALcPHTLe+M2
cw5hYgWFr5oKJhMKu34nGBUy8oGIjIdD/oQPdqsuxOgYtcYD71XEwMKyJ4QTSKNQaVg0QRdWIfUq
PnTf1XfqsNzkNWrK6exlKAbxtU2ZQuBhNW1+7PzZwSk06QwgZ2FvySt6OsItxFY6CklnfrRmwUlE
HknICCshzBBj0CKwdKvzaaO03lE86eGBCM6LuPiyo4MAFMmJkIhpzgZjofKUUIlHUQ2+L+IgIbtA
IwdtzpPZaoW2d+8zd+LvM0u/v8tE7WhZT/rf8D+nCkhN/fL4I4OwT6xHvGdO8/FD9KaaEg1LT4Re
uBzzbSBMctC1Cfprg5AEmErrTyu5UppEQHNMjUwD1PpgNG8qqhzAxt5QgwKjfSGkP10karKAOOSA
zC5qdMfyPFBQK11Dg+6dxmXKZVGKDgL8rF2c2BQcWsJYEIphniTHhzIpVIjBkg/po03tdce4d2pe
ZLH9Z/Nw1R9ke9MPJajzXoUmJO3flJmn3VK6zplSLKZPF3Hz+y3PWCyxa1Op4m16RAz3fdqw2Y2A
PXHqIrZJm9HDMtusUOjPExaFrMZDTVLKKHJHBPhaw9R3MHQ72qwjHCLsLbvcjsQy2cxeeEBzRigB
5TkFE3SAXfbWR4if/m11v0YGM14QsL6FPn1cRSrY+VzRvnY4R/mVRCVLbNRVBWVDQQLfq6tqw6mw
42dELwkJbqJIeFW/DigBCcW0dEmuipo4XHSDR7plnTnx1wy3uJkQtj546D0XI9iSxBwwpF87j0yE
TjFIx60+vH0jWvJoVWNLec0sYX4yt17Vq/DfkXQb7ElUMwc9KHkdzYDftMuqIgYBaa94tZ12r8LX
RaJivmYhsQ+TAeXYBqwEE5bIt3cGms5bz+re3EQwMaJ1b6iy4kD1/0D645QWdppa1BoUp8H+rr7E
eHIOgEpulMJhN+AAB746C415MHqvFZrL/EtCjd0hLx8FENo02TMd5EBsS1osYtQ/R3+Uqoi3FH3L
8Xxsat9HVTw9Ah9XMb6FdUlCfHYbh85UbTnpIwBvFkGvZ7/9v+uCiOyltQ519Wf62VY8TateU1x/
e6l02aBArAKpOt+hKH/0INlj63ZI0+jvECH00CmBeaPARbEwDZzpq1WWaMwfpuKpsF/EBLipf+4U
rADDL/BLg6ZyXfP9oI8VRZAraTVjeHW4lCpbTO+s7RlkOIXonoWdpjke0Pa1fyNI3/EqmMLRal9p
3wgdN8n7CuldpQtTctEbq/yTUM5kuLaEWTvBAKdxXzy8PpjckzbUfgrUh2AJEgmirfKM952qINI0
AR4vDEb0BW4SsVHoF1G0RbAJ5YDwSa+vQsayRlXCEyj7lkccrPwYpFYwdsifReL3wscfR5JKQfCU
2KgoA4aZ+h43bvzu9pM6O8fkbC+u2OhXU5eYLPW9dR+eGAsbkibTyDXqYHxgZmXsaKnnRz17nwJN
p3NXiSzQoDs5qJVvqpEViVu/lbWShrmrb1xSjVHuxJ8rcvfxuP53AKGt+Xe4m3DbKC7XVh9GxIx5
UZbh1/ypI09xJjUdkpG75udtcIb4HchRkWV8WkTP0S4rqJ7iLUM+8ORB8voywqzgHdhAm5Rm0EdV
fqW6WBz5US6ESfIa+gOTE4/oZINvbIQ3wvwata7QKlTLnZ536weVXrixi4B3YFTuku7JcXG+LOGk
Z1YewLB/tzP52ILhoGrrXOymCQqM9eWA6LnioPQfnXk+tNwmiFlo0oCqZlmcUXLaG5UziPgsglyz
1ZmqbjUnL6l3UNCKX17s/ceOY39TRnL3h4qCr3cznwjVa0OsZ1CoxPjnUnLCxcS5ezP0vCx4qYk9
EayvvO4RP7JD5UdabjMSZVxEQX0ltRkcxC701WOiwarfEW3fZydJ4WElxlt40rlASBK2FdzCwkkz
ZnoHlauBeRcFV/+SH6g7y53DlLJ7xdTfKgq0nU5RtO5wcBHSdjJg2L6242bss2PDeIENs/M9nGJT
ZxPzUOS51e8WPMvbtMc9Ke1/T714zQ8UO9KbB5WjAUlYaUwk48Y7+j4PEVRYA6K7ZVgxlKY3TEyB
Qigp9UzsNcWenIG4xlknf1AzwvnQ73ShkI5PPl1MshO6HD2lAmiPkXTpMn+nXZsjsL4uX793+ndR
1UPUZnj7pt+aou1j1jpqk2Hu9jlc+T+4vuo6f9y8kGtp4kmMXJLDbuyvsjRPQ7bQk35xxG6JBk9/
uk4tOx5E9A027Qw8Ve19XIW9+bkMXHGpyCckhZzwXay7QruiBQK2DAlyOAZ335rpjfUMfVq90T6i
5wMCZfjNHOOCaXxCC6Kd+SQTI8tpuWaAcVaK1DJLBQY2/holppa0mcQ0S2zopcuFvfX9JTcvWqfY
hG7NnCqj7yAwYjHc+Xus54ciGPXNYkpbUVWXZnP3HU0vznogAO6EVEAKSiPzN8UUetT26MGGUr32
ysUI9zuAS2byWNunI3XFYl3XzZummwZXh0gXxqOEgel52ql/6cPr4ySX2hqd5WRZVRg+TZDVvCEZ
u5pTJjlDwXvb5tKC9j2Crtwe2RwbN2HIRpSMA+yJy32fgg3Si/b0ScHBWm+qXU6saxbgegKJqgkO
lzjPohd4v2ZhiLHWMZNH3RtcZP8SePP/LXUyp87VyN5fxH4Zh/8OADuUZQBniyDZYHCWaRxS/ROD
Qs49hnRRjyieh6e0oWOC2M5POt4w1C1P0hL58yMcmQum0+ARry5ykH5QVFFvATr8hBcggUfX8Evu
oeQkx92xChQkiMRkJBr1m1u7wBWOxcHJG896RCXDxmgvuoJ4ZvSGf0kj23bh2XrZzlsGvwF//RGC
Mg8Af7QCeQswNEG9ma0PZzeCQlMzo6MiokDdEPoyyE8m9Hj8zz6nlexbGoZJXoBuj5QIHSUL0YlL
8UwbzKRHTopAmYd7I7BYrmbNoMeI6GW/oTgvdLlZ7SZpToKnemF3tPUw9cOA4VYIaw2u+ZADptWd
RwqtuJZH21ke8uM7yppelpRMbk7sqUL2KemVAQITcfy/30q9SS1euGiwK37V9knrthCuZuYkQchA
HQ+pa1Fd+9qpdOHzwWCG1uHW5R7ZG29gDctsJOHSu4lZLkEdGfClcHnfYfNfaZgUSb5nxHdF+yTE
b+Y1PpFGVqTsTy4P68xz7s/aW7TZQRCRp3M5n7+HXDxCSsMb4SHOsSarZTLqKTTo88KRhz8uvQmn
1O8GHveMGFG9pU/QwSxMrVXwwv/c3n2Jxj5q1xOLW7g2EVIL7hW0wClAviYOHgXN1VgVRA58aNpS
rtmMKQwVlZZ5FkwBcM4jhyC8V4o196W3SmSW7UTZA8Z68xR6SPCipCpBcjjfcpC4HHP8d4x2aedS
lldSA7J2MFtkpbdXeFFIKikPoZsobM2YQBO5hqSum9BClXnPxhqVwYu4DpEoVp4q7AQ75sQRLD/d
CrIw71qtZiZMEussKn/aR4gqbuKU2FyvjwWVV35TafDPn4g+mk3SWUHfg/wNihoGRTsk3Nt7rFHY
NUps3eIqLiHzLq04ko31TcTh2w2H99nRMOQBn6FU+Ls969saI1cUevhSvAL2ksF50O2Kx4HEWYBE
+n3fnzsNrwtEX/QJP2O3/PkbrSdkSpb+vz+t2C/Y9tTaDyk11JKuOXZ22BQrAAm4h1ABJG3APGCx
L8qAyKZLOTDb+T26bKwFPbR+UkaBrXyWHnAB6caBdJOmJk/ZuTX+6xh9fTeN9EmoqFAaLIuwaJ75
cCD59yMLTS9NwbiPgkcHofcf+xmRPBEuHloMDBAI80RS1x4AW/7tvuNJY3aYllpBXhbis16egURs
Ppa2QSIbVQj6ZaawOn3ho0Mb7naIVYICcf2Tz8A/HP7B85TdbXjoZUBoKqi9nyy0gMpVuF1KqUjT
xRqt9FMDNoXmdF7cFK3PfW4gmKVgLZpHD2AuJmAx1bMsrRYdXqqv5slprtZoXMl5OTTUcOVjO0kF
/dhStp/NptCXAltO7QcwBxL4+RMR235t0MelCDJPXUpUMXQUTlSZSkoZi2oetPu97nsyUbMUblqy
fo5gqq2+LZLSjhXuT/54sCOMJkOwgdYFzqdra8yBB2s9sYsgecm4j7FsenZeNrNwYWFeORGJ7NTH
uEnjxw/wd3VLTVceM6RNqsAqigKyToDKfazm/iZqvNznOglGaDbrag1TfABfd5LNmd3s/Nb4L02h
7S4mUCNTbrCVBKak/zlspQ0I6TIKNlGxADyNbmG+FQDqYULTALtTl9fXHU7mNeubyGdsQcYZmDAs
CpmkFcjVa1c+b4SAasoASw4tUiRphVapPIlQ2hGQphvLUoGaQSVhyhiZsV2tN22MhD0lBGUx1R26
UxLsqT+qDHMPK2xexSeQbvc9apltLYcVfJZiXBaRlviORV/+z9QofP5LabQ0s67vqY7iVVr9RaOv
idQY8/Cy2zIXbcdrMu7htxe11JjowVY+2/120N30sMCpkJwSiLBqgHXWPcMGAxHq4FxNgLOVRRJp
51+/Yys4foH0Vumj5ZQJJyjU3cOpZeYKoQ3VQ1omL+9muc6rqhF4Re33I8adGR440DC6l9xlL+Yv
hN9gzBr1+aTLIG0LInktsdt1McC1qgHBoNu7Dnha2O7hdN/4gbpR4s+OBg/kmeczeBZccIeMHMNY
bZb1UQ13WKm4PIMA6Vcn2pv3B3L9462ma5ZMQHqcALLhUNpLMqhPot5zX/BNPsG8GUS5k//tbJjR
Fwa0bMhnaI4Rj6kmlLeJ7PcqaIzPkHU1u1bN+7iDup6jlI6NFjrH5uDnPj11Guor6DEkaQKI/KNP
+EWAyz/ZBxyXHY60nTJuAIgLZBjzdgQfmd35KgvEtkpBYyHWQahLwh87bk8S6A6jGCW7s3GpRz8W
3EfTvIMrkQFhxxzsw0lKNNvK8jj7QtStB2G+/1bmmJgYF4coi1KrG8Z5b1Mf4Wu17sz+1R6e1Ys7
RFhxm3Pomv60rhmYZfB5U+FLExtls8YX4z1I/eYSiRjShdP9ebhKJJYS7csprTKyDnQdGNz4u3ta
YJp3SaUS0aV3w3vJw2g5hKx0VMmvR7sdW9ERBdW/S9sUbhdqPOGh7z7NY5PIQa/dXq/EifyHVQvE
88k/rddi5/cbgm03vjKuc+xIvHEmhvqqa4BFh493+CljJlr23FzWz0+TaL+pzolxjYegvkaEbPd2
YhNLUGPwMnE9j5/J73PvB9OYw6u50LNHTt6Egs4aycK5UTblVEz5PxEiWXbzYNZaYDECi2rf0MRX
FoD17fxATdtceR5uUWbbxpw2O6QNzCScLlBvnkTLuTNVmjc4tJlBcdfgeyZzZ7fSToFJl7lVCTwe
f/ucV/TAOLRjbIHyV+TBOV0/5TWt3foRBq00Q8J++OhVYf1bpjMyBKz1Zl0L59L1L/1gd/14k209
flPx/O713ubGTP73AvFDy1Q0HDiMHw6/9m5S+83TPwvMCa4sJcX9U9LWEnBgMFhmvlBjG4UbqShN
WlOUOUmTVU2AIH+FINcv2eF6i+rx5czO9M2um6YN0ip+95Kz97N49LEqWd5gsDxP/FNPvaUOn6ep
iZLCzev65zEsiTGGivmAn86YsI6YI+TN7C4UaWI0rw99LqLg6C5+juL/+cG/46jtPvlbqt+3zxjg
Jw1mKWx8+JpYNGaNme7uaQxbBgnaarX8ZhLwshuhThZ+OILA1Xk1HSl50t5LwVTpkNqZ5ZDgPnRF
BVd1oZ4r7iYxBidi3pUYVP+Ox0VBUF3jjl+pXJqJzT04yrDL9DUOWBrczKgiq8XJ6GuAPPztP0Ji
hfZhfYhVKlDfsvvx4RYB87ahwtBjDJn5TUQPrtzdBb8c1LvDuDJlfzKqepbgQlQqGbKsY932Fqjn
qWPHwWUigp/sVCGTa67A4KBG1jjPvSk7GbI8wjRVjXTfTdTlsNMfXAQzyXH9pTPSV7rPbz/qPXG3
TG0fjThPUoa2cbgL68rLopr7PQjtlTI2rnWZ5Nh0CwfF1YpxLIgq/yigU+sRoTJCZ8ARyQITukND
YD8rR1T0WgERd1NdC8802YZztYDFkf1eyWGeRM7QV1utAoDhBGwNk1JJBiE5ZV/gq40EUjdY+NkA
Q97AQyEvXhdrzhZsMXUXOYc/45LYJ9a4tIvclC81FFNvc7jUnhQoXqNdhFOVwP8PDlBXNlmUtd0k
GlPQVXTBoO67RvUm3F5odgKIWB3wahGRZnnAh9eEm6ZSykVbZ9ua34VQ6XfLatQM90fUx6cxFOoB
VF6Hf0IrGjWTnYcSS4BbLY5mNyVwY8oQaB6ehlNEUp1IETrI14yWpxQ9PeGESQj8PGEuNcKoyquM
HWzmJW4RNkuTfXW0+qeB1UNlzdAtCLkN+jJqQdLAX/5l/dNfMW5M07kCyNolUi1IVzlH+4K2Ze7a
Y+14mryDQOSz2uM48BnfGHIrCRW8Y1IdACv+9wQUiUL8vIU3JNiiNjY6xzzM8XaqHIJqzcIxAbgf
F1f1KVnj5XINGqo3kD0Rdcuh05SvuM7YjbsiuhYIGcqr4iRg/aaxaEfYqdrgceNpqket9aaIksmt
QDe1A7H0t6XMtMpOurtl3SjgNUNKH5azNeIX6pbkC2dsIkzem80YFEC9rkMq9kH2Ib8u4AxXxR07
l7ERF/x4UZfBVPefJCr2h3Y7KPtFjHeV3i9THxnamYVAxZAhaDmUMVKCST/SxoXzSRryiIeEse+o
gJU4oiwstF57Avc3a5eu0Rs0AmIO3IWU0pUrZx79oAQfFtyWPYr0MzW56enYls8CbiOU4lmxHrN6
7eev5p99A11gbCRBw0nGpcsWCMJ6ytBn+OJ7scRNaVzOGOkiKnXGgljC8gl/fqiy9MSqL70k5NGD
BBrAXAQneX01n5f08TYc9hApLdtfKDWGYtdS1RgsK0nUl/JdXIXlYjMlup9Qk1SAtezvfRt5cXXY
9EQCjxlygV5iE0eDHhO8uvCRGKeRrA7SLXA/fhXX567D7nSsLLGTBSOfkNhg+d4kMM1S24azedKQ
4M+N7DQGdwB/Ll27V3Fq3fbLnUROvoRqd+u4Cqb7Vlswz/QPxpLiz6bvXly3QhEjYS6ncoT+3/xo
742yIFs1GctBNceqX1Vhh5CHsI0Qz/mN6mhNukC35fA9mPMKMR3LxIp5pvkvTIZffSXXOqLpmqKg
I1Uu8Icrvn2LPRTynXEIsGcHBv/rIGTD/dCcjpInK7I9BnBezBMH5cbKEYPJNphfWYvMTwq/mSu/
8Su+MZHw4HLxOrrP/IicQWvY9xNFgH3UbgSCE4gb361rAP7HQhMNfR9ntmteG2pI1kXgvGXZW1cu
vT90HMfGiJ/3Y/qJXwluwLBvdHeDGENw3iSkiqbKwgGPCOocNpt4EU9PCTMHwNF0rgsZPJmKPrdf
kZBu2eiq6UhyHpePPFlgBMbbTpMlFDS4pYtKn78NlzOh6BpMWi+SmTbeSQsHZ9OhMTWq00jc5SHb
+2BxYycEE5YmIIL9ro3Bdo4YHJ/m0AGQ/mZL053gYAnT5Z3xqSfGJzX1z5/Dz44WRaeZUJ2nqFU5
QKYuVUGVdIgENH1jFzud0H4QFd92wyaH6NKA/OAJF/6EMi3V+EawaKbdvvwueYEQ5yQtXbGKWbax
b77KeciiVjoRoe1JR2w5c4z5w9d1x3fz09nz6Iq7pm7sTEi/AddKBjRLBczdL2q0ndagSLjr3hwK
3S9HmuYoh2x213zb9bViiDmjrVCNvc+eS2odLsqSLmzof5KZl1nJFwLuD4xJJyqVRgCY+crGoicy
6eIq0ulf5rEO+FNQZXmz1rKufnJKzneel19Hlkf7z7ItR51Pv1YpNEp5e/GJ5a8Y8CzueEI1Tjjo
qi4Uw/Kpy0yFcel+zPSRnnMP25Nv2ucIyzO0urkINCU5WCZYq8WiNpnTY2D3jO8tisoToWI7QCPD
bzixZ0p6tVSOu3bR2xht9fcjK22qjhtOh3VGtEq0LCoSMxXFBcgD+uWk+FaD3CUbCNy0kW8Rb3qj
SakiOdUEC8IJhptNt5oz0zjIwDoJU+DgEM/hvzTQ7Oaf4YVd8zd03cfZNKHP9elOm/8VxMeDdRs+
K1kCKm8xGA4aagzyyLIaasU9M3089W6V5RYU+jXspxqaIX5yI/ZVVXnLK3ILTfhPpsU1bmWz0/kT
coBzCZ6KoWHsD4ZOB/wQjh9EA+m2JWd9fhRR/PGlV6ljGSwZnF68LRuiDVm2JIYMmkeRbLTpZbjI
Of5thSb46wwfnaV0cuEmw1rrdQYfGWY5g7YF9ODDbNp9dwYXwKPnkzlQErl0elDHS+NvY20soBaa
8mviNtDkx6/MJlhh5t14FkBkTv9Ak7Np/bCOmocwcHyMyRy6vmg/dlKVlTKxdaX3ScrBi86xFtqZ
95qJ4kh49YzyvwYq7nbvvbnynUDKBItWIjsa7X+z1vAULs3erF6UcJDRrEh+2ozYM3fe0gYakMEj
3tsCI10V8DQ+TXjfODBo5QCV3A2gkarsYQ6rMsZZGH/ukW26gePopIF9+fTB0Bzsgw5UOkC/dcLI
/VHpyDYyuK+RAdTAOMP3CO6a8dLCzJVyGWAyJKrcSaqEZZIo+NYDTet87NvMzuVZxDxvvF0suaMf
vYcUlaIXNOiVA0HDixXKUPbgh2jaehQNCIylxQ1J/rxkXPe6tmxA07Bc9tb+suLgIl0j3OQqI0t3
pa92XSzGAEP1W1C+4h55B6zWWtuBVjUQydyX9kr1g9UiFB5hixHuDHoQGJQxvGIbQLqkONxrso39
wAoEEszDyTS+tM1pVQFc1qEjv4TWfpA2X1P9pZdjAedNJ6eMJ7NEsUqZAZRx5d4FCpkOLZEAtgAO
6OUET/JNo3pTHRLlnns9DMG1BlFxRJDkNYUL7FDNSlt9JxBMuxBmFrWDixpOnNYhbpX5weDUDOVP
iHslcaabrWDF5VQMBj9eAaAV9GXA97NwOagNx2Xcb+UZCer0HFZfCPR+jyE9YrP4do1JApEqnNaV
z4IwNei4C9vC7CL3wZO+wmg6f33Nn8hACPfgzeMEkefe6b88ShMKbdBOziBvAfB6RA4ZAQtC0DqK
3Xs4SNi9XeIEMh+0CM95o0dRM2xFuBXUUkd8+Ks0nHCaDgeKywzJlceomFzTOLeRhbTCviCI7rIF
gFS7sjqukqqQweKZA+84VXEjS6WISBc/FOK8BkVV9IiQ02SbIZEVbcnNybp//Yci14DNZweEdrDV
W4jO9jUv2iaL5+klPEcZHWfxgmxpH9ciHHSQ8q6tZiq86FjQTQRmxAt9WUK/dA93iDGIY+cutR0z
Dt8pcojRWuGusWR+wfh7t7v2Z5W+CPsrf/jLf/xmwIbZyEmd9E09T9araP7u2SVQ6zdZyN2nMYJA
X+gqccTTY+psnnVxwcis9GKXpZVtrYx/bFVq/wSKyEyeSuG/41ReNk0I1Iq8tllTY5DsmwNDpYV4
1I2Y674hWDS7AGtXwOWKT3eiKJ48GJuK2ux8Cu1cNkyV/sbh2DqjoLRuzPQFOvw+jPwkgvIv3fIT
TONEF32+BDmpMdsP6hfJiyUFZxP3E08DlBfvcwvW4t8pYhLeaGL9D1XyPsFfoJPeY4GcYQLv6zOR
fP8qP9zU6Pq6F58bNnsoQMnuy4CykMDg3cPrwm+R7hy0lAo+6NfH/T5ff6chtet3LLkEYamAadvF
7ivPudxkXalg7LgTUzb4g1uM78iMgtA2qbk5rAahhUUz2cLPT/n9dkf4JogVeMq8ZPq7SGzzUoW0
pAGn3tJdThiSjV3bPyKM0no1FsM4UKByHHTJmfSJHYm9uXvsesgUGCYrkCBMiCcXvezXipKVqlDj
8dpp/2KtIok+tzIWL0vM0YBOln+H3UwVD8cPJrJ0xfOwa3PJ6PAr+S7m8tE9dFvyylRuFi2kWOaK
io80p2apw5Q284mQjqaUHeyWrEUUHQiFullYbOuy7u0d9qrr3S9HzYBeWatlyl31M7wzbSJADPnF
7gzFMKr4aFwsNvWPribOu3Or/hFbzXnjn92y9gPODMg4Gr5Zmsv3pbJ4CQfM5WVT1tO0jobLYcTj
cMcSaD+7D1Wh9WzYDhh7ceRRWtbRAfrgA60bKvSVrsvEwvIF25PI/pWUD9tLh4VCigTXgStYbQqY
1Wn05VRmu5nDfJe5OShetUPewavbHXZZ+Qj0pySxVJD+QxLWUPX8cIHqaIzAyNaAP16H1QR0AzCD
ZdyziTKPkQrgvOEq9i0G1+DMk9KAV4Az3OrsZvCm41WeTFekMc5rO2ZXBwpGZB2Y5MszlFPZ47Gc
pYgMkMeP7byhKyV8RhHuK12DY8DcbSEmuKexvWL4EE/MT7ibIM516VQXrk4LNogv/Z6QZ7ZWijsc
pho8OUi7lt8IvgRRGTdUzSMxRZtoSV+Syt+xZQwXaH0xgeJmx4eGrCYJJWqYI90cjpf2E9Pe9Vmf
YSN8GtU9a1I6TFsCKApNDEt8E2WPazm/q1mnqrItTTYms92qI5+bU5kiaiyZmOj1ZiLKUMgh8jp8
ut0w2fUwSO40wxoT8dtU8RIbdGXmQCfFHXekKvf4kTH2/abhhCYzjxlwMNFisVsJwAp3WRNFXLZD
nRYQ+3Bk6s+72uj6+2Vv65Z/EB431Biu3fvZoZdfAPjsl5QcbckAPMPhy188zajj0aITWTuLbw1d
TZ5ULUuoypOxmt2XChxByk7CtdOEOPbxogo9s6u4Bm6sjJxaxaeM7XKTTtejuczTssANQ/hmgLgP
CuzAFgbmsCRepm7XLAfPIHxe29IX29FISJzCfeZxm4FPkIC3fOpOKcGZMhsjG7gQIgNqwp6zcP3F
6EXYJL4trs2404tJDW9ZhDx+Cce0gOmEf8GBDw2K155eUi/OQmAYo9BtS8ckbda2kL9G0cvhaNCg
9+znt0+JcNXWwLWYdrDgHM3HHCne9U8fxtfH/RU5ZVfk+hjSvOZt9NILeNsQrQ+NrRJ63FHCvVXH
aJVNfoEK8lXrTAREXDBBismKjklHZlU8Wi19HB/Q+A8OcTlZPh4IKSFOUHEtqrTobQ9fGHfY+aUZ
Qp4Kg+IRg7OjBVrRyKbVEKT1O8s/SqgR7kOV0ZLhGPIOPbwmmORS2JPllibOLtbtQRRO6o7XLqY0
9nmbzf0VoXJlLE+YFAp+Z/4Ds7zJInQyeELScHtRitKQN0dyxw3oeL+/4EvI99FGtl4/Sm370qMv
65uVu+JCEYEkaYP2HT06x5E6AA2YrZZwMyRIFo9Mo3g1N0srMRt+9W134GYdsYgGQoiXU3TrFzxT
84tqyoUJFSEHyYaAXM+TiaYFaXieshv+BC1gXaOXyPAj2CsjbaKa+vYRV6hrnCmucylP46OGEQa+
LlIOZfG6gIm4aqC5CyR5a4T04viX6DZ81x4/PsxRqOLr3uaMjzeZpn63utEmQjkdYrwA0kIxWFT6
S1t6f3kFk+iuVzi28hNUXUoq7KUsuxiRhzP2JfE5qcaSeRPr+sXYlLLEuQU8+MEeJWJ8JZsc9r3A
zViVyaty9FQj2Cf7hgqTgpmKP2i+Veq46K8lhXgzHAWVR3K7VnvdVkEkIrvdVvueF7+IBG7HiMXO
kcGWhH9j0fABPpIBjFacIp49I1rRc/E/kGzUxeebD3tep/sfrsXkMUf0HgujIk0lNtAesNIzyi7O
xQvmbMubG7tqDtXIhUVt9gS5aT8w2YGqTqXyiRYudW6PE1zvXOzeoyM4o43CFMAlC0/C5mi+WbRe
d91idZEj+vrPeqiixazT/grGzDql901G2+TkUlSwZHsC3ibYOirTkwgkmZUkLbCaY6fmxYXZWwZl
J6CcWIifrX3fk7uou1lNJ6q42TTWjTX3fMV0detSBt3F1Qq4Vbw1ZlJr0uva05OMdAQtfL8z67ap
MBNOP6QLrXQq/w/vNzRfXH8YVHU00VJskxhYKS1OQZutJjiMcsPQf4VVjrZRVDERmHPpaLCsGmeI
hzPeEWCUU17O8vYYpaiB5NSSgjokxc/ggtBTEgJh2jGSI/yk1uvEeiHk5LJU1IQsFyLeH7S34H5H
ORcHdM/FXolxCJmj/RjGqvt0UZeU88mM6onYCKIyeX8RKwvlvtz29TZu1QyGx+OBV3m9MJY/FN45
rSWtyqXlvaYz10jMvc8oooAxZ922JZFD5GNIE2X328tXIX8V0/Xen92rzJU/N04U6kqF8nf2yTEe
125J+aqLhvgwK9Jz4+xbz4bjrOdJ/HsyoZHQOoM+GLA2TGuZPHW5J8dG+tlaGoj5234A45Jq/070
rKgYt1WQeAG4uw1OSUlvvV+B/6t5Urun7DzRgtmFJ7+vx+b8MSzwHI93PNLD9ULQ4vn2whmvDpsf
0OjTI02mR7eP4AkIPTUZuXDkQp91vbmCOh0U0BiP12k7qoFpeRqPvPwzijkYkIXAYX5k0pK2onQH
dTBLbjidxIeV4aHbjZiNeWnFhzq8QZBp10CmPYLXzY4UDLOZcPit5jEfzAmApc7bvLbozUKfXexQ
58Ksu+Mjdby9W9v+4tVXbwHx3stEoApIkBtG45+MGyy/iDuAt95I1eBmlMMI7+UkWUjtkKHLUDdM
2qh6cLNrTgsUJIoMEsaamYpg3M68Q8rGIoxzf64riGDkm2fOjejekhZJXt/ujYFzmKTfOo+wSoUj
F/BYiJF6ODAuUqCXIG+Hkdf1Dtq5gTZUQwXyMqaOPkOM04lj41KsZTEzS0Bzl73s8WNbbyQe4+VL
srAtgtXnpPXfWxR5DClk7xSP8/ZF50QlPDC5sXj504les7I25CD5Yc8oCrtCLmf/ELxzfE2jH1yI
tEjdfCbceZmE8kRzI9bLdfpkXpgrqUs+VEzC3uwxStDlLCcsPNREEVVuy+3kIXdO+tcBBRVuB0xI
+v3M3HLl121VIydl2juhVc/JFkeqF8PG6sQnF6/6g6DvdIziPJgx4nIhLJNfz9KAHnc5m/m0GraC
Hv+cUfT9RLSTZ+IN360ZiDvOHQ8/Ijbsv5kWbazROwG2e67fErwdUecsgDRzvNA9AxQZFoPfUZAl
snGhPpNGoACYIRh35YKXBaZfmpCBRUJ5rQ/4nF1jFsNXJ5wnZjz6EeqiUfwtmnPwV0Jnw/PpgIgw
2fo7CxY1rQZcb6AuQ62PTPmRQmPeWsXrudvKwdJk2gJfkwLNGbZrPKUiPoLzI9qgjBKxVbO13aAM
ht0DmnRr/AjpSyKmeCX9ypF7Ywz+K6OmmeIJvTvzvkIXLSc3yatnQuj2+Rl03HnSOnYN+1cTn4Nq
r7/d3XJPv8aHJQqg+7lmLjqy6/c5BMwds70NV7PaIDrR5Y2bh3arN3v0nEhAMNKtNWe4atydEANw
7Z8It5ZhexFH0SR4c1HpHSjS0bM4g3G+qKZU2qySdyvdnn3GWnYI0ulBblnin9Ceoep7Gn4VpmAl
VZ9H+/pvDz5SMzA9iHm3qvVeXyPJpdj2zQhl5jIyUyNvkYTdvNuoZi2pzN6QbdwrTfEStm0xeFrT
3PQa43sSKoXP5YtuKZ78ffNumNkp6TWPQz7enDl3noT8z0c9lgJdaCIw7D7Mo2xLIpPh6atPnue8
WSjR769NH3e9M1h+Cz8kymaEFSzODUPIsgCFFLqx63dY1EY+59gV11jATng+GB9hFbIr4+WI+Jft
dJ0iPDs7H2Zy+0i+yGfkxSfAbm7/t67tvvgN3YKDde7oSKPq8kWIhrGuP1fKqdbG+uOXVaSO9Oqd
9/WBxKnrhJIUFQxRWX7BsIITzearwT7af/jE6x13DjsjOEt0b/1HQiyIS7FS8r6Mc4D8je0+bIhk
5WA5rFEhFh6wQdSfpgXSJi7SG6Our63Z9uVNxKfZHby3yyaXihMctF/zNpIAdx0rvhFuAHA2S+NS
9Z+AaBQEBH49SqutOET9tn8MvPrSNGNeBN37e6pb6sWpxDP0tDRddxm6tOsIR4c2obPleA/mBtZR
zWyyNqyJfixU3fuOo8FqPNI822DZbZbpDgZTvgxR4YJR8ISxwhVCwOTUlkfqVg1ey3ChnRCOHWeI
MnTBvgt06MuF8ViogP9pDYwV1SUx/NoAFRJs7PrbKNb56m1Yft0QHTG59Y2tjkqdPU4msaoCK7Fp
k+LpnPtz4jDAf5pl9MJKsJcLNSkX06MNtW2C33gSTxOrpXMYgoqK9wBskfBya7hSRDWLdJpFy52j
PpkyVlVPqEi3BrFrwMm5Xnu1AGJAyivgAsu+NRejo3lfOPA3wMt/Egx9jf+iPGtgyxfiTeRv/dPm
LidlKJu6zRuXy1Oy2GjI9ZE+AqOTUAqQstNYvW6R8MR/XVbYG/4ZMGXyumBLZlaPNqYVGdK7VP5U
lOTnLwHTxJT5VTApla3I5N7+FevWRp+H4odzZ/pYPxn6Y6UxpEKzcUVXxk2rLT1X0BfZ0FXUzfse
t1X1zGmt4NX8vV/pvTmkGlmBIOq+f/WJo35IrkQJVq2iNtJNQArpttBvE/H8Y1xJ70dka2f+SfkJ
L7Z10HcuHfY7XKmJV/27R2CDuy1Pi3OKZIUCnzCBrypdoLkXfLodAmBTpbg7u8LC6/w13O5mjMu+
nEmMzoWtfXjgEIDeNg5CnnZGNq0uM0k0JxnJdZ8DpbkEd5zlgNljxp+xQ6wUBlSoVQdPBGcIZB5c
PO6qb4bkPG2H9ACIXXMZDvlVlO1KlBI12R/0fnpsq5xMJV9foQVuMqBNCQv/Lxi4oYAQs33TcvDl
CtxzNALCpUCKd2A5dfXZ3gNmz5XN4LanlD3xGqoFti/neGu2GwONTfYB4JBQDb59PyZDGZ77E1Hd
0eK07m7gpPc8qCsCVYlwj/UWpZsENhGxIew5Kp5qupm4vEawo/1+kj8GysDz+LaHM2/h+dWIRFOr
NUPWvp8vxM+53WvevQgE5atdSGALXVVF+AroWihT6cDR1fMjctp+T3v+zszZUpU9Jpw5O9Y3deLV
2N73pp0kFBHrx5F8GdSIWqXOVxOE4jdM5MKhaAWXGjn5N2OvOHLVYyIolVfLPAqOyCD57OZR28P/
ewusmrQTkl53PQvBIBhcl4IqpZYvNCVXnoo8pVQ9F8QCnGN6OHlav+8Z8ERDrt3vo3yp1Q+0S1RA
F+ciZaSi21ZWiArGsJh4T1dal/9DIp1LcaIgWtvtIsIHshghibMk8wH9a55BO2AW6QEQAO6gaytt
xt4HusiU7W0Y4bpG2S3pbFSu2HCbGcAnzDgw+BLbymsxQXHaMCWU3iOpg2NBWpv1bmYbf6H4NeRl
1iY6acV+bbQvxO6vXS+cH4HIpfDRNiTHIHsS9XAVfg6QZk6Tg+HGcIZqWqOBC+8XVUKvQypWZFTc
mfFjoAFUBuCuNjT6eXVrdhGmGxw1lSsZveo4xLnUS/mfByUwufumlPqzZbNaVEts0zYiWvY68xPR
2QYWJOZop6U95G+m20Lt1Fid1j/6sUJdLvhLOLfSuF7Ozi1kUbKMuttqUqHWIt82C41W3LEFtMUz
KTX1OjElKLVv/fNQVGIwrP01vd6gBrtfa1ivuIzGF1Z730A1Yx4sMkwv6bArEB50QVzjbB8FxOm0
xertSiOl8WBF30q5yb/8EQqpd05FDEp/h6/AEvUeocZTnulgNxeQHFFBHEF2ktFNbyhP+oSycLqN
EzqKGBa1GUtDo/RALMC3haMPNl6pDUqgOsDs8M0E74px6R39Jh77yjtv3rvjTDK1hVjxh+1yvein
R65o32dxQnPAkyhBFczkudCWLTPAl+TZB3VTDPg+z1lVaRWKhpM8eM3rTEpl8xmmyWg9EDe3rOos
W3LXyDdewkmN5O/Q4Ct0aDxhqTOlLOwO1AUmWnHb/WTr+In/T6CI2tnX+HBa/9fcisHxtNsv+s0/
zVSzeYuMvKAsSnGD9n4ZnKH01NTX8gX/hXXr9hhhVPd2rVT0QefGi04vDNAPz+10JLDCurGuY3n6
L6dwibezRxJIHdR7I8wDC2rIcuwxio9D1r42LlaMR/+jRRY2k0wzcmQPHs69hmz3SEnHiPLVLSWb
1ocZIYET+xXzFNsVGXU4AqrWsl/YrJDZ78D0SgNomL+08vLg4nK3+IIuxF7baMg+M85wGqH+C9b+
511cmW4Z2/IPUdGxmUJmu057YJ/CsmYWBEs/wXYtsCG1lRaW0ggwa9nrAUumIFkRKh5ZRrIl/yUv
CIM8RYiiZ4GpyHdWT1M+3yDXb/7dGKQNIHUlvFn/Rxb2dl4ks82ifXjo3bP4Pn7YuOo2eGCSd4kP
RYrZruNSJ/LEBthMwb6a4VR/U+Pdv5IxHLt6gpFkoncbg6WC06uemvr7LtodVmTWC2tErGFjrgaB
u+IV1IqSsN+TLH75P6YsSt/ge9OdfQmw/k68CoE0uo+/rN8n3jjPq8r3eT6vhpSaHZ+Sxidw1YPq
8oMa3wzWCx9tk5Uje4LyB89/ay/grAxO7aIn6Hlawr8l2pnLhWVKPS6sWx5gT/JoP6MDwAQIH9nV
wHxj31mKmH8mYJCA/UhCU2uMj/UuT5MaZosA1+zZ79SNcJnWsaRTGYnA6bvCGe1eKRY/jGWeoFr5
e3I0Mp2pWFoxGb+Enpf4BnXL3Y/MuJ7tAbEh8E3XQWUctcAAMuMSK/osyI5P7RLlZmTpyero2o+V
2pJr2zrhV6UCxUGiJin0uqqlvdxsXZGxVzadfE+GygLAEYlzriYehY1dCEXT6exg/AifFA4TTqBp
eQ9yfQbSvcBsh1UyOt81M9rLQWYTFvR2GLAmgdkFaHIz0jvTDa7U2WTaERzJ06OT0nM/0nGlCUJZ
+iknK/64GGTGzll405wj2VXRRTrYp7j6FinPtDuZpkM3aTLsXK5t3neT//hQ1OHPDq/csgTVSynM
n0Pjt2n50QJd6v8ucbSwPIcVR9iUasDF5OVCCsg7wn3ENKTnVJtoRm9TMPFT/jHqQCWIP935n+Ml
F1YQH7V8eGyNqOt+1QHNgRDuyo8rXx40yZBBj1KpLQnNzNeWV3u9wDewkEvu7Kce0bSMo025YOeG
x8sGIC8T1nfJh9qbjjqsFbZ2tUXs5PuuYDX1LiXhV7BcqNK/rnSQv/QgqgESu4FaLi2LRbbjJjq4
38tQOjnxFEHX35L0ogpT64Feen8Cbk4BvnLq0xa7Y1NPv/MBQgp5mxTKc26cbVKmIxWoPaVsNeZI
8v+Ow/T5CAyy5i5f2Qnu35KS4q5J0QPb0S1kSEuYvW1TikucoBrdp21b5cPlsnwaT5rdMDSg/LWI
BbyP5aPlnOW78eXENWKmmGNTD6o5Qgur2rUv+kQsOuEP+CQdRvS8dhFr4kVp1bdyOyaO6y/xmA2U
9kl5PJxK7wSHHikDLPExShw5dnlG7Bt8Am035GVwJBCVvqMRpumKU4VVKXf2tBMvJAu8b+kjGAPO
BnHXd1MdJf5lk0udqblJk12GTEeVzY7dElCkx60Ur77ldgJs19jIpOPOXey/knaz13hejuex4NjE
44Lq9TZp8yHf/LcmmZgpQtBKZCM2bfrk88WOBERIHAU3+8iQX1CS9X3gN6DSY3QfVSc8kPrg8E9c
5+ChAGK1befrom13Q6/kPZcGa7up42BmTmDOYH9UStikGmnLocsW4l3/XigZLHCcJyuax/isBenH
oq5deb9tkVB83Qiyrhz3VunoBPzoQwBjFbgZvhrDpBm6o/LFsnMwEI0XHTB+FFMvRobuqJ5HWOLs
QcC9pIoZTIhhxk50hlEVWW/QD1XZnc6IYqcMTOG+1FQGOXmsTKfW4w/i6PGM11n6/2a/gDdH54eW
XCD/kb0lAT+/OID9QpY7Jyv6fnBZNYX0C4Q2dDWrMZaj8dD84zTO9pfzneOmVV3JuURf7I9ikEyA
oQABtI9/72znayNdZ41t992afD0W1kF7v4HER/I+H8N9Ncc/GD2ZWyTSeTelv0SK9nK+c2EL6N97
Tuqz83/HkYNILaUcHW0hwFlwDLdPvT4HiJfI8RCvEsRD4GLm6N+G1fvBvdmkvdzDUN5UZLIaXytR
joLXhzzDquE0YFpf2FtUjd32ecs68/QEwBXQkdgEo8Nolttf5rLcfqXuzRbgv2wd4vsGljJBMNrO
pcK1b2wSiDbDNEQbEGVftRZ2tm6sOkP3tWDc3LL4b0Jh4pX/qQMwhj1LUZal3ggQGKFoFTGx6e4b
020FAUZptTykvg/g+w1D8CBYoOUD6UlP0mAwZpM5yWDTtejFi/1qnYPgVErN7tQ2IZBT55R4ocqw
T2SS0tig69fvWmlObfLWLte49khplqGLr4Et0UR+b/0knzSABPnFB/vwWljSiz+Gvix6aD7SETWo
mupMXTBex9kMGvPHpbY5E/kY444RfJzm77iNhpX/yJCX4sl6lSX1suknG8hEVKOY0nnW64oBtcub
LNuciOfglDUzxo4SGMpH+gsVPwBULYf+Qyzt9dAoFekYMSGC7otn8MRAMBiEixT0dlukONsV55+3
AzfVAnvyQUdlcTrMwapCCoa8WhfljpcgEFCIEJlOFszfx2jU8jyhusYfgnm1c1QJjUYIvKGzg2P6
wUhgEbfV8ZRJRqnN+tPBtqJ6VLwKDGDh2j5q+GJQeXPKBWZMfEt5tRLBtD4qIVxCzBXyN6Pg26kw
2oaeaE6KBTUxk7GV/sucNCTdVxqzLEP5GAgH8puvMFPLjUVvmGYRPKFJQVIg7Yjzhz0oJtqJ11dQ
w5rAN+ddan+cTYkkme/Jk/d3uA1EnQnbNVz+1z9i1KsHHsvy11xSiVI5srzPU9WPA4tCw9hdXr0V
NoCyIHlMywzQDh4xZDwlvkDDfJs18mRdOLrd8iw8sLi0VdUbFYZJVqKHzL9InkNCTcn3EmIke8oq
vTYzoY7QdShNAN9HXHl2w7pI3SquHZCRISlCXbpMhH6t83DVsXCuBbX7VdbfpzxpgISoely3DquA
cMO12VWs+mCjN10jFSUcXkBgwA4dGnDzQCpoEsTeQlMkuuVWplwfx1O0fM0ihPHRPokxhvVZaJxp
IH7Sf9/Q4bbJD8heghHc99ztu8wFH1NiVS+bzXH2/U60/5bBGx6glHQuYW1V7uK080ySBd66SDmH
xiZAgvOcxKQq0SAoqk/VqdDo07Xs0SeHccwOiXTgKrA/eInjAtOxae8n4iEszIN0jx8PvLmIqtbP
iR6NaRse8qXKcNeWXNSJIiHp65z19sChk601InlvbrxC/lkFMWVHkb6N7kaylI6yrGMrNCFPOb/7
Z1J4IVHjlgsfSnUh9e8x3ua/FOEQ+U9b5J2CaXRX97w8lR0xM+pzLj4peEJw/N/wRHqC+YDynWBu
Z0SEUobe1BjLb7kkbNUuGM0FOW+JrrX6nHUyryNGz0k31viQ2KNwfr/gsQiWV4w+HfErVwOkcuQO
0+ZrmH6VqhjzR+Xh0+cIcCWPTURGXfn1DZZbxfKytjb4iMg+ruGROMc1uN40UpJ5czHkAcRMJTey
hbWqLrNpURDoRXhwrt6ibn2X2YnCPtgyud7gTzdqls8y48H8kealSU9xONDLRzx5BfrleMphRpoY
KBHftVwDg0U+9cqy5K0fyY+z5BQ0hnfZ2iE86rKgJmvykaECzTGS3P2JnK2DZxeoXvcZgEsbMDOK
TrZitH7jZhaCKSAKauJ1QK1V0MDEhLlsS4Lwfl/NXtFq78PIhQG76GDp5Fyf/IHqLytcSd0+uUEO
uSraNore2dlSWEGMsDs9FeQBqxuQvxsTnvaNS2Sk6mMvCIPPwxrYqN/o28P4nAv4eyypQ/aPzFPq
RLF6Y0M5FSWsWkHnCYTs0AGfcolhlY3VeQT2QnuwzATP2d/fOLVz3ndfdxxoiM5D1VGaHZH6VJPX
HwOw7XhnMUgofbz/jqUjBAYCQSRMLr6fEKa6v8akMGIA6YfJDsP6AeyVQtr36OZJv2l4Gv4RxTA5
a8y7MOOQtq3S1ab8wy/xfijAb6MUKXqXzY3f5WcNEmRbajnlb1LTmrP0i6KNlBtWD+vAPzTPJNxT
0NvthgKB182rqQGBBmLlKrRUsnjGRzw/9hU6a+OOIZCsVVWPj6EXNTJplaQlDWIh03AuQ1WKrcPA
nfJAq61ArZAKX+u25tZUqdZ3HrI9E1ec02G2UgYH5wHVEST/OEo3FbnJCdy7U3HprbX6idsDYmca
UPY1K8mQiUCm2HiLCe6TY8YVYkOBWg6/qgs1uTc6YTw/Yxy02p6MJmydZCmSpJ8yU883+zwFb8Gk
TUU2nPrfFQ9Tlz1ftalZLMhB0bDM9uuRF97zaSJethnPCL8Tz0QvqOI21IhfozmCzo4g93gJfvHD
CrEgIe4ocu8Rvjzt2VrDtwRndI1oynxtZ/7AVzMaiSREPPbi6qLXgBfv/GDtP7UlAi/Rk0b6Khxd
HLiI1Fis0F/tugxqqmzxYBNOpfQDgyHEMskdCKnFp+W77beyl5BwGgvzE4bY18oyaSPiFBVAfc4S
MHT59OZOxOX3r3Tbc7kjUQD8a54qZaVr+KaYRHOeT8uqTz8pNlJ2yqYej7r1xzOQjAa0qt2N19NO
Nj5M4O/qeF5uJ1Q8RmEXXMw9/ooTVC2Yu8l47HeYppdaRXqskaSvu2uuxAs8iXHPqcMwpzm3qH7d
6G7h7GAZCgnZl3gmHj3N0vDAyjPfL6JQneTy8lDJH2BdTaCMEB44z54bB/6VqDjMp4gTViQI4a04
1x443XMXIczRdwdbsrC3MuBysk5ECj3KcmGkcmwnkbXO1s/i7k+J+DtT+zTUFfBxTSxu8prNe0Kw
1wlVMAOn0yznlRIFdh/MnMTDfDrgXzw7dqEJAPJCPdMO2wc9bRylFPHbFR77HkSNDXPyyNJume/X
ZDwygUR0YHBZZjXyc3d0miHnjp3VA1nZKornBh0f/qz1eLmF1B2X8gkx1wAXN7TbblCaZay1yOt1
CMouci+xKkIVGgy1G4jcXgoktsPHyga8V9E+HLy+Q5gwI7jdOG0laS3QtYb/zyRXx0zlNYbed4c8
jwke7Ho7hxhv9gvg9YsYGJA6f6JkrR4j9N0sseV2y2mJyN4Cb7xAbbLcMRX/CYCox40GXmsO7heY
AzRgd1dkgmUqafnQ8AaHAdd8siAb2VfWG98rpQVGBf2XT34MK1cT+j8vr4ReLzoTc13Zmg+wAxZb
ELQJpU1c32dKy46/hNNK/nz/rtF/okW8SyDKMe4FLN6wTYHmrpoQg78f1zCMYUk4s3OCfyf7bbOL
AEH/beJUj0QjpIz2Oo/gL50Xr5h3p1kpvBqQyVEJzESlZv3Hnc0QNMwd3PnGpFb2BWIrFuRJpMvM
57luyIS6CfFKO/5uTNVdpNww7+sNRcJS97nySvknvj2pAsdc8JlJCiA4Vj9CTl1362T0gLgXOhDa
/9gcvL1oOwo+/0aqEaE2Pk94H2fkX8G3dk0/DhtmrcLZzBrkV20mfPeKwVEAJoWbT+Tl4qK2rNpC
kmvdUZnXy2BWK5YEwkxJDqu9p9xLGz4NDf/XjjKWaij+Mw6brcdg9fffGV/hu6tE22YfOkDd6FDa
gL0jmeHC4X1Al2uEy17Yl9qCYPV57nnUzGXGBMQFoXKjvtfAOQQR9tBoxGopKGtcUoyTPAnx//Vj
pEx5C4Qrsy4uzpmigqtGtZAGZZqSzglEwHaOU4v2sfpaAIeCdHJgxR7BLAZ/EJSuN2k9Tk8y1Qc1
xZftPrDLCD1Fb1n5MOD38vMLhacTEGWN+EbyvRCqHZT97qTLMf1O0LsZrP34LQUthepr/kyueCCT
i6KaYBjHybZzG8lCWIA94uqwx26Ni/CcLXaVrSDYacEtTxGG25lN/ijWbsMlKebmQSjKpnEj2RGF
2sboPS2TA/RC+R27LaBfZSJKi7pQNdthCFoNIwykr2A1cz0pfkPNyXK6pvCjqw35csefgDV2jw3m
rzJQSFEPGE1HB2HJAaPwOGz8J81ZAs0LJILXoQCTU0mZ6EZzZa715MJZMElsoxDkF023TPoD9No+
El9/JNyy7SNIT8n0asyCgSqVlVu2zKjtqFyNutxZtAm8gkik5z++7A/t2yvX4G7QoBHQtj0w+LBy
+HX5TgwM5253kN2fDk+ZtKY24BmmvB++W625wH5i5YzRj2ok2SpaRa6pJZkoBJUn6u32ajHALkrq
1OWmEuerMdWNzCX+BjJ4FyZFp6bRY9HHTj6UrDYz7H55gzeesfN0fFqReSq3VHpbfRQQCzaaEw+/
rvcy971x35lU/fetxKYccuzVZckU4grue6xnBxP144Bc34IWFlZt+dvOWoK6RrF+dXC8WNt/0cZ6
RIES8xbkK7QVqr15cLVfc7n9HWRrZauIYz5l9DMHpntngnFtFRr1pOtz9ivMiOQApPyQmA5DLRa1
fTEdUJxYfGlb6KAcu6+KsgeUi0rJMKl72JD0nLckjMnUhaUj7Jtbz33ng9Qh99iRhf9DKv5I0l35
6bpEpuAMUEfxktuUJsjBzjAm5ukaAjP5syZdWXKm3pbWx2aHy0etpEme2j5VOLEvLrY6Hd8JxHed
/GgjI2QuOOFLz295enVGGGO6ywbKsrkP40dl2xdxEyvAKQ8qflbHUxWhZfvoQhJGrNQgxJid9BZG
W1CSRaC3yQQR/HuoqEJn4VCMXNdF+bQscN4qmE55Or9yG8kKq1Rrv4ZIPX19JS/Een1LNfzNZ+YJ
kdSWUcrcAEvyUbNdjJQeoujdDidvZVkUAK1nBspMDukpMgD/E/GGr0+7oMqwDV0TjXBRX8P7pTx3
hmCAjt7+aI5tlneEs3UCGxDD/TkrsR1uIo3iMVb2UE2DixQG/sJh9Fn7svyBHEuSco1Ew8idg6w0
4ThpZcUw/M8WM3Rzh7o4Zh3L26r5MKdkWiaQ+Ilt8gcChf8ahZr89AZ7SCOMayp8JdDA3GmwkWt6
rsVMhgHg504PM3zpfQoaEBV3uXLIb6n17qu2gfq4dD9QzcL+pDJNu1iR9sb7yiRvb89sU6ltCjDS
2FHoJnQBl+DZAxEcrI/4pDON+g0rC0QnzFozer1xUY1s4qKGczOZ4/mTJ/MrJ19G0VlCpf51pCGx
cCyP6+ooo7ZcCn6MpmwEuJ9ilcpGfswUSV2n/rcZzX8+2RWvvgZkzU1ICn5jqvCOCFDmuhC/Q7sC
+b4BmncmYfnGlj8SJgc8v+1QaT/6wqbGavkpL12EwenPaJXRnFg0ToV4gec4uJ7J6RDS8PJDrm+B
9t1Ow1DTQb8U9XaT3g2+vQEpjp8mHLzW0wpko05Tz5ACNqTC7nywIGuUS/8cgTPUcWlUwo7iz6C1
rVBzEyci6c7CZYdK/a0j/ntXpa1ieepSwuymUyAb0dnlziI5RsP6Pu41vnc2Dpx+rKLa9PoNU41p
s3TrvLW1Abi4k5YL4ps7E3aGFfHZD5q4GrmQCT5pXAeBJ32EXOuF9zBJ9ijvqaQPZUZXycdKsaof
8mq2RBBtn+7eaXqzM3Hzb3urN17sWkWSedM9LSHxsqq4zCffJd9ao0XOmsZENBOhra6loWQxanaG
PstSFF6QchW8MSnwNCSZZ0EHBKW1S6sdDleqxLd7Itq93lL8+g26teY1hwGTA9ISZqTUeuYSbrLO
qJnUuD9ccyWlkgLYZ1J/8VwhuyMK+5fs3Sg5nxYhlpzAYv3FHfKwxSCNuRh4eJPwjAeQ1LsGFPXe
9pfnUPRHeNkxMzkL/3hNS6/LhXg5X+PnVwDRsSocOUUvzbrMvWFOJ5ejYJNFyrY8ZpxBS/3UwEBU
2PuuWmMzz5pgT/RtlwCtoXvx4p9yUkx7d3IdHmV6jxK3fv/rRiJSJnp0l4lnKE0OgtqGwuSuPa6m
RSrM1xneZAiNdCZ7AvndaxA6QlDc2yVBY6ptXtcx+jMIIfCX1P8zZh2qTFvx0zNAuQaHNtjZDK6W
ni5MulR+uwAC8srRLOr/EUgrlnWN2sWm8oJqX7jqjVg4NASY59e+XKRU+jAQQchfZ8CJDBFrNfmh
nXTGaQLfqg1AK/pqMO9X3M8HQEoN+wTLAUV670lJMma/6wwlYf/f7ECVm53mB19cO3FMTYp86E9o
jXSuRkYUv7+Yyr069Yco8o467QqiaZaidnJW2KZDs8xURLNVwrfAZ57AnF14Phf2jltFNiSZeyR3
2kE1smbB88/z/1+Axg2mTUq4rhwzK4bZ2oQz38g9OpCjqPvqDzYL7am8EknqyB2F660VFMjX815O
0qv9r9HvSYJCVfswu3Dm3sSZpgzOfq5w2iWXf/PmOHiLNRs+a0glG7oe3ef9I7vClyDGotJpTqQE
I1F6GyW1wJc3BFbL6EiegVsMfmLqp456NVEl/JqEqI/JbELlWVUrvpE1lacVcoR0S7GEvBr5Qims
0rDWsZwvk6oKFZSPTzmQ9hIB+YNBeng4qigV+Ssj2qGK15Iz3oPSLejjY/3NByJJkLepw+JXsN9K
GHOeB8Cuzqe36NA5sqbCDC6vAfSpEW+grm/xrMbHqxjVBtAV79zEE3Qy6sxrhEG3A7FnKCkmM5Gi
icgYZR4lUeTmmxJVgYVcEIK0mMDSBzlwi1etywqkuGLFSaOqQJVLMfFOI0BVqqLVVDTW4k5Y3xm6
iIA8ZTHM3kOU8qXkfrzxzqTRaU7D79TF66hnhr7C6dAN1WtW3Fud1I8YXOzZI8R8sIZw9vN4lnyB
nY2QtAUX5uRqWiSvUPcZ/NZCp4hj1/u77z4u+KFCtQ88S18vp/gIkTHnwG2kmuSAQPraEunPr7ey
HnsZ1x/FTLuNLWJFOaEFjXtx/yjyOoaDZ+HmUxOcculYQAsk8jNm4v4VJyviYy+ilx+5g2qOzYke
lAgb44UjnYx8bsk8ahRt7TR4Rwfa7/7Qlt0bZmyFVWYW2lacfIaP2rSSCoLYEOqWV6cbej+KtKk1
I/TdoQ+KreAhZt5F7qkUxJjOM7miA6lizQkDbKqM9Mxj7O+V3PrKZBxtSHx9Yw0QRC1IFrlT4VH+
/Nze5OO+Romz93U0n/4h4mky/2DtthKjTwtBqZ7qpD+ZVfBx1OZCxc4Tm9PO3MklhmVbe4nSpmEW
vxdlytE0/WK2W9DO5CQ/egOKikdbXoiU9qIHLfGeWWgaj7KzxDsHFjU9K5NW6C8bFE3AMqnmqSeA
6dwyS+HWJMuBOe0bx/Z2M4Pua3ZTTKIgNXc5KK5tU0I7PcbYCW4wmRC/unsi5xAUAfmw7ZXhaREC
FJgfyP2JZvhJpRH95/eynxYDb0N9vYV8vCE7AlkglOqv1QtwMa77z7ylGZDIFHrQt/prQmA8mxtX
5bVtCTsLEuJPmwKymFly+TlVPXYMhbXDhFV65bREI46br0IORMNgnLYXB7IDMrUv0XjgX1Sz7pYu
FSJmif55yzVl9J5WL7mj/qkz9k9rI2WUniyP1WcxfwhXPBn1BSy1wlKfUpbOswWjCvThfn6XzELC
43jEqsQeAncju2EC9MfE/fxwdObtVE/fQHYSxKTENT9+NCc1iO9sXRLT03AL/E2NIr4LReWuL0ub
Qh5FXGFt88zh9rdVUJ0lznzkWPMkumoBUxfpHTbgXTDhAYQoEPGg7VsHtbZiBrqPiK71Kqo/WTL3
/Htdbvjey96MIzOBtYn5OfXGPldi3p/xW75xutDzd0LIQeGO5qFdLzPs7YN2Hvi+jc0TLEqmoeQl
5WVOjCnyqgr8HOG5JpfvbGwVe/kMSYzBtcMU4ZySDKvtEO5ZmLsFF3//mdN3fwx9YdVSQ3HRGJRA
THb9/5ojUxw5CmOymolWfiH8KMrgiXBqUzXy5qA/2PGdbl00yJ4cL/pVuxukyJJWKRKdaHuRk+R8
vA7KYAl6VU6eK8Onvs1gNzUDmPreD/8tXvSZIgm9twToDSqB7j+rV7kLJnzpSv4Kr+L0DUbyYJfJ
f30ilrlfnC5Eb4ymVScP/F6NlWaU3sC0Qt2nn0aCbMqidVzPWEfI7Znz6+80Iv+TnyVOxDXRpnj/
N9Nlska621htDlJSubHbrRPn/YjsIQmPOoXYBfHZW1coG4BCFOQjBzOksnwFG0O0DS0IwG2GukgD
KASKYE66wtqiz8710DiUUemj5+BY9uiCesqeS5hQnXUW1nn+9owB2zWCncqF/S6xI0hBf+DCoHqV
qAKKxTN2hHTELfUnoXWI3VflnJHGilHTrfIw2mb9rIIvAye11/j7ovhRyzSIiLjmyDUi2Ckzr07m
W6ODTfPV7Otc/SXS7sSR/PuYjDxe9pwAsmRekeku4FE66Pm7USPwlI/yjy6ZAk55Q6y//DabWdbv
O76A27SM0wI87lzHOLAw5tWYPDoR6LM0gtBef3tpjqUZB+gG3wf6Oacs3JdE1OXFELGl6Oxo+rTH
fp7bJf6NIfYw4tY6mtjruX4CwedoJqUX5cXqNIdf2jeJlEm+AqPw70RS0qYcRXY1A7JweDALkAaE
nO9sFgAQ5n/7Gfm/+QT9vNN4/A64vmrGIQqoL2/FyY5NE41veGmmwN+eblP5YyVDsNcF9j4NOTze
vXjd3ZU5PLPu1nkTK41KAG48zw3fdgPkNHzHAdhmqIhlsHLgRbNIE/nwDPSOOi3HITHuAj9YYwQ0
j+lKG+5mWOtWkvlDKQzbitM5SQriQf6lzbDN/eVmHXitg1stPVMs+/YUNk8To1FQzs5k5d+It43f
5UModyFYYigWZQUJts5c2QDq++bnTWU2W8GPvNmgaMD+OuUn5rAUrVdjww+gYW2r8LJ85QR6X7N1
JKBHRV7tLZCXun3TX2UJtr9tOd3d4mAQDM7nOoGJLatyq6fRObmQwePE5gn78JHwxu5FGOUwkcr8
G+C7KF0+BVHV2ucoOmgEvi4vuhAIesX/knyGM1j2vPCllwOBglURGTfi4qnIPckugmiITB7rEwIB
O+NRq7phUIDM8tmvjbjXCxlpM+u6omZNpajXPq1mAVsiveK+F/gzX1I1jfP1+6ldlpbeW+BJFxrL
CXw5q/CcFYRziRLIUPLizErM57VMRA7SKExpHdSvhxKdcJlhCgXLA+fD+YVYBDtO661S0WhcRkBZ
dAmM4rvtv72S2307mlXbBNKs19Jd3/EufN32CuD3buOexrOT4dsNvGr5Xnut6UhPBxJr/Teh4kKh
2332RNpq4+bc2L3s/TC1JTrsBti0phpk6RlIavJY+o+5WQpHxSIB4b3HWotfcYEyYs62FmUK4xrv
Xbaaw0yMak+NYJiFukV6KecPFm8FRMeKi2UGzDlMLBCDhoix8wzO0Kq75dIAsbSMLmmhK6MmrnZY
h5NlXICqdkXAfFFIzPbV+uNC1nmKsoijp/jjJGty+PuNbxg6JWsrhrUSINy6mGic+O5y/0OzVepA
qA5ZJWSJaHv1P163edqHD2Kjo+JXwd5WmBTVKrLS/gqcxWgbyrCsyyVhFwLTpm6blNITYXk6UjFk
+2nhuQTy8ebqtHfuxwcPplkSqJITqnQApR7hB2eJVHN8QKEWIXG+Af9eX3GHwKtFBko/rKOBtofU
BsqoBfSIY/nfixG9N2mIHVV4oT8lUNJPgNqzVNm/Ca7uL1BOzRbaPMweK3LLGZTDCcrT2QIOVrIb
MTl19wqTojBXyvAPCAESsb88xcd9BQqqxY4KkIgBcVIONML40vFxpY2bVFoK5+G8cYPOImBHfECH
rcfyBK5F6yWYyMXvd6ScKTTGSSjhB6Smjv16iD+ryKdTKwA8YlmkL8sw3/hzi8Vh+FmJbm1MYmym
PCSJkPtsUKDwRvOZBayeVi5YQR8TINl7Agz9CqhXgeTvouj69zmE9nSUu4gpQessfblIQlF6i5B3
SMcw3mliEKqZtRVouTB0wkLPklcS0pNFcFRZ4jFCaiYXpKZzyvZ1AVgipOQfFcu4txK4J6F+/Inv
FGPBV8Zt51Jsm93YiNX+QXn6Z4BmS/lk60b+MLXi7zw7vQn9udAwdDfg3i/CtW1u7+/jTj+qVj7S
ThoRZiU1ReWLjf1+2NdpBfAjxLvA+12uubN/Ug4Y27bU+gx3Gt+QWihK/PPMr4PrVXSbeSQF6RQy
DH6KHCzRPc/7N0zHucfeE4LZdrWp1/NMqCDuMRLJOuiUSMUfeCecec/+ZXi24x/kz4EjKpSeIUqS
Rjh+VqrlTEnyvKOu4nWM+hlVAlBHZoIZdGfvjOdQI9VQxE1B07lSJk6LYSD12PmfOzgTCIw4W2QX
4oiHx/z2z44o+VahoBiFWKyMYgluO7hPSiius5LFpQ4fC5dYLjUEzrVx6NR4Yvgky7Y3PhyYTWZb
JpHe8KswMXj1T5yo4qiWYUBWoyKKRo4sRiFJnPtHkNHdrx25Qf12KGFiM/2+EltVm12jHPsqYbzw
NOl6NvobDwlftt+sndZ5KPnTeORwlBDoNvR8VuARSgLzGeWUob/Dj8wIlm6Eo9B0CjWHuCQI93Bd
ii1dg5POjfuyeb7/LNf+I8oufrnWswI4Pze8MAlKp0Ngv51ffG/HGaAmChaBtNQwGLxxBTdTd+gz
FCjMnzm4Jyu+rZls/dFjbIoJTTCnhOR+zgb6FfcTGYmHEb9/t94xp8qkMEKuTWDfkf90jP4Q8S05
DL0GLaB+YJABdjWQ2VNCpxlOBliTubLSMuhULQwh7psmRNGu+rlHpfja9/gRMRnSnyVIqkvfESP4
DqEv4XQ/DLLBiSW+Ly3a345phEbkuWkrFHfwsQL9PD3X/7RUDGrEKADOiROrJ+nGOJaZqoD/akB/
gQubViWOrxMAYOIcSrVcioIj8bDnmuWSYGfBmFlkEujN9wZwW4iGj2mByO/IIt/0EJIt0tztiRdG
rPoJEO5G1sJrgz4XHiZfmnNcJ2FoWmcUo5hi8dgiaWu+INBwdr99WyhPkubhJI4T+HAL0RMUnL4a
dldkGX4xBtFfQ+h9FOUP76p3dmTRSbJkcrz3m7FtRcIEH5L5Hiaeeoe+J+qvozw9Xxy3lvTDr+xl
okcbdD9gXxKn1Cf+vfckRUF8EPGJaaJB0H/apQiHXutSDOn7LAPWWb05bwptQa5JIP56KJ8u0S6l
pI+qpeoPMNpty6Dk1QQ3SZ9xErDT06kSuhlMVqiKhuunE1XQmzJ4yNjDMO8Lx9Fmc4YWF7ClCyuQ
wqJjWXl6DQu6gCSdsZVi2yetfkpZWpcBz2kR4wHWxv5eQ0xZ6z013xOAMz4+Q8mLlKOrOBLVZOVp
FD6wixjKoF7KpDDixO2WIfCmHFVVsVSIfzhwAk0HuRCrhPwQOyOufOMNXPgp+6Abl8arxaB287j2
sb4LpGEhj3IdznyymVh9NznCRTTJ1HLjtNb1LeAQIB5GpuVpOAylKBwbrg73F/WYqjzhdGZPjy6R
ovQSgUKpMTO7qikn8L2xzHJWydq6GNQZYUPjxxAGeNFGsyywLGlQEZ2WK6cadPRRcr568CsnINML
XFTM+l3Hv9dQ31zA0eeJ6QsZKkFoEmNTZU5CfrsYz/ki7EucQ3bWhRHIzn7hbENNMRvHf3xmSy4J
TLQAf3+q61KVYelWYBJCxiloOT4dRrTp3i21dWIu8170A3PLsRsRoj/e6S/ahWCTKbQVm0nAP48A
GUDH0m3vuyQSSZ3zRyEKe2Y/+XkLv3uQpruvcvJL/UqvJLfTsnZ7VezS6/LPe4s0Zea0xOshdZfp
XosYL+Tb1eVlulDyIqrxVuAJOUML+qU/ipREsYdFxgTELximxefYokouBitb8sOrtaQx1Uj/7OoJ
8XrF/+JdAvCWkgyiX06/uGNnhPYclMruktqSJIha+oFd5Xrt0RShzdDBPxgsuoGnEqMqnJP8X8ay
SrIsHXi3UjrxTo4GEQ7utz6AUCYJr6mhtc5xLlNI44TH8W1L80n/pevgrr0qvpoJS7jk33WflyYl
6QSpSLOO3dAOhoq4ygfMdURRHiRQ/25H56/rWegtPicmFdwxLqhjl5lMp2Gg74APgVe9dhH8td1D
ldsJW5s3gyx7KOuteUnE7XlOa0kKyp+Q/zKjTbArXrzStU5J/LG5T6pRi5yUbdtKJfpm8s26uVLW
/rLzlfMrkfEse92wfdhbqlGhO2NTTYsQ7kjhXtAseUv3f1T6p9zdmIjQSSsdGL4NFR267c0mb+gd
UwH8f1duWf7BwPtggokgP1EPEvQqf6RaMGxxY8moDszTHstkB6NcRzEH5J6xDvLGYdUEDQW5Mco/
IA2vcv3EkbfAzTaalSsczCo1Po1MuBlxk0z0yUm6EcQO7yqJmLTPdQGGGzzvKbAkua0yoNtbnciq
d8dJeM2JXrDUM5W47c5KtjARvfQQcNYMPOidVJS7wZASexZIAVTX3W3SOvMBmco2MyKPmM08JHeQ
2yOfMDSEtFcJoXjRmLr/XrCKstkmB8v7QgX1Of4YotUz259cF7HxiT/tsIt2Jh2kne4WBL6Se822
CyyIUO5zO+rNBZ30h0ohW8fBfN0y99eS3tt7/alxBQJ7Mybykg+SXMB8cnqp7T3tVr4QjO18RFNe
mK5h4616i8rlC2/qas++dQEHQSrpXAN3SDgiTf0+rydlsTe5DFHmELWAPAdUTVI9BKK9yyu8Ml38
deUHQfkCTjxxtq9l88yoFTlz1+prMmBi+GdY5vtygwon08ohqxEDgiqUd19vRJnNNyX/sf4bTIIs
2BjxZzyBbxqJyLS9/KBDsOhYRl1K3DWAt7+YVPYIThznv8ncUh4WqzfIa4KRuDLSQ6Lbro6DoD9N
Z0DLFWHNGrpRYrCUty5CTUTGrpaxWRKVi0GXX1oyciKlxCwRYsN5VkkQ1yW+VizRe6M/tQ3okGp3
ZQCrONjSD0V6q4wUMQ0+KZsL127vnBAXgvBJDnnAeLwIONPIO3ZZNrBNv1QoWJSB8zv8J4LE3JMJ
skdf7HqSI9Hqkr7b++PrPwiGqrEMVQL6EErLN4F/vGTH8LYy8AqZauWJbv7aBMvxkwo/QtipPNyo
tGrT3u+jbxcrIDIMggsoYBB+Evk8kntkOfMe7TKcoJJA2Sr23low6m18DCTRcbff6WGREviuP5Gu
rI+o6oJ02C3AD6lVMr9PmUbrdRlRDqIBz56RVHXhicNNrCJHWNlhQ7RWlZ8AxjqQaEt3T6YCNRqh
6hq3Jsty0TTs79TmHKnCSVeuvsIoIQrBcoE9o84P0kcJuFQKQBSmzZGmSQp7iheVwhyecOi214ri
jsORaezpo+mNnwKmz7NN0xk0gWDhSJFx/RR/oyfAM8IkFEqsj+g6c+WXui/CGjbpxozFWWb+jLCI
KAW9UElrKf6bLKDt+dIcBiTDyFdAgd/MUGgjCirzYatsgg0CLfFXJXhrugKPmrbKYkVJO0LZDr29
N0plEMETo7cEK7mwdMxWm/zkGazldfeFB3pVT00CPMHFida50/3f8CWK/u/VH1Dhi1n27PxrqKi2
0eOUv7lsEKrVmTg3E+AY/Wn2hYz+4G3n+mmgza2+AyF1HV4NI7itB5T0m1voASXKsnPHxi2I9tfY
zMgWEdjAKuK1G+stJ4BQVEQOKeT6hlIDxPlH/izttLioCsDhsrc51TaxptivWnbemVSSGLTTtdth
9LHPyE8+bTkBmITNDZBeemlNFA0QguqhwrBS47mKxm8MFJwJDkCC+vM2QMKTuG+di3oV1XNgCeWv
XfZc8pZoORYer/4qO52/ZILT1/YcbSsedS/mFMeY0EJ0+f8oapG2lIASygwSATroWXaP8CjaD+qd
d8IbmfYw70+d3aC6h+D/yFVFyvfAYDKkVTjCftLtKkDxMRBaHBJW5xYS6dMKZ85cIRklbGdvCrU6
S8JXXDcSiRQrlKl8E6BGz9coyg9rbipNhzPMp9b6ZeBIeVRJ9hox2RC8JOtMRVhLzpwGYOfo5Zr3
L3JeBe+VgCtqtVJSvipJEiciTcF4/TsAT/O4HfAbOmrtSaEWV7ycsQ6cDORx1dov3QOVbEM4qKsP
0vKEXQZbN/EBbUco47V6Y+K2dQmICZwzWtL5m5OFt9fDT5LB4grFltqJUgbhGitBb23VGzNWgjKQ
Z/dEdHfWAadebfF0UxWUG8CuwvymTnwgg3XyFpYvq2cAhPeOBXtp8Ke5EwIPI9Mrcyvm3AhlKI+g
DBtZF5T33UWcHMykczaqqYKFm2DnexPNHDqNuH86CQFL5m92gzOkm+zIOkVUbqEuVQguczxpTYQF
XwJFNxwdxcjJ8Si1lvNH/i3JkWaoCY6iSe1C/1OFkXFRAfDicpOEKA9gCam3X0TCHZICCOfMHCa3
3DvGXvXinL3Hr/hzwW1gKbjIYeQdDlDOR96tvjAd5cHjNl/2XXcil6HLUrgcI1oLaXxtQljX8PY7
KAyWgYNeMp0ijng8wTyO4X9civged3ASkOIhWJa8+xanMUoNQ6OMepgcX4XcjCtEGwWeFfFA3ogk
a+KOm6eLTQH4iXTjYed6U3W9xu/w/d/JRSR/D2wfd40UzA+EDX1mZ3ZJaHR5TiQftiN6LF8KllVK
KymRYKDkWINv+plSieELTOjz5WBRgarQ3sSaNy2gvIhjJbm4Z/PmneDfkMwABdXpr59oZy7fpDyr
H6x/AzAubt4xO2XUZieVZfkQjpN9vH2Wv2p0a1Bcvlp/fZSQv8r6ky/ZMV9KbtgnXyzY+p/DxMNu
H52uKDoNv6DqbVAEvDaknXMecDGiQ77H1IKReEwyY3RQ5/DMkVdGW21SI65pDKmxJZNoZ/1Gz1mC
lo1zZFl5EXm5OFYZx5ylaD0+nWqXFOuAjAG+Knu5FQOX38g+ZUzUekt8v+dVlLXHA088xnbf+zKm
MKOYm8H+nDXPdLmRg/fhFjY7bz+rmbaFMpJ/IdKgDZNoHl6kdNh6L8/gxd9v2bI7X/letLXVxZKz
0rUr9XF5PXA131iu8sR86uHSHf52qvAkTAPHqvw94LSHQoR2pl5MYBLi/9G0sKTaa7QSsltMMOn1
astDlCNHANypXwcOwesG+2t/klcIT+gnHCwhgfz2JQ3fP4S65x+oooprxnAaryqibPka4IlVM8eY
NCzSOHt0vgJYqOqQ/POc1JxmRpbowG6HDHGGIBwVli2k8OGlVeuFACRY+7bLbwCI88qR9QbhqTpT
EGme44MOoPkLX0FH8IedfHRZY6s+5UaGTulv73DO/hqmkCcT6HWT4eoYvcGXG1JGyYrk189y5bk6
lgk3qLwbG8Y6SZ8rfKIjt2HomFMNIgUZNqJy2rL7XDnYtMnNphMC8TLeLtPtU6cmcEUS+P+1C2pR
faqeaw33Oy8w5LS2I6xFfqDCV0G4qYJy8VYRoHCXxwnUKvJ/zHlGmuMhU9/b7JC5pIG0R9lwVMtZ
dR4Kpfm9qCs0ZjQzky4ifmc2tCkLij/A1KuNYzvqF+fdimRBV7z4GRQFMP4HBm1SsOrk/ocm5Bhu
1eEX6sVfjPSSpsmogf24p1EOlmnXzUsvoEDYdBLgPHF5RwwgZEhXw/ucbxWeAsVaXFdzS2PTOlRL
iNMBPs7m2sVjOnRtt0cOmjOnbZuvQr0siNnj9SshcscHFAq7I/npWE36fN4JCck5ANG65LSIrFzR
P91ve/lJpXAfyE9bke3K9c44sNfSWRq175GZKlLgUpC/fy+R5FMe1WMlQj/UM0v60P5n0TJ6zW1F
SxjU5OhNVtSlJFfsswWHNw/TTxiVlYdcqbg10Z8aR7SkIo/h2OOE7c7FnDKVB/EusKm3FmP32GiJ
YeeEeKrBd1f4UVzdX6DERPdrJp1jVc3HLw3yG7YCshiCQbFCiH0LF6MZV8kMOO+njuMWPDsggdHA
vZbPGPAcK8DQpnjb37YQZRJTqf2u37R4sLGxC247r+2VBaOUu411C7kwSz9Ni3aCFzYL2dE3zXe4
MlangiwX1cX+0WxIf5nMsTOp4kZUNBI8H+yNUnYCU60X41m7Xb+J1cldJu0bnqx3S2Gf2By5VPsa
9H19KESmWOfs4TM/HhjitCBm7cxDKNOQP+v8qFxvL9vtO8jUT+t0564j3f3BlVLR6lgPxSR2kX4g
/HPzeb6AwgHYsuS3Mg2nu5t8L2qBetJ6oU7SKNcf+4zpacDTusGvc0x7ggE2lIdX1gfKP4yXN9DZ
JXUvUqEqePjoqVZqujQFRkxIYkPQEfBKPn1StISGcH8TE2rOZc/tUMd9pZcG4doTSG0oXL4MOI6u
EPlPwS5MHe6wDc+mff9gaMixJVps7acO5cuRx9ntUF2ssY2tE1Yl2t80DOlEELgSf0+ueSbCf8tR
qfbBYdf4plARe4eSq+LBTdag23WPq6cHzaghux3P48KqKIe+bWB0nxP7xl6uZkk86EaFggGGUDg/
bKrDBqY9Ee+bE3x5nYByorTMKGEA8kUuUcLXlc9E8V2m4G/Kp6pvorIoSvyFua3DwvSDRSKpi7t1
S+xgwqcS0ibZngpqfoj7+JZI1DcWKY3QfCJkF/YaOd7QllbrawKE3VRbPQ5yPmh4KIJV9zWYQ/h3
SH2xbZoyCtqsT+8ZSVK2mVffY+2zWt33++Y5O3TCAEraUXD+9Mo+no7GuF9FMrIr9VvJzZrSpFNk
AJt22ceaagQtaYh/QatucS2GbsdHLRvRZrPEm6Bfr3MZBafTuScnfCNHDDmxTLkr9ssJvkZ0TIHi
lxNTY/3iuDWODt0jIYp7sqLBW+VaHqpAEfLw3jqnQZeqEUlPfwTwvYGNjJ0p2IQ7pI0OVab49/qz
UbwhYYPN6n209JrjYF0XC5OZJN+6jgev+5v0OvBoRNTHBONeog7mJWm0YapChNt1Ch779DL/Dmca
BlIsdTW5omi6P4DX0y87Etz6RsTmHdRmM/DoFpp3uU2IRR8D0hlqvLzo2txRJiEztq3uz8iiLc4F
T43pEn9GB4zj/z2ICF1VdnsMNatrPK+wCl4rWy4xVIsiLuCQgxFkd54bNEOBoRZs10+Pgy1+F8NR
9xeJwdH8E0e7dqgRtLIkMBApScOLAjJbCLUF1eO2dAtvPJJxTii6JdHRqXz5mUZ6bKzq1tzpDa/d
BP95bpM+wRSLqx9LdnabIwdff5YnI3SHPREPH04qK0L8NJFX8CZLP1TiAddKQtpV6x5b3DQ2Lmy+
DKtQAxbDvqd4vr3X7W2et2+CJm5zxyE6RON0QD+kJUtpRoBVjmkMTdeXQbakqUiGrKYhz89hkwr/
EX3af9ZhfxPLZsQepI3aSwSAhfET9aXwnOrJvy+f0a7SE1NcCeOpMFBeVSgKn4EecxLF+fs9uXvT
ExBH2UFdtHqqs99K70LVfACOwi4FDyjpSJFz4zILEmFzWdjI5i8eriYHO5rLtxZV6iCIi4/oq+Qe
Zsr9wpz4qTvUJDSgCnJlXqirlC/htgCjJVMIBuBNYKyxwNq6sssXPVTXHwm+6Vq5Uu64SVU+g8Qh
vuhtw/ltOdKt40kdnNpMjmQPuDjp7s77MIyZlca+pF3nOmB6VTXAtyjBNC6xmB2gDBKQcWTY1bs4
NKbjJq4XkzZk7oM6IX90TlCPetn5usa3zIEApkTUYte251gRSZhhJUV9qPbnHJ3zWNRGXz4ehekY
6k4oK8mI/D8QgLPu/mrfjCfen9SYJt9mY1bq3EElmr7Q/Hc374Nc1hthE4CMqTd7AAh15+F8Au72
PcT/WiHxdeyHXdPq6dqutS0LLRQEi2C9tFKi6NmeFi4EBIiWzT1KEUgaGya3Ggh7BSIgw33pwOwr
S3orS2AM4PW3LkSDFJiZaWoJdEW3q+86IuyHXfrwr/L55jjDiTpOM0HsQC7Uh/7hlKDImePY7LXV
k0KKYQdapoH2AN8muoRKt8QEFE+pwFl5aUesXExo+9gRv4ZBNxho1GqpdbA0mEEV8yXU653eTWvz
da23FN3LF2l59fXpSb6hCCDMY4kqH/XlMcIk9jFHo8SSBwrs23uBnoDbtw5Gram4lgs0jL3EMo8H
xMXD6nSY/7i/ruoDBvoIDk6n0U3WpNC+ni3fwqTNLYhWRDu5wXGYCAlAQMnPYKp20h8qBTQf+qrF
DEythJ0uvrRpkBuESEthxiFn9qEBPV61c7tFpIKLC8nY4n8vlL3a0Oe2xWVQzSVxENmCdGYhNlOP
ju2vUZOb3SdDNYKzTL1ZTbG+c0HcxeAhSFskiCHJGuJLorDULdK4PRQiy0AUju4uKQYu7qTcU1jE
aVndkaBpZnJJbYGbSfgJXKZDCAvKLa7tDIbOqk0CugiPBgj3zilXAuiilvyqG1CmA8FxR1CfLaYt
+6lAPJiTJPIf6LYnSh1q2RjjyrwIsjDkU8O/mO18G+ccb22YQeSaGYulQnarMP1qr74TFISSlJXo
BOi+z4GlG3cYmjabtY2dyYHeiX3EmDLlzgnUlpiK9kMYFcS+Ff3Tmi1x6PQl9NDXT4rra9kijIaK
fudyRZWaRNxFWF7CB7M8D2iwgOfXIibiQsNGcdiRbZUrRjyikLHKdPpCplsnyYpHeD2MkxLt6oeW
h8FAAui08fQ1PX5k9PUj2FPQcmYOBmGjG7HcMh/1JllVAIG4eLebrtROV1JFF2yW19LTEh6/DN7j
ht0aY2xdqKiUD+bmH3y9aLAAt7SP4CSiDLvmDKaYc0cfVziYltQSjOGOkcEMpV2UNqSaIuAm0EF2
hpnocfj/r158AGout3YSXPTZFYG2XGbfyorsQIZYN/8jJbUJhGIwxtCfZjuDiUTUDIU/+/J6FiGP
m4kVztyVhX/1uavmNxFSLaM9o/llhoQ8AYZ4tNJIbwZjWHRqAEZMzNuvD9aGTThGtGVn8Ga8ygwW
JDXq9/j8KIsVd9vHM8av2j7NmUOT4SHiPlOFBhaEpkg9amtKw0Hooci26rfL8XqvlUaUgfCUNw7g
o7Uv8uJ9QBacnz9Kx+Cg5TT4uyYgheBex7WUiv7Cy5MlUcAuVTLBn0YW6+56h3SpyKiCBRd9wfz8
CsHr8RN2W2tu/gytMAegAwb2mG96IbMv7PkoSvBdb0vEmc+yWtp8cizdmyrbS1wcX1zVMGtG1fT0
vJT90MYgi+ldZ4AmUV3yYR6DhLKowTIR6ODV5b/7eEa7CqX4Fyq1NK/ecpyqC7hiPE6KSafha7eh
mro8TSNzSg8lnY/cvnEZdaHHFJ/wXLW5HQybszNDuFuh1v+NCx5WuNf+rvEEuC009TvkT99Mqvi3
KJb6Dki0Ogez3TpD+2lyHdKkXCrvbr09sKx6yBi9ZzFHNpIvyOVFt/Pi0VjU+exq1NbC4Jzzgiac
uSdKeg/Y6TOZwQffkTuye7jPNYLr+4XkNbOjBa3RU447EW8hiRQiBlfgzEOqw+XkebkFiAdarwZT
WcVjVcdBy+UWUIxuaUTVeErKdfnyCx0IX4dKJtGCBgbWsUAuAJq60ovpeopG26z05FW4uuX51KJC
URLnfWVexFVGIaZNf3u+LkolTCD8QHomMO33JcKXmYHv7JQCTRRbtRGMdgjKMMRw0r6VpKDMOsx1
GmCCzSbM23KF+7pBJbQquvrP7ImcpevMO2AcRXvoOEM9t6gOhpbU4T+kHcAVWx8N4nDKtgQlf+M3
b002Daghb8cDF6l3+qh/Cm2FDmMdySOYZ1tVhNhRVss2p6vRgDC6iyneq+MnE/FvsJKjcntaZdaf
i/Lz5mp6i0awjuRUEEFY+0XcUlHVh2Do6kC5fabNQWBULiwmobJP/dbjU6K/wrxjlU+cWN2pz2cQ
q1fqU7CKxakCU32okuaE6UmA9PLMX9f6mAqYJM6hdQoGEbPmf5U+8tYjbEq9pf0tLCfJXPnrtNdx
pemx9Vf+0jVEHPmnAcMfxvFtYQIZi7iWaHsaMYYcrsY/WKxvI/XUjo2DKU9ZQs+nIWMALDINNkQy
ReLyK3R0WVAo87jYBy7fP1UdMvsIpm93jMQOk7J+GzracUBTLcLyqo6vvfA8+XCg8FmKUNm8RNOd
neGMWQeCV0aa9gda2CQsVYlqWu2XwM4dvZTgutdpPr/YbgRMrW2hIIN9MyzuD5x1odIdjYaoQjYj
Jc7IGEiyGYaGT0xQYChe9Zqhe3fJnoZNQJxMVNXLDNUSqGJHAThLgSdIs7c+1Tg9zokGz3gZ81Dy
q7GLet2j24RbYsds42/BHdaBrAbgYpmwaTo0G1DhJgrS4sDj6EBhbM/GgAH3UJwyVpmslnXYCfEc
H7P8iSrfEOp/R+AZ04ae2WL3U/oLIh1q2o+0CBABsjNEJEd5+4GSxuLZexcPCOngA48JpTPzaZMf
QHQeqQfHbLSBsTUKYnrwMxnkrwcVbOjDUWyH18XtNqP7UAPxRFVlTd1NQKjpABWgAyK1CkbjXhzV
AnqEiwzjRNGqQX0rF7R3wuQOQ5wsvsbbCkd4ZUAoa0BAbgATv92DOhmpQ2WV16GiyJGZWGgDzoHx
e2Va5fVubwwRKfPiOQMqnOvjqb/2Al6mH2Rptwpnbbewfdws0NukBfXdS9tKybNfHcBmL4fZcgrp
vvCnzBXhgH+hsRz9Q4QmPdpXMNf22ysVDCxEHlhTEC9jjpyrgTeQ/5HD4pDiHShi3mM9XLPjNND6
6gGpbwEXMag68JUG1hi58/s+bQwwWIGCBeY42Sait9vTZrCT/M3A9l27hApKI9e9c3nmS1Xfu3fs
aY3eQzn3+as7N1kkPxldOALUwXl9wmtCFQFa7srL7nsEJoo7Rg06vT5uTFMZOBmkFZtaAWlPE/PU
QK1WKm3PYphHyOemWQxlVP4flB85DoyZohafXH3Zb3SFeFYTnsZ3fjU4bOuRjBp/xDAxSnyiRj4+
ofPfrzlfcEUAmC1wIKrFpaGIum1jIhRDQxhNSGn7stacAG+2F1mFSW1v4FivHWcNVoRcl+2M1uqa
iNawy9JRtbuGSZfjwjZTFbSQcgj0fHRbthNTM0vo9gY7sve4aizY5Be3749qsaJ9x54z6oddSCZw
Fjf9bHeO/fVQ/6zYtFRxmL+CO2EyG3RRAfFBcrWGOdiqDzRB+4TdTLReX/3IOH7FmSaHig/jT0kv
LWgnEikOWdYDjml1L00so1a53YdpX5MUcSa5EhFowJuN4WDa8ARfUyoYT5Mg23aDHhgUnWgq38mK
xfSLkadlggibiNWeE68tdHgqo2pBo+XSHHpR9qzWMO1qlySTGz0TH144SWJHEv0H0xEWbXvL632V
l2ypB8SvTMmMBG+VDhhXuK4ruu6GsjG4PzgnbCSsKhzOQO/pTFp0OioNF6e/shMeGcW1JPQv6DnQ
I4WEhZnKbSXMm+X/ZmpHJSP+NWZfWTv8rMH1626ZDnZ988Pp7doMG3eHGn2mH42jRjIQalRAZJQR
msypJE0RrZ7Xj45aUY1lxXt9882i1BwB7M4DbKI5GW+dV07bVJM96uvsAjIFRMj4C79sXjGYWZ3Z
I2t351ArnIULfTbtifMNh20nvG4+C5CUj1BHQn7D6851rkZ4DNkZCqtCQX4XmY+RObj6V8G5MhJZ
91PLnZf7N0YAQskGB+T62z/vlkF4xtazjhDDsiAz1fOzNALuHhcO6gLGcLgVquDKTaF0inGsfF9T
WazCnVJwARj0QdeW6P2Cgm0KbIujlBk0e+F3Py6s3FuAX8z3MQvZk571QUgI2dfDZ/vrgqwG8fcX
d911qPMewENlBpYS5Nw/P4nqv2iE0M4FxjzJRe+n0OtZUOjo8lw/udy74l8YrehUptfjdn1Ibu1X
fB59vwv/+LODCpO1YTHCwTvtCyBRSXLIksgcmk/yVIip/jY08E5aPpRxLZSe9LfKQjk8TT68Znuj
61f/IQDjds7lMvOwvix9ZOeL7LI9y8F0HQzlsGClTxHt51rg4RCaNLF+H8AX5Wd3cNnIZ8ZHeo9/
iWAkjIBBea4ZxgAZER6nBUCVIIzMg2Cl8HNw7KdC3HYUOM7GuOKYY+4REizTSvOLrg1m7Te61gR7
KPMZGeyoMhbywCRFyKrRyp2dVNrRw9tCcAanf9pNwiowwJ2UC6fTXULgWT3IPAnD8ZMNcEFYgSsg
0LWVK0adYE3vmlZv4lURKAYJVHpC2dXazsa+FKOvXxjwQogUPiURM0kxYJvkjMOZr6Njt89tk+cw
7+yeA3HyvpK/PqOAVfl5o9wgvAi857EtASUin+/ErRzrY+6ChGSyMv6kAT4H+JQAdGjahTwIVD6b
RJgp+qDnqNn53TJZGmYI8j7o4z0UQkXOX4IHE0/0xmj2LCniH9QO7nacfRI98gFjkNvXWYyOIY0X
UI35QnYRCxOq0DuwyoPh24Jnjv9UFs7d2KQ5A1mYixCmsWRnHU9BERak0lqP6Pzry9Bm83va9d7F
RL+jl+EwtTH/v7wfvLASsuAN8hYATgZGkp7bWsc4eq/b1hBnGGOwHzRtlOGHKJOWPAMn8CXYaqWp
SA8DwgnT4A5VB0BaM+T/u93aMDbBf4XQNcJMcjcGsxIhdKqVSMcPwWrs+IkI2vrlJN5b3zherq8T
hveCaBrKSjqIlbgMzuJ5JLUUMrnMnyNjgTp9/009J14PZL4fUPsrpAdoo4x+7U21cF0CwTuaaWF8
OGZmoqVAb9RjGqUW6xgmy1gun1InUlz2acBLyUFrsxiZzVGA0rs4YxW8R1dIeg0DQpJczzj0lIXZ
+gPDlxqrEhefxiDPLfhtRvIm02gYPP4zbGi0BSIvpDtFcr5CpPmThQPezed7AiZQ2VV+0C8elp/r
lMRB63+SRJ6l8E6L//OU3PmRfBSqeD6ie0YBOctgWNU7kihR0wsBJ9xN23vOJncqezxC2NTSdhIv
4vCIWMtv67tQHpNGJXOHRCUTZArgbIlCguEiqUy2/Ne6Prv7TJXde/S/mFPy5WRTOgYQfBkF1BR0
k8QRi6vqDrPcUzSfDOx7Qk8A34bpU3C9RfSGzO35CQlXOrSFqRb3JXVFs9vy4hlsFZPceVQyeLug
D6UdgKQ02nzkM+6z/akbP8Dzy1XB49LUjYLt9IpSa/OJHq+S4kG0QjS+D186EucW4rbu3CICtv/I
8ChvRPGJHcI2yZs6ajzs737e49E6SNbqGFTKa0wsvy+BpzpLYG+EtTzNMSBE7goDIxIKQohpWIM1
IAH53pFcXoobACuId5HkkrR83fB7gAIW5KAm78KOOXdOZqYDB3I1pYgsoDrDdW0PLxlvq0IAMZVA
iOsfzNPM1FWm3Db8Qq0WdaJA36C5Zk34rETYvVRvaWOrHToyapPicKr2BCQJF9d4VnccfsaEiFsb
2G9SxJs4OX89m5+YqwYpCYUCwlYcNcqSEjDDMsq8VBtUKu0lQwjTKkiJZvP7Rgjo9Of+WH+q6gd+
KfTj0LZjoVEcGMqjNjRQiM7fawK5T62dsCIXy0UKuwc2OtG55Ydc1R8l3KH5hlUQUXOJZ56VUQdx
uAA6/eX//xrRBEdI7Av+3ULI+qisLgSQAA38wUW/QP/+L0o2CHUuSfd3Yk6RIFuODsOh+GrRzjgN
poVgBNdTICcNN4zMhTRKGcP/hP0qAxeCS50hlCI5lrKhjGqf6kcjXVhPbKt1ULMtqEZ9qZ0xss/c
/oezpLEGT2MwdZs8O4y2SCgLnLkj+DCAD1/xn3BfohXfzkN8EW5H7driZ6MIkKaxQKAV9QGj0ly3
TCX7aVZigNKttnwr8uVs/jdZXWIDFk6T3Xxc8VsT5DfK3vJVlhZLkG48XM3PF/z3GthmTY5mtAtL
BmJX6TWhGHuiiL6xVgccaX+lNSo0HWvUFWZlyQC9eUCeF1SuK5g9uZAOeL8XTXGbRvyRtBMrxDJI
11phjmt/jCwMzyrhbNDjEfWrRKgZgv8ivL7Lak0Dqum7FknKuvDLIcI0OF7MKxrdvnMZg61lP0I6
e9N0Pl6NtbvyttFX+17tVc823QNqUoXv0YsxIecLk/SvmkVjIgQFx7eaX1m4tpnPDU2Z45USGox+
99kfd3Rm8XB9eh7AzTz1lqmXzR7BfrTVPugiTYq+lvigjhUTw3iB2VITS+B1L3HeEwJYC0ucGYCQ
u0JdpoUpcrj9lDlWhKBPQ1aS7hmUFue7antnuMhMQ+8wJxJRCCH96XImAsuocq9sUilkfXNEfksy
NFdOFSvXBYIYlVq+JyqMdl/aq046Wu0jxm6JQKSCIHAaAxrnntUXSikxgD568YJ1fb/+rgggsvAE
UtMBOISNRvytJ32T5iFMy+n8MaQwEdRouS+LkaraABnvnnm3Skd6zyFCqKrGjvCsfMbhPIWwtAzQ
JuDMRES/n7CRzW+gfSeX6+cRCWKCzhJotx/Pqx4EjH9AbuLV0qkXmVczUVqd/czuL9xaTYoOmVcR
ffnRuC6MYqxNZKgjIaukpYqhILRdH+NMLBO0+dg7meIUPC0UOuO5FZikI8bAJNAbYOtGZr2YYEjy
aZziac/ESX8E8R3iBjxpfDXrKRdBFbtdPPApBNwMx+PHFivkxC9ElVx5Jfn8UgjFKacsWgf+buqS
B9vMjzFh9b8S3k/HulW2ECnAF+F65teyTlJnykCDNZU8ATQJ6iXTZJ4cPnicJokbh6gdSAH2OWTt
Nt+Ljz1qppf40aCRzrFhLSYSU3Sn57qjNrS0eEEn3t4uWgJqF83vpOkPqW5woPwc6hS+55pFMwnL
v+isIaHthoMQnSlsw/rLeYnRxa3W9mzM1o/ry4z9Ps934XzulAP7A6WcTlrN/3P2Hfd3+BEIr+bF
K57f6rqG1fcKUQddzR2zdjJj/xUn0sZNaG6Ebz0AWXIEcPXsd+jN25FV4LDCiYQmCjWubC2KML1H
BSn83zcIbXYnL6kWJ200cFu+Qm2o2SCPx4J4nRcQehq3wip+PCT7ooOaA+82KAC17e0KEnn/fB2E
tNWeTYi0p2rQNiHCnDvgaB9du0imN4NoVoaRxkeDcDs1O7VGMd5yzDr81Cf26VoAUCZOjyqdawUo
EWgEVKxTJgCMQTmG+eVvxsxQCOwLgjS78ERmlUYV/LqThLbRZYbFgbQs9jAyWrdCX6jYglgQ2EHt
aBQxXyeNfs6k5wB+oEfIOu6ga534gUkQebQIfxAYI/u8XXZK1MfeP7ozTKj8xoGpBrkrVxkjDXtM
eWAKHVoYEWjUyhsf/kxMMc85oZuOHFX7m+y8rtq89XivmIr1bUtY37+eFX/fVFrIKiqJrbVZZoqT
UrK9CVUjinuoUSFr9HkAcAEcsVa4szk7hQ5mn/e4XarLUbznr6U9TTcA7TPt543X2yDJ4uA7VKDk
S6J8L+MqsVRVTk2l3UHvXnqKNmEHKdbHCwEUH/5vGHqFEfwhJ2NpTjKEkNhKvxxsslG6ETP39lyD
TZtTauVKa1mVUAK2oRKabW8z3iTjDhdfBnWErlQxSfdDzloUIq4tcy4Sd3wrIrQcBOVpzosKk7Jp
ON/gDpgohr+lcNyQtN6hyCsxZCCR/RquUHkvmlyHh7osgcMfWdDMZ8HqguRjNrOAarLQ+LFj/JZR
rmNzwYiKb24ehthYa+5RxSxAO10eUF76sAYcG9w1sv7737eH63dIwHgCnU82Oa8ay28YdD0s8TLX
+uQoNOK75mwSQjM3uU9eA3/ro3CEkB/V35rk5k8g+Gd2hk7bIucblmx5dbRM4Bmgk3RHoioWjf68
kky0TUeW4YjY8bmoq5BJqltDrtdzWTs2XYf4jhMlpp2dY6ycdnooQ7QjotEiB68yY/DJVALjsV+q
KQisLD9q7fSxkis26rCCm/j8vgagTz99AroICmGNyrzW5PN2zzdIPCC6QPWLD+0KqGnlp8AQF3Jp
/hbGaC1NtegdcaFIA0kGcn+Bpo4U14Avj4a+dI/R21FPnPWRffGsV/WuraQMZf4iCtYIeobDJhSv
IiZusQ8C2N8vWTCDB0LtbOes6bT+yJB3nwaifn65SfZ/8v/5hp84cy0JIwqA9UmdXS0iMRDqR/+d
QRnBYWf84Dandssk2le6rfGOHg7Kl7QeMb1gpY/z1Na49FDzuU1KzZxTm3TXtyqNayIRzKXLyLE/
wh1hPi4w0eGsA7UiMNiDGtoYOLiEgc/Iv4en4hCHyy/s/4G33mGSRVRUVM0JBKCDYkmuedogmZzh
PNzEgSOfironEjL788lSB1oH2+/ccpP2fSIs2rnVjHQpNfSwZHMdemeRV+1cA8NyzVSI6AoM2kNQ
uUZnLcpoOU0q4uKBMQEwm3JmvzEFwuz+pvIMwst0eTYS0Bk+/t6795KAcr2kOnO//LOZH7Ir9xVW
F/VgZS6GkLNCiz/92kcPWH2Jb/9a7SPS8gp39uWjdPi7ZBxtkl4oytvKuQO/qga8dL0htj4qGsDa
lMNKZdAQzcbY6sldh5W9gSPuJ/MGiXFDs/+2ZmWYD1jxsU670cxwrGCzUUWdmNyfLs74mgN5vDAU
v0j3PW/g2ccxxY0sttnZMKyELkxVs00gACbFQmJ2le6Mq82p0Azc7XtSRLBQoAdubwhU13Lt83G4
igulIBBTIpVammRYayUs/Mj5E/lHpy06cCp/KjrYbJih+E2OnPXTWVFfDjyoRvq7A/8mXJbipX6I
qLyXxWHrnpFoJOv67Akgech2HrvLbvmhI+YaKrndZ1wyWOvCh+o2tGjyRqI+pPFrLlZ0rXpNy3a3
7yssMThotVhTRjk1CdCia7olnH3gJEdkT2w8e3g78ScD0SMPNQE2VY897T/JIlDoE1T+56H/TWeQ
3vO34hVRdsalgTjA+xLyI4VRkYiPoILCWZMsxXfAOUygu5haWSj+dhI94Wjs3KbosS7+3Kd9iQ+5
wjQyR5ftllXmeH9IMHacQWzRJrislnVgAase4vknFYuhuzg5zCb29ri01hQ8UlHn6D5370fz+Ywd
c5ycwh37Lw8VFzdZUwpPztyt9ezo59MLIOTwfOlv8D/j84m5bQrjX/izTWR1poJFgXtPTMfacsMf
Z6MN6KQlaOT6PxNmwsgwLYlAOl81y9Cc5ngVHk8uVhoORw06hIxice89JPw13LOs3Zc4U2WtrhMI
H7LQhXz9oy/Y1TeyCX3Ja/MxGUnrfwg+gV4QyET9ng6kJYFaguctQCYj1J6pHr3DgJlEPj6sCf86
wHl/8mk7P6rNdXVQ6rmxlexyESneCeuDQbX5YkEciIqtH3EFuljvoRso18nUYg3hOCp+oOcw7AhE
JtD5enKV9bszs0RQCm6hfQcAT44aWg+wZ6eMmj3JnpC5PcseRcvqRGjlw78PwHjlsGJJLqKCwuqF
hov7RIp3b2G3rHodNALF0NyQKrudRrDWExjnYhDdXVub+R+6Cme3KNlWDhBDjHuXCjQ3U6//J3d7
0X6NAHS+OHJmnRkmAAnDpfJtN5QzEh7BLvjgdOKN08MICoeyXfe3yqTu7hCMff/CqMMSsMDpl+3I
8SkHxTa12QqeMAzO5a6AAn1SJXz5D4/aACqZfq3DltIa9bdKZSYoFXwQJygGrRhy3c0Eqa3pulAb
sdCbV0DUtkpms051mTBpqGCGqXONKbLpJ3rPpCSEiKgh7f24xrwF2QZcP8c93zR+U2EDPq6O0tRw
L0YxpO1zkd88V3Qj4WplkpoFOM76zSAkVWAwoaGm9VqpAV9NkLOj8aqjuTntvn2BNlIusO/v3CTu
2k57U8woZAftRmsJPyu6WJP3QIX2uHxZAxHC3Jp+SDcOkNAPY+4J2UsrqDF6p7uSYy+mwr3KYIIH
BQPCbbYgt4JvNY8LR3fZ39V/sbhe+J1jfy/dN/l2D397F0kk7EPMT89jPXeWBGUZ/ZKQPxsPerKN
ICJHQqFTeMju0uGM5HG7ke+Y9l5UtHaWCW16opUZ/pAhUF2dFcvVvWw49yAaaJxJvisNhD8tcijm
awyCmfc5gXDkocu1Pv7mUXZoaXDs0twy2HnPOcOJ4ptJ7lp/lPNQmajNnsQLkIZNP5cO3vMXgZK5
qmDveV5DEEFXAzsoWeYlVw9Rkd6CCmsBwdBaYHxxToCE7S4isRRP32DdfUZZKQqzahs/hZYy717h
jv0IlFQkYBIF4PMB96FVNvHGrNxqsg5ttnwypsFYV82x9993sLU3p2hU/RTV0jRwee3rZBbzuHXp
3SaT1HbKnnGKxSpj/Sv8TtUjnAyjanMocxvqR9i49vXdq6MdMQvuej9yf/XD0FdTy3q4TfQn7VGF
obteifjT1PA/MlnsH2aBIjOWDCu7wA3QnVEmOBVqUrdTjYcZTZnxExysgfuRSBJ9Ozm0DuYmWJ6c
NNY2ZagkuUtJI6RpseHrhgeKQGZYjMq4hBqsADymYBN9F+jPinj9nFrm/cVb6j26YIcppxv5/HpR
M0cAfSGn2iOyFukABVFINK+y2q74LKsjcNpuy6uHbxUlj2Je2BIjPqlNwdz6/Bs40eKnu8ZFbR4S
qkcNgYSblFVA0FvveYRznb+ZPZjS0HwcsxM+g4WNebvupPmUjjo3ASmowuvEh3yGIdIFY+9TVkGH
LSNA6h8LQtA01mNK9EYVJNat1UpA3UCKH8zv3+AoLBKb8Fu0/Py4SWdoVWkP9u4ZWZSrTgrL5r8c
nklfVNy6VgpmlgsqyAfK64QqPzJkzeO2M4RQNSKrUy3JE8PlbFgZ3Bro6C7x3Xd0fM7uqoiWEd6U
5PWAqVKgg50Lyvblm0+10hclXv67D7QQB1NuO5njcs1gdXkqv4SB7W9n7+m4fKY2URJf8pdfqhPT
6qJfQUk4eIG6DgMK6jpzGl/iO5e0VnGxjCGymZd3Z2KRVRTkeqrCLZidq3hUXnIPPMJxAfXZisUF
PjTTIgBmxJH6ySr5z3DLl5vda3IUFqa+zTiRddAS9Bs6Njv3vRFTErjOPWkSPY7C4sDiMauIgQK5
9fIfU1X+uyQZQW8llCxlYvv/Reno3kn1mfc+WVwu0TJOtQQnsQDJawPbh/Z5dEf8l/pjZVSvB+2g
TY8K31FlCVib+lnevca/75FbYrc0r2eWiszwSaFOuK8FTCaVt9/ovU1cCW7vw+xn7DzarUvu7W/7
feyixLdazNPd7rUND42kA9qRRBGzkZ3PxD+2oK1ArVXv6BMUa20HhzN/VpZ9vRoFRnykUbRSAjZ2
QVR4oa5XIWOM+A+huX2w6mub95S6zfHCikvkN7cqV7eAEBokqEXM58TBZbwE7stwbcRaW6E4WdKq
1FPyV85djuRSTMCHmXBknGT89gSkBS8zzSfDZRYa24r+WyILjzlWMqabk39rV5lEaTjL5RiUQlyy
zo7RLZnY3g8k9zanl6a+zz6JKvJI+3R8TJFBp442iIH6b0h04RxSxqCjG3JZGJBNZJTvAq0i09Wk
acY3Y1+zNiTem8npCmraPoYma0fsE6ptANnteIXNCrt5N3jp7fUcOE30JiF1iuPqkvBnl/bsHdpf
DaaPQSpARWQbJLNcyILAWnPe9F3GXwMRvolebAUrlCzpLXVUJhR9SqJBEz1Utnq0OC6/9vMh2qbV
Iguzg0P1OAqlFQcm+DgxPlYZwDn/T+FdoLx3/hg8iHuV6QD99DWWhGsTiQLzKTRuFaoOkhg5Npmb
B4gOUhzAWuRj2NHJ6wvaaPZQqFLUSlSKaOPALWXk2YJXBej3qJZCVz9G5QSph4Ak5FwcCv2pCwY1
46ePDsJvNh7rUhNZH6WO+AsJClwU01TgsZlmWJbiz3GUtQDwQXDZVD6B90n+RLxgIpWaSVVVbiPe
6FX1blpYcCic/gk/TT1Y+tL9ZEzBsXstmq6dMr/I6++UwjKP1toZsYKgss6CMEMvE1+qPx0Iqkwm
JSbAsTenpgEfY3Krdq0+KjYcQdyzON5wsbt+eZeJ+VL8IAmmVZA9M+hdKvOxWxx4LOQ8BhWcdPeV
0gPUyL+h186yRTWXZ12Xy8nxBm0q6VPMs6qvtsvCsYrAo+b/gplcJKHd7+9sbGxI9bhCyW44ZYjC
HybI6G5E+y+dkxTjx5Mvp4b9jIJNMaPmJn/NxzAHY9WBecyA91zpW0ywthA42DrN5T1VzPiwnDLW
qbRdjUBCDPxTBcYTH93B4Uakk7ZZC+eBZYLjvq9K/hHrStiFnS/HTOPLtlI03Bk7K50RJN1/XnE3
X+yphtbEYMnWIJfKnZkZ7gLFPN7csDyY1zMgnQCCgl4MGNysGskS4TU0Bk50PCi5fByMCBjlSDAO
xLELTDB1kCc8jzRpAjRVmIJhwh2yDYZ7+S/RBYAJ55YwTFURTJyDn0VNvnBV7SO2bp3Xpi3RtE5L
NGczBlJkdaSinqm/1lCchTkX7DwPYaQ1d682olK09yWUjlVJxySSrySgI6r2xQYtntD6t/oNxySu
tXRn2PfgkVCN6HDQXWHruIC/BpNDM+D/GurfvDo8DV8coBy2ulkBgGkimTIogRFuLny/jicBWTPc
cJ3DeA6xBGn5qbVWfuj15rIoBYZnUyKnfIevYZF8EEBLdm1hh5QznI+mNEnHkrIgcb11L2es1XtF
5rV0UB2J8z3AEI7cQH/LIVDtCi0iRfzwGXfIwCnS9z+HY6kj/X5mUsr4qpowGl/GVSab7CX3aQFh
HlYfpxeoYvjEzBQdkGyZcApOguv/LHlX62YBhBXEzQN2sPzmwl+u5d3E21vTxQ+Qb5qqh/pjfpKQ
MZJXc6bzdPZ5ak1pJuABGnkwN0r4gA7NEETWfRwOjlbib8vObeeHPkogoDlmII/dWZ8FdzLgJVyU
d3YY/76cxNe/Jy4BaABfOWzz1RgmJY+u+yeWUpbvSi9c2rEPHxPNK/GAEAzaeHp7C+MqthNqm/20
z4ol++YBXuod62/mIi0NsjyQbScL+RnM2S4Nm3BdU6MHQBh2HtF0inn3IA2+tkzsQLy4nKOh3JwH
Fyda0mbxJon/scBmGH2T3j8ILYE3pECV1urxEcxrIExsQBHLaEv9Vl//3JR7RbELgIg3dZv81P79
M76BSUyErrngGUYeWI4xEXQj4itRRVJpwZ8afCVqIcHGxeAEHKhwhdIGngcT8I0xpvdHb7WzQ+D7
eIVWg0pyiQUlAs2tCBYFskIv+1pHhz+bUPKFwftGR41CJsFoBmrp9YzjcbAoawpQJp/m+0DubOv9
kAx+f55d6MPBNWTLEwyK0YGGieSv2+B1qfyP+XIyEFNtKEIeI005YcPz4+QIxqjRRl9JANbM3wg9
XPEZEMcj4MU7J9n1lm9wvSxdIZlj7SrbBHLzRNgEzgJtAJMUMhE3Bbv5HeCTbfqcDGOHafqkJWhb
uNA+w7liDxCjeJVyHmKExIxf/kFIhE04IbHZDTTniCdbZaBE7Gj25fJbOSzQvMnmtJmkbJLvXg0j
XNSoQerLWwwJ9+8plaOy72JoJ2jNqh+98sl/QcH2DfdsHD3uOZampm7i/kZVan5aMF6LHOJJ9OjF
480pS8eQf5OK8sdvepiJYomml/jVaIshYAXMWi+8gcMmjvi3HxVCM8A9BG6Q2OcryZGUVXJkgasA
jAyrDFPefSSSkHN0vaqVd/2FMRWyVF7hCnMh2XT0kMEMHsoKWvs11h+/dHaqiszbxo0RLxIsblu2
Wv1BuB/QaU8IM7u8Oegry4nque9mrSlipg6FEtfT1kOD5x0m6TEiumxfvCuWG6T6fvCtBM854qui
4mzlaBOwlGgWw1epA8H2BUL/Y245XvurwNzWt7X27mU0rC7qVzjGxdW8Vq0cFvuh81HZeNnpKaTq
2gCAq84Fcz5d6KP7gKj5AV3nZ4/XrWgfD5OkY+NeDh54CXXFCEBFmH5/t3kf1F3mYg3KpJIKVFuW
CEG6kyFkZnaeNnrKSIXdDcvtu0tPMNvukvDXZeGq1pti+k9/xUYiu9JFOZC0rDB4nYxWNxLSdMMu
37nNSaTcxc4NJ0hNWuExT3n6rfgMzYek7e7aFjgE9afE3r83dDCa4o6xLNfSDShA0t6QXNYaPwh4
F8/pAvCvr6zSPbzKx1sObzRRA8bMiCM2SKlE+kd13sYkgr778CRt4BqiS/lyEwLTJLm8TDzNAhhz
22b0l8y1W9UOVKEGLggmWNHjUeQmfcYPQuEy39PRHoiT4XH9QBCjw+k91e5Uipg2SPnAZKfYwYiN
HOeOvMnP93nuXDwFN58Irg9XAZMqnuZtxK3v8eAl29l2J3XELZ2y1l60P3xTPLz6Ae43p9Ht+wk3
RVYRUdqIo0L3A9BiyA4JwGH0JqQ3McqgOlwD/YR9HJCIFoMtU8KYNlPvfsMVk6m/l2dh9/ScofhA
T0npRTPAcCwFhaH0fNDWDWyAWCeV46ZJ0g55nxFSGVjHIASNMFAdohdtq2YvLR1MN7kHnOiR6YvJ
yv35GLJQcikpbFTAttgOXymxmZqH5qzfynLyrPy1usGAWlMlsrxTDz8IirvumJ/8ATkqlPMTYPIK
Juz6M5XRVC7+X0bCgUPnhH7eRXkhO2U4pKFjNpTPY65vPtnqkulW7tbQb+hWRlyx4QMbgv3I1JCX
K01RymT6ayTVkj7T8maXlkgEGWbuzvLfQkFqo4rFLq19EQXesLyHRpJu3uDx1LBWM/ybJYauRo51
ZptU10lqzimND7vt3jyt+HSPm9jSyCVge9pHZHoPG4gTfBXK14mt+Nr1FQkfEXQ1MzYps8QHfdUE
P1HLT74dQHaX/oJbtEwCe4jaN7FLczpfbaCL85qXRS7TadY4eI92GwQy4EdaMSfWklBCBj+jklVr
n2luzGEQiFiocnlDtrs91SiKv94XsNbQici0NU6x+L4lJBSzp/mATP3bDSLypcAvqnGiA+Iv/ZwV
Tr/4FQt+7526S7k/O4OGxNvcMcR0GheUiJbOY3SINiNR5F690akLv5JxU1HW4iG0PK0pt92nW8SL
/KQD5vUwYdziMq1C7srguqPEAmq8TKiT5mZsSG6SIlqAPg4xav1OjXpxHXykl+JEiT8Tx96C3Kvi
8DVCXCzqnvDmoOHUEHBaEeS5JAhRxiHdLmhfVNcAsDKkHbRHxe9/1g2APn6q9Xm+wUYwPjFV90lO
0eB3xVa5nxs/ie7j2cxABLByUf2TBJBq+b5mvXvVN0+lU6LzmbkwR4dKe6YZ1d/vHNd6zrm3rwUk
ugsnUPkstutQnhbgbYmqB2I26yrefLGAttvQY/ToBr9qml88kwi0M/PbK1o+Q57YHyBZFLukj7Yx
BCcqWPe993TckpMGl50XUlv+8QMNWrVxHYVqjNRf2mD4BVC1E2REvSSLIGJg0EDLQuqRm0kTJ7ZR
bCuTPdbvcX9AhWcRzAtagt/eCWqEN3CIm+Zlz6EjRy0yHBxc5pe/XOV05LQPQ1PUeXRiXyI4b6vY
dJ/S70UWV4OvWf2BFInEGgnndumorSsoTJ2JFKSKlD7+dBR5rnUkMP7AY11GLPyyM6srGBUKr90s
/7UqufRaHQJfjxsPAvq9Z6TuA0sn6KNSW5uzCxC/kboRQGPPfKG7ZC1mzqwezFO3ATLMYa4T6tmD
GyfujZxgEbI4DnQ7jzogvtJen/zO/Ywrz+R4pVdDVxR6+y9eKwPDXsJC5cF6l2WxRhnBpi2I1hbx
8fdPSMA/QklrNEYRJ/crJWFQFZ+XHx8VyZC2Or9B413c/jjkKi4t3Btc0y4KoMbipksPUPsVreeY
gkQNtaydALsUhCaEFRsak5cjZioW3HCUhCKXCU7bqCzynV+tA1htGalgjPudusEiDv7Ty66VtY4i
WqL0BCgloniE9fPHkWfFwAJ8J/7iF9rctqDnEj5/iWcKMFoxENGlmcDjelGqPwaZfawvs4EATHHd
uVS5DfZfL7Z9RFZfvgIPUa1VmgCbR0eW5Em6vxxuOgzmsFiWpABWlF9V6TiN5NMdVPShUS0NyQA1
l+8mWgo7oh4IeZ3PjzKj8kgFJMCioYrgkeG9lqMF46yJEqM8qBVNwd6pfQ/B34W4ISGeyDSQ3B8Q
IIhZ3fLA2m0jSxlKvEFTRadElLPxXd7DePopgCj7wIp/UYYIdxeSHvdMR9jBWn4aoAe3JYukR/yX
HylmLi/YgS2fLRPqkAwKk8UXopiI4RJ/6GpGGmuzHEUvvHBnzSIIKEYREuk20USZuqmt79Zmlfy4
6XpxssvCq2BhrcLtXvTGPorChPzUo8OcjWr5GRnr/o3MvPLEacwHGZ+Nr2UgJaB7D1IOlu7ffwLZ
lwPAS4aT8ClyijJhGQdEqoPIloznth/ud5a5o7wcGlQkEVTodcGOdhyTwBbCfO29cfk47m8h8r5y
5FtA8uWr322qd/b+ZRtKqkY1Ws1K5PCeESD7FAQlf6CI59OrSGn1JM21RsM4nZIa5L07Sx38Nywe
jnGSuX0WNSY8UlarpdMoVQRb6JOLKIUeJfojENMJbNaVXuvaJ0vWr+vzgLlt//khLa12Ewn8MZuY
zcJpYOX+gfqxr0q/8ajFH8H+xRbR2vyJ8jezDkhLnQfmcQpgDnpnGGGLEokopTMoQfHRTQxzcM+n
YkkpHx9lHDcmVn6WKdaIDqv5hr3IzyRJZMIynAk8L9N9E6K5Z4xS8K39hBUscUi/OoUNh2wkoYFY
ENht3uWEjyx+wPfNoSZeyBVAw6t/7Hfr2PhFDUQ1zUayMvXQ59DHQ4+sVNYVAsb/kddil/WUQ4qZ
84FBFmky1yXCEPJWa7s/NoJtA9vX3zgmPL0PVDtrTjIv9dASSPnYf842yIj1pJ4E2dsI42GKXaM+
koaRZlt6ScaCbTo5KBG1fEhS2x8uto0leN4X8o7FG2J/Okkvd/+IcSsTYMO7NoRXgPbxYxI+gZPX
f11QUStBzoLGnMyz5TbT6Rbjqc2dGhX4SUsylC2sc6vvMywaXPUKbtQZEmQ6gr6zjxjRh7I35E+V
4308jk3J8sl2BUN8XhAEAbGME4ZH4iNLo+ifgzWIcnkdAd+oAfwHj1sQKncg2JHD00ZH0GBt5bj+
CNoyiIELa3G83StYPE0Sz5seq2JNNDfC7E3sihEay2RfqfuL4fB9CdnkAuG2IfbxOkcDimiDnZLM
9Pcf4juv503TxO60GqzU0ljyz4OsY8lYcMyFUxxH9tCRH5Xr3Bn5S26e6swKSubTG9a3M5/2HvTD
yPEATB5OafT/+7p5eg7yGNwACJFSStS4psWQ08jRglTuwxNCiukI58c7V5PM8pjj26UJpLsnXS9x
kwPzX1ugChLhlr+rc7vxFFTzHS8F6UpTF+cPEYy2bQjERUDD9IPGwTmIvsXD33UVWp4IZkjo4KvR
ST6isbekcEbXl60V+fCZTeHiihyaTW1BGkJKKHp0xMTWq6PP+J76stEeXRevFH2NgMnzB40s+Y6e
YzUd8jLUd16NnQ0hWElN+n4uERGFFQkU6YrpBuWEnwz+OI1pv2/XrfQmVi+/hOGyvDm8PocV9+a2
miCzc3hOTSAYcAW8ImFi2foIvh3pzyTjr5M++TqI1kbIe4m+ftqWEAwiFseW29ROGZcHv4+FR3qw
XSjNFyf3MJuq4hHdxNZSJcyf/gIv/wX5lPeLNnU1IJ8dpE+PDO384o1iSZDx8yM5aiSCmpUKhz3R
WLWsDWscuTcWWQnBhCdpeG1yZk5PVgHJ2i4X0uws9+5l6ETw420Sy0hueZ2Y+QNd6NnloBfG9ZHg
ottrxqxicbpWXSeyvqNlGcAf/WcpmkVh+SUpgdUUqa0Rr5r4tdNm+MLpBrMAT2nO9+4SnQQMyL/x
o3zOc53e60weaWVG7WPN11dIUWMF9iJRtJDgyuxO6n40c08bStom+GJevRmXi0PBF9cucYwCq+It
PeJu+G2Hz/vO7Ii1LJXrxolyGGxOi+OndOhrYICegTOj90N77A0MISjCOvKrSEKY3liAW9VB9C8W
BtBEB5PJCGBiCpIwThNM3+dk+U8wQuiv9Znb+Spo8tJD8g254ozlleAMDIlM4saC2vLN7W8QlDq1
eQw5Sd4M0/6cIJpnJm7/MfBt2b4WJudiuiImjzQOQgSIX7LgKcvVFf5iaKNTdB5c2iWqDFRYbgu8
ohVjOFsxuizZyrUv7IES36GSJIfOh98ecMU7/8MiBdqBL/8+2vvW/hIPQT8Ndm+O9GznL4H1eMOI
zVaQtlkE/FKsdJLX+JojjrnRBM7A0dvhVEQE6uLkxN9dA41yzCRMpBGATsymytJbzC4TBsMM4lL0
RyroW6ZuXrTfB57kVLpsdPh1CyV4DC0woPRUloPJ6Iwbiim749ie891jymenuj8YsocXjz61UGU1
NCwsLiE82cIFHuz2q4kldMglciBZp6i5Dlv3a4FKxHGaSAY+Hc4KwFlNuZy0CMSCg/Tv99/Ms6Qi
7obsjrJkw2SFXL69iJpXNoY5FWx2OojLICp5TFuTnNPxKuvTfKhDyuAHrxMNjgxGS5MwSBVf94Ej
F7xk6BpIXEDaC691MGLo1z4LKHTgNMXECeD2lxc3HtMgXBxEDsyZISE6OTwy8s/3CLGtoY+PBzsy
96uXG36QkHADI0kxu8nBIBd+LA0U/WTNZWeDGQSaId8636MjBba9hHqB/qYNrSl0twaAo42PXgmW
HXrgxW69eDNkGW0CNrVi0OzasbZqVV91b3/gBRZ0z0qwgmWJ3/Yw/4cOzl+QCc383lSCYYdY3VtH
3aqD8oc8KDSyLpIMkBnlZM4MY/IsX93aNHFMbkjkzraQAYuO7ga7VKl5U02sHoP0QWql5q9gGx41
N0DZoRDkCwzggTAck6xJnGTM5B0jALwAFN4Z0dWCN/Ky3ZAUF06RHlwIWUH7wnxDwDxsaRtUmZTN
xL3f6M3m0O++LJG3tchaevXaED5aejnWosd4/e0EPkgq1Z6IfTddTCzIazrIqkDBUUHaQjZ/WL6k
HdrQmtqSsvEXl0NN6Dspf+tT8MxEt/Utdi3airKHlzydpH6u7NV+zd5AdSOiOuW9wVxCeY0ktrqP
Pn/j4bhoCzQOA50wTTPzi/uYq7PIe0NhzewRTwWei5AZCvqjRyaEhSYovYrDNmwWfo8UcjTknbvI
x+Lz3FU7HCwHCrgFVOX0sxWWdOWT95EY+apsMb033YjosopgtMQB4BUn1WHX0ssF3AjJ210uNddt
usH2VNpZDT+eFsH1l1/n3R0+2HP27udM6K2zzBWmXQa3F4gBKwKXU3P2BUEzVpjehc4bwP5EoQFa
+ngjsudJsW50+VicIxWt7FWbHEF0Jpvjqj/WGVt82S2dLiPhtCp/DEXEcxVDrduhqWckD2ap/Xt8
g0KHwYDvYTvcOk1shpapDZjpo1vtcYkm7Xga7EPyT3cgUS4ya4GxmEhLcoeI2mnOBxdhsyKRyl1c
4ZEeUl8QEB5FoQW10P8AFL4DV474RwJn04CtXaplkkqVgOHO/W+GWQM+ykdJfgVL9eD2qveMkmFw
IoT8ZpOSkJU7ExNQyr9zyfHFGRMvfgUTiCCZkph3ARR862gww8/N6cMkG/CD7FTADprRS8I877vn
nQo0sriIB2hlX1NsqPA8BY5S4SGfXAdJKGzc/I5zsMXJt2T7cbhhjYC4BBngUt5gRiVzwg/tpkJ8
XyzAqmq/u2hfoG2DeXecMbSPIVTuiV9/dj+9AsGvnx8TewsCUXcDMN7A4wC6Z6OlhYD7kKvB5p6l
syjEzda5Ajc69q9beBxMiws5Xeh13FmfZrn9m1qEgvsa982B36X60B3QUcPYJzMvK6BQvizWGtf0
1tgzoit2M50pRLyGbIuSL+dbFbK5nDW66OKtc6AfCzObxMSAbzVStN7escyBr0jK4fyz0Rj9vT91
QYzZMz1AXe8k9eBwlzeZXBloNeQrGyoBgT257xwD8H8imD7s9SCEUT1KC/mL//19nLg6Q16LBfSS
jfLsMmHROSpMWdQKhr5w0B+Y4xsm0mfwmaw7kzo1b2Y4FCeb52Ec/Vywsrk2gEyBOlrf7DIjZeaF
g/E1TCeOJYWPrKUoROiVTEpEntN/kJvr61OatRjZD/z2g8xb82XeidGbnbgVDivXQwg9wp4NjHDH
+FiJu2n/QR/l3rPLu1zBK7Q/xCkDV0EyRdEDTiD5m9K/36Ktho5B+CnAijJeFZa71HLMLAnX93PD
+78kgRIXQaHBQ18wQCoumXUOeA/IgTW3tXNbwcOZjdiTsccVC5IJQixpvrC+FP+05wYKjPGXWNuG
48Bs/Lso5zBIZoqxuebDPNujInKOtJha4MmvUGzYWPUplh2ZjFrBgp89nIWk3jvWROBIszCQddAb
fUWs49XBUK5YSFP7qQb1h/Ht6Uf0o6pl3p0/lnvHzzLRuBoMGb+syr+/NH2rIAZGE04AVaO0gm6S
OHWaHcF3j03RtPFe5PEmdvfCJYJ7mm1ZaRzSk+oaOTho7m44uqEgjlgwmRD6CuMrZLr7JUo5ny4e
ryiI9ppwi5BaDWDd3jJT7AOMNiCvI34tT4iyqHmQagH1I9z3+it6D57IJnLqSiVPX55l4fsLBX39
1hUAJe4MGbuoCnTLyKGxokbUq8kDIkjqe3NbNnRtYVGsWv2Wv4TKugqruNkwehcUhXPrYYbX0JRt
PrIwaeKX9eXHPbD6K+2nkMwUfaX0qfZE44BZ4OHFnW1uSL6jNv/bDTp9DvRZ4lmZFUy6uzUjC5iK
OEegbTXviWUkzfpqIGl3dAFV3lYLq2KpKV8ZmX+z/sFPwaIXBJITsj1CJ6CPoBYpfUL7G74uzev7
0zKkRSyEhwwNLlEAIJPvKNVMHMq1TW6jwEoapmf++IFzax+3XKRJgTD0GtixtVT7fn7je5GT39dp
N75iL6AzxRpd+IN4tiGbvNMH4gLhikAwCLwHJOCLLbSO8Bs1cxg26QIK6Nmm888/crVJVmdobbd3
Skp+i5NlZPWcZid4v4u1CDgqKRO80Rkb9mmJ69Jc5oF6u5yRbXg4OEJj7h7bqBoNJmFylS+ALZr6
BbJIvGNx/3iGUR2Pa/av1+NanG3i+PSiPV24q0mJN5VwrfIzd8VAcrQt5ZieE+VLYM271oRi5YQ1
qQ+aBNncfShxKZR+36G0WXpA2CgeO71iSq0Maub2zszzxpux0tdhpm10TPJADfvBEkIJu3nOHgRg
sMv5SghcH0fNKJAUVcZDkONiCALDXyUSi1TEfSdooX/PDN9zmPpic5RjyFTwur2ASIuktp3hdlSl
RZbpg0d/IhCuEdr2bIlROL/MWN6DG35jQfR0YuxAgETXbGZNEdnH6pBSD8AbvOFQ/g65FSTJ3WI4
+QXUQFYU7+eUt1u+YTFn7zShzxBIdR+fEN7Zlfn1xW++al3f/QFFbrUhH02OcZ352XaL1ZUi8zGo
5++vSxmsqZ7TciY1uTxUu+WPvl2t8b9RIUXP6nxAcC2mHdgVK3Ekq0ltkmO4sEWDjYvxN3sf9ngC
2KPmzbhPl4EnJQDG/sjubBs7mnNAHXtAF5G8W0/Kt4ollRTYheyQbZXFE58zs4iJ3iOzy7QjGOpr
mJoa6X5svJ1Qn2WicYHTZ9ZXxQTrXXHwop/yHPnxMdMA4brd+VHf3kDoCsf+pAS1h1PIigCxHv58
6ruS8Dl5E4epLZOAtnvIE4vTEe9/MHZ87IGxJ5Q4P9KpbF3YPOJ03gLxu5TTz/9BrpRKtF1h6Win
ImOr0DcJUUcQw7L5IaWkuxMCEZto6tj5xTwq4oq+ltGHjd+YDL0udPTbz2Z/xtnZpRd/YNiLckkJ
rQx3ZCrSesvoLk4GCOFFImR3Isb7VPP/Ojdakppt4sQPdh2CIyaf1ZMe11Q50a1kmefQFwMwPwQL
8OZDGYBeVp+zt2skk9I/O6H7EXcvdcs+k3SU3eQTuGjTi4x+5q5UTEw+wgh2+9obfCOLgs+ineaA
YlItQq5aZDu9+Jyw36r/zUOtrAxt2RARsXJwdzm6ArOx26Xtx4oOU+W6UFcVwAaveCsgfQs6tpfb
WzheofZ6j/VGyGJkBNCKJGIhC6BQo6rpXkve2lgWabFGXNdj7D7tqsVwuoFQ6B7Cegm/uIac2g1m
aOK4GnFrnBPSg7030JmlCFYzNMypUOmoV+bMjfrSw22tFR+x8OAkl5Bm19oeyDWYLC+ePAJOzASP
DmSn3SH8IfIHjHSz+h2DAmtSNzB0khG4Eb4LwuVjgEcRmEyiTInfl9wSUWNor1i0OkknMqlbTH7E
QKgAADaon3mKyVA3nbSqbCQTGAUfeOPBPlEGsu8wkeSJQVhy2uOlcl9l5BM8N0WIOddX2tjKQ07v
0+CBYhn1jzn6xPkGeuPZE0HVVogk0wlcmOSdX8lZOu5b+UyfvxWnIrzWJFjHeAyh3DuS7pFM40F9
aurdHroasFk3Xg5gKZgmrj1BAnuVwNOwHJX1G2ekNF2CTIMmLBifKe3Pk3tC+HajMNW3Tvf6Fs+q
Zc083tlX0jftcWWi70Ef0qKwpoCgTmStdPh1wXUeikxf5P2wSeAhSNHzkAswNRRl25hF34Wjgra9
a45S+EhNPBze8VfbT2JoOXeARMDD2WAgMTAtk1VAU4MXLBxS7ZbqxF7hjQS+VBkfZ+60X6ZgXqdu
O6syWmgtogfoUWggXMK0Q1Hytgj9WtksvnpdEim+FAXIjVzFq0JcgQkxhgtb3Lm8G+3pfpE3PGuJ
d/z4IGhj93aASvm2IP6IxHDkjg9pSQL3lE92DayVsgFPmWm8j24ocovALoOLuuah6P3kk4ioijjW
rOtqrX8onMF5xJ2Tx7+51YBLdu6HjvMOxVEdatZ3/4D++Hb0kzdTZQ0S0rx3dbJnznCMP7cNLFUY
w559KBpcdDnbsD8tJZGksCXto9zFhNFyEovu0SPPNww/V8pBvkiW9cN6wpk+V+WsbmoY1WiMBExE
jcg5Z3B2g0oSItZyJTsfCnuGNkoElzrPr8YDA/8DbElkxU7BAmPtG4Fsgt5P5AuzM+Nluae2vt4A
4uhE4L9vvyG0i0wtUqCdnyGf3p1iRqgVoUl8cvqk06QLZDuSRhiNW4y65dhewV4E1S64DQlD2i3x
RtcD1pCjOWr0wXdxz0KT+ZxRhv4AetdJkDlDsYd0BT1T84X3oA5cTCbu3ZdPRLBZ9G9VJnxag+dD
Sr43blbA/gHrc3UmU2kwYpsZyZfBbwcccaUZTEqfgi3l23fFFH2YcRhoZs51l+bkK69AvvFdV3fJ
OGP5g8oTIYaR6P/egNljD56DafREG9mEmbHZHwaulwGDJXNEes4dhuUvnzNaBwucdVFahiUD7k+5
5p8zJeKoM1kb1wMD4yqQrdKeOP04aH9Jf7p/SR7KEiEauGBS6htd/2oXJQi4q4v0xcNiTF2/2LgB
d5VmGcPRqtCGX17CRf+4oxlUCq170Mjpfdf93M6NAmxRcHnJCmUyUEWROXeCQZA0y+UnRdxpxtsl
V9th75Tt2mERD6tr20X5tWy4wfOqtikNtRJQG3AtEsnXmk4k1NNZQ4Gj+osw6C8XrBESq5etUYwp
7JexW35JsRFah6sfkLwYUOm6PTAqZjjHfo/JWHyA0Txrky17GkEDSs81hOtvS0OfK5gZZXLHStT5
BEeyqP7upv1kg3svnh+pH+AVqfWpPWazXU+l6pHqokRaQSlffVxfm2ACIeV1QAzdeL5Ge1P4Hy3L
xjjokyIY8qVIt4ieuG7xZBnj5um7FkrfbRXQ/OHjbU6ziC+sCML12lOPApRQWzalB9WrIOVC4OOc
c2JWR3IvV/4xNUxsZpX6XNH+cVNuFIVNkEg+kM8c+gzWsStC+chEiUK4DYxvYXLHT2qOyGiuF1tv
QMi1hzJatVT5Ypfq9Y/MCh/Oq3U+BDBNkb1IW2EC/KYXLI1XzqmTkpp433hUDC5eTblw0IkMnzel
t/xtw84Vgq+S0NqrIPcrla2Rf1oBZBKLahEuVUfYwXd8PwertCsOa3v6t4rsaCZISzj63cBvMay7
rPSkb5FCQTrr9IkGBoCT6/xSmEIBizqLHXdx9YKQibu/128mKMZpqOO1QatjtUj1yjAkIue7Lvfj
jqSl9VV9EnqQuBgmmtxUEk/5L9yK1d94tchitOyoeBb9OFrEgna2qKyadUFxYEODp8j+K5M6x+vu
w3Cv9GhZcziHuRVLMvksq5zFCbU8b6eH86/bleG2qE9bgvg6St0gEnQZ+/jSv6Se4kSPsUNUExKO
iwbOjKRxBu92YzA4xYhRu7Yn6VlVjT02H+gISBBx7z6Nc1p3Rg2+rdmRYCJ3hQNgl2yt/a1jIUUP
9PisdNwcZhhQz6qmLjwD59QY1ie7TMS8M5CJycs/nscigtRouAG0kLvlmSRLtY5yKp1ruaUQaIZI
5LL9toGLKZoCgfgnXUrWecb7rK6FsbwVw6CSQ5CbEfn2tTKAuvK8Pi2YcVt/Q1coYCllZ7ChMmgP
5eCpKXJqWm8H2m9ppvmVDmMEkOhau0Gn+/f20jnEb0D2G4CGJwrQjqgDyMI8JvPBGp1CP6/5xdFL
+/6e2D7GwwIdwBS7hSeQ5QKGC1xLjHyOgU0TopA0+XISOlBQlBqkrk5zqf46o3irlW5cJ4sueVkw
SrbsIU6R6Y3G6umK7VUC4bTW8rglIzRRKWri1RX+Y83rB8wBcYt9TZuTnw4s2+y4ejF8nti2FZqt
ps/+BrYSUlK5IdwNeuO8v1IOCiqqes+v6HzJsUD9CUd4ChvPhIiuLUsi+0SNA2r1JD58zNrFMsV+
u7sJHhCEoovMO7d1/pE/GpUgaUz4eU46Uxh/kObXvujLE1qmOooZCjLX0ismAWgSTv+ZPP/MZ1jI
V+cesdd+gELM9BSXLxjOPKILRW0mwWn0+rO13OfBDufO171tLWd1/J9oEv8gkKZNQJrf9UqDjAnv
uoit+n5jaQAw1rrrIeGza/HelQybtSWxGHfQYfgdpwujjEYNLjbDZkSqamTG0AemwvxeiQn9RY1b
WE6jo36r11vCAduoKRwd408n13u6umV6Y9qwZh9faBiT2lIqIKvZS4nDsJEHvO1T/nE6N6QjBao2
1CkuyGrHBSnrZpZ2wKDfjQD4GrH4oEAG7tDKpHtlDzahgu5un5YycbLgjsFdEt9uS0C4ts0lVx18
LFmWBTxdoj/8urQxJw9SV45sblJn58em9ER0IOZhJ6Zu1GWRWFLecj1zFPak5+OQ6FRmrSjbWoBh
MfTZwQF4BF/FYp1XA1mpjFU/9I07llBcIIVoRYRa5fDhS4L1AXFVWclbb0e9lsJyaICZeDo+JNhh
WZNGwFNb3pa9Lss7HFsd/dpg5U1ao+dH3ZtHSR/SnBxcLPHGSY7BsDVREozFQ7XVTh+UiCoPoP+v
+XjyvNBaXdrzRAJpc43nEoCa5/ACNKcv5dBPB4QpUg+CrlhpdSGMMLrI4GomDvnLAGgvtOuyqRWK
8hp/RxgHX42KXBJnFsFuJuRYIPDUDXrVxqKQ+C0W13dqI2FmB5rbkkj3YlxRk176HYhqvwzid8kE
ukEowRH2rVwWi18y3CFRmEFodVd7A9bOowPmrI3l1Jn7ePibFxTbD7ppzbx7iQQivx7U2Qy5PqXy
vd4OxsaKeFkLW3n3IvWaLFgMr7H3uJPD6diCwitX01UhWjXlh7wSQOrUFVf8F9gdUzlIctcIN4iw
QmlyjA5ZnQUnZqQA9qNAeAP0Rqeoqs8oGRS0DuDH//cy6Meeq9w1jb/18Mz429OtKOJ8XGFuXAnY
lGK3ociFWTmxj+Inyl3mVMgDD2Q/5lIXa6m9rPciirs6sMMs49BmiRGwM16uKCyc0LLjkuzschSa
CpTTO/hrhqbIPDBnD2nijXqOs0ZUK3snDCdBmmoYQp8dY4wDRD+LRH2wQQylGhI5BlUMW8Hr8hyB
2Mb6wHSUoF2WDRd3gZPUKF4A0prb2pz1xP86+aZMdVkIeWT4aaG224paK4/9WDnkkbwxQ6IlSxeY
iI0ltNjvp//ZJ/dVhMX1e22gwnXomK4gEwq+TQnr39ZxwDrYd5vA1GmF5gCQh1c0D9BDp7hPgw+T
ZGiiFJGGbantaaZzBmQjHrpQIfkiVMTGIBUfPvAeg0GE1R0Dg9TbwtRfR9syk9y3fpJO0R6ENbZc
wU630skFpzp+RnppOcmS89FrIOsxBAxQTXOf5ODKChLFo1oNHvcheArmHJHDrfVmsS53zkx9RinP
tW+c3D0y/U+LGMebHPiYm0NB9pxtVCafBupIILxweiFK0/UEdeZcBMZyfwkOtuCv2KxUN/yDZAyI
spsp9fZdDZzzHkvvMB535C4Xk+8GObOoObcMW2ZFvhX7Q+ESxZ3+nPEilyFnGgsM/y4OCgIPT7ZL
pMWGA81t3xwvC7w41d+E2AuxZjysDySPrBT3QuXoTjW4Cg4yAh4xtzay7rJEmnwKHFL0fpzZ4vG7
/fBOU9vbwi+xczX84tsiL2Z3YXgo654QF9gifH0cDtc+CfUeIb4/T8uoqtQ5q9O3hu+qGSh4J2Pw
knsBfvxpuOwK0oiCY7hLZ7s61tSBm6HgMd4hx37sqD65zhV+N05BssPimGLh7xykCg7cMw/lJXw4
RctZbp43Jp7a0PnzISizWNJIF4eWDqUC8A7VO71QMT0bmNTDPhAgyqn+faBEjKKKloNdzcgdCWHE
74luwR9UfboDGxdYflehJ+rO31itz+Lnpw4ICH6H2VI5TnBGhaMeiCT6wNddia88LhYi2q3IAtsw
5eS2u4EkHB+xW9C2LFW1u4MAOk1Dj2KjXPc6Pqmay9lQkw9w8kme7r/1o7Xl9xvb5o+cZer26eFk
tSOjlu1+hQgijTDUDvJmPn9Qn+5QONyEToLT1dCYAI/2uAxcT8GEZiaFewkrtB+TiTqXfwy6Y1iZ
tsxWpztT0kzsBDey6WX0GJtk0Ugv1Mfhn+ISaIS2On9Z4/kG/flfVbT/lGQJGuAXFWe1EjJWH10t
8D0uVWhi34jNW923Iq+pfAdsaXP9IvwMsWQwh8NJhDkdVfCREMCXXUu0+FtuWhOMr/ctApa3l86u
X5szshHZWvWB6YJUDHlYsvOdm6a17aNT0hP7b5N0hOaKAMLXBiOTp72P+f1DKcgJwolDAGEu4O1o
HHiqYMXICysuQ12BhR+DF7yc08AOOFgTWYaVsztyxHl1vO+4mk6aXCZeX8NvAcKYRN4XHw8W2DYT
P0tJyvAPYjIhgAnheEMzzxz2cjCvKrKK7APO9i5BPAyrGxNc3gM1X0qx99NmJYSkCmjw2KkUV/Bq
BO32YUueMeXFio+qPK1Y1vuaDkhBk1gPg7+GLAzMmNAszKQWG9rWTUlWawiZEbwtyQ7bPE8WXVpQ
FTcPIp5HDuVFlniD501O6poApNbPE/UE4320Jir/aZQzaIzceiD4saIQkWMFRzcI7x7x1UExfgbG
bw6cMA8L6qbcKQRPrpl7CXWMdK8UCDNzOUKeE6JdC/qo68DQn+ymRE6fl7Cfi94nS6pUU0h+SxPf
4yl8dqutR/qvx3zIdRkZOCITxmtpJ4zV+eofpqMJG6TtqF/U0h/O+VWRv7UN9IkCMxd2yEqOLrb/
cQHBZRPo6LvZGruPVOdcfP9ODAW8YmOT8kfKFk2G7l+8JtvAYxRPRS7e4UyBxZo//EEcfzojKB3P
mOi2DEjLEnhecYJe9IJdKMZy8TZJ0UK+XF4dzVxuTf7kmhw4tVUcIjyqQTeFiO2yDIh+AliiOMlO
JGGcR0niaLTbAQsoNfjply0RD+cGzWzrCaBlp0vfVP3FUthhBBASPNw5H0mZ6OIinfbH2mB0Du8S
sh420z9ey4CIsfpk9Mk4Hah2ESzH+PXkNYz9DQaToxZUiCa/ISEfoxk6aviCGpTTqvk/JDyRyoxa
GrVjC0aW6CfpjVjaBwzzVvA+nvhTsOoeBKz3zDLQkWejk9DkJgMNTZ+4L1ICeYJdkD+qCkqWDNzf
3j7V7ljfOiqmkSMhACBELcjiOmFz1XVRna3rMbCYHWc2cVkYgx3Sd0RuugQi7KzLVgtyLioA2eP2
wdqDxkwZU48h2QlH0xSgned/vsJEkre50TXIsDfk/YSdl3y7NfyQB/FpURdDeeV7o50pmOT5FnMx
dMo0qih9AZEpUtrx8YQVUa20ilk2vglk2e3+SHYtAiIRWPkdDr/COvIuZLg5/SZmYkavQLa+uR9S
p/LBUulDxM9h2IOK+2fEqEueovRJWgv1seiZC9psJsbXxhTThw95uxbpfbUJOF3AvyUFhYZoPkL6
t2WVEe5RHET2/k9h5muR4aFpJffnao7M5MMIoRMqiQOzUmxH0KrohCP15XkS6cBeM2BIMVVitmnd
h3iZC8CXB2n5cAbpC6FfOU9uU2kjk5T+apZW133POOTCjH+zys6qJ9CDI0+7D2EJPo7QIHJHEKQx
AaZD7nWa2ACV2/Qm/staW5sS4Sz0tJfEyCbBgxENpTGsy4+ipqH+Tt9K3uad3veCRTylnigLtamK
62Xru0o2unfD4xhTxZB5xTy9PWOR1glK6saDrSQLMcQhb8gZDAFUy/HHwaUAU0+hnAQsCm+FSMAD
4NuDGSHfBDwnlGPsrDIBQkkY7P7szIsbNX1qfs1EbldPEJS4AiOJPBrBj4tLQuwOMzcP3hvEl2zY
D8KAeKLVRxTNeecGDMEwzVUrblwsMPptNdP/KJQ4fKawo6pA2yOXZIWr05xx6z70ptnRUqbKxi5P
+pLsanIP5ieZTSolRB3hhWDGX4V/m0UBN5CQHKm6sHqHX1l7NsvQxSs9RZJtnVBDYln4GoRYH3pK
J3/S1VXEisYDfjW+w+J7hEL96PB0TbhxtI+RevxlI8Yg4iyZLRxkcEvhZvxutWWRTBHxmqT9tqLG
ZujaNwCBwgCppZJRckeuk1KquVPu0S8EOOpAIi7nWWn3p0td5/j2FqMGK/BWQai4cwVAjOhtNnnY
E8yKNCLrVAteaztmPiblOkFZEHAXpSgnphAQK9FIZ8iFCVQpQ5Gb6/FLo26pRJbxH9c/h2jj3zoI
PjNuHWUbZS8BKW1CDMZN6MZg/iUwrCgl10jOIDUcglklJ6WgcVA4SJAEGAJLunfaXBombkKNgf3J
SxM8kCxgxhJeM7uoFl9jKTXEBhdE2ZSDlOyVQ0gKl5DylNeuqUnGDxHf5h57P3K7SNZu2xKtv/4L
NBxwSe5+4NR9yMDDPXIpDt1u9R+xpTIqirB4XIx9mM2DKfjeBd58N8+xgp5D2egxcMW0auxm6HcA
YtqP3jPNtAJp5zYv8lGnISK7KbALPe5pXmCK/X81ebzuvMSbNE8gpakdqb27+eNtnRa/rBIT01bQ
AZkzN7A0Q+3ZED3hv1auma4f3ZKHhdqZMGQrvSFBAeVY8L8W+kzbBoNUr2LnfXYW8Rx4/yxuEZ6/
ExP7VJRa/mMrlAGDRwSlAc0rrTsok5TLP867xPQxa5FexkR4JC067GThqU6yKJ4nwMI+GaoKPg35
Eaki2U3xyWTS9SOjXvh3hXndqbvCSComcpdgG+7IdY1ND5d4MzT4cR+oUcxqa1Nxh0c/jFSpHUH0
Vm8oviG8DE0I0REBtGHq6fX7Pg5uwVPgsGTYpr49LxmvwV2LO9nJ7i9ib/DvIz7DPGZ8t/amBXD0
/9bF1htBTinQSOBWXJfQ8SMxq5oOCDVBgkK6EdV9IiMbobTs7XkiRCcYCpZqwuggjRSMvQgxj/Hg
unJFE/AnTpkz73Ailkkoke9YlpnRxms89gZK0e61hAu9lFYmEm7yQQCNP80Uc/aPc5Noa2WPhDOj
08yx4rkOrcYFwYUjdnE1foQyQVQ/AOY2E7ktCbel5YnxPX2IGzfkWxiFYUVmFrirADJk73jxdyZZ
8xUFQahkcQOiMdEarB9QkfolS+de1QLnhbX03P4fQYh00b5Gc9t5/WYvEwUCUJCaSyUsh4P+q1c/
LvZwld1Uovorw2Qda/k/SVspWLvjXDBl+EozUowfx9NFgsblnmxn6Foy6lqFtXwxFQI8ZjQmX93h
Qh3AvvZuj0DFD0CWbo7GzfzWfOGekNZF8JZskAT04DhiD3VHjFUXS4B/ZUtVR+HKy7f0q2Fuxljx
GVcfcvgKEMu2haqDnIAyB9CXEU9ohLrAOMHn2JWtI2NDOUPTm5OGR+DcX2w21JmGaag1WieCtHDk
TsGLzr4q1Ki3wgE+1gwI8PKZdlc2170WRzwWePCvDab6tknQONeCXkQWvZKDAuSE8FBCGyAmcXNq
Ab/pdxIFcnI2rUWF2/dX/as8iKhYt8HHmrGWjL2ZX9+RdOOZmsFF/lObdDKmiAEvp7r0N5cJLPMo
T/KPi79yKwlvlCmTdSUg/F7+TtjMv4Q9XlbRsc+wKRwpVUKyD7OhcXs3hMLsvas09wSYIAn+5Jwm
EoY0zx+bD9nbw0qQoNd0Wxl2lUB3hnKdSA457U8b+kD0K0RXBTbeWHuALX4AMx+HmtK92Xntpdvs
e/ZH64jkTUgYRjZ2JDl0MI0dVLH7E0wFr1h9FwGEPUr09+XCIY7cf562EtYxs0hNhQskT/RcaAWI
JesvnFakPkTCFzpcU7QgFv/yPmSsAhm1C7Uvaa+zXf8w3tAS8HmSgIPdDCERpmBW9+lIKmBqWqGG
6VryrMJZjv46Ds+Q9nAoC2h7umTjtcuNxfH4i0VN1VJAWOvKk9/4I217aqKRNKEi3yrBhhruYkfT
JOWoF3jgt+Zr6hTutcs8sZjakN+lL97Yr8u/yjCynxLp92sptvLpQIIK4ySHGKqxTLDM6ulo49qS
SKSSX4/jF+C4J4WV/kh8AXseVYKKOAMI7MFImYmoed+VXFvS+aFc75PtenXpqNPqny5lbxIQuvsA
kl2pbncUt6rfaL0HHiMEVatXp3Qd42DdlEJVf05cUTj5mhc6gZidSFuTxttKHdjfAY2YaEAFhXOW
SekGzE+r/zlmic56YbkmQAVuKqNZVRZMB2Er+a2o0ySimsWud7enksUhyMmS91HCUth5zI2/rtNa
Bv25gfubNjNV4l/979MKGDfpZVI9fFnGj88weJn7NPh2UrC+Kk7++pok9N2MArXx9EFNs99UgWru
Dg7RNgH+7ZsC9l1F8rypJTwIrItAWM7jOgPUTv9Db1Pgh+zeJodnj8jGpfd5teE3NR/6Z//BzsMS
a+cdJ2G4vvuCbdatxq6DLqJHOW5WGOzheNH0ZbJMX9xyKXkiiJ97gyN8ISwxZQbW7LEdcqT14VD8
BQoQv5I4qlFeWCFhtBNCO8k3vVsV9D+HYYxfuNooYcogtFqdfc+XLioDOlg7UBKAhUxTMC7X++Ol
LH0DM/J+TNPvHc7QzQfEPRxPBp9+G3N6KoOjEINkarVm275tkIiUbjk63vbZunxNpSSR0REogXhI
YpVbicz7M3vRe4EbK5q/YiCc/lOFmIESRQf/Ojbw5+5DSd2LKepsavqoYOY3bDlw6bLue7Rek20x
4+jgo+ylQoSmjF5KTI/Litteyi/onUKIfBk8eQmSOOVhPeCqboK0dOTjDZ8EcuQ80UW52VoTObF/
cf0JHjnHjDVhMuZRRjweeSRgubh5bnzUvaf0TvXZd401Roz7tx/O3ipUVxfQEyiTi9cSBs/zjhV9
P6hnKIDGZkESpa+RAWNbNDRFNklJ8O0LCCZfLG+gV4Hytr4qV5ln83eTH0oB6j10MHGqhz7TaCEs
DUqoy82yduCNQGxYQp4+w0mQh4cnQpCXxEftsSLHXicITXF3bNb+IW8SykJB8FRJRMQgv+SXVKAr
cbHVVz9IWlv1ipb2XZxJy40sqlX/ZQgI/TXDE3fyNevdbijUwBdboZ5TPMDv21Wejax0uHjAKs0+
OFiUBp+uTtLx5RgZsBJ04GT1s5VUM4ZGGAqQ+LPnQiSWeSkkaik2m4gdGh4hjvfEICb93Ali1VsG
/CHydqkePjHXQBI3T+lWI7b70XZCFiiiW48+ZFBQpoG0fNNjYjfLewSzZifEcF4Eoeho+2hsUw+w
bWWQEXzyUqjzjMFqj/cHuOWkotQv1v5Ihe2uVCKWXesCvtJwDWXtvekG3fm9IRlN1yLUnzi6x6Ft
Zrk/EWc2VmNeO7UP4HlUke695hkclavGBqsbYa/q0dgLhQ2VlPEAGcqqKTSHdJAkloiqd/v4CbTB
4oruonCEtZh3nFHVf9sJ0XjVO+zRvlwuZOCr0aTQyMxiEJlofuGXA+/JuwyhdchuaeW3IaQRZfS7
rsf1iuPKKfbKVFdwpDffvEhNhEGQrHfApDHod8O/mSjIMogwvWMp6/LRQBmb5upUENUWSBqx2SJg
DMvxPuklBLL+xr1BOrZhe24qWcu8W+IUeh/AgMQ4F1A5cbqNlWn3lM+uRxVDIbXuIakjpY1/icCQ
XDJv/PDioW7pannKrTyF3xjqMCOG3VmLWU/lSxQKeuZADOYo5ID5gTAxF3L2RiqWtMenTnwhqODM
9L9VaZ3iIdyGQ0i0AgUZVDG0aI3i4HMHOHaQHItleCHc2NEGKLib1GPYZH04EDBM5vmZm9+J1xcT
O6zzQQyPzVqevhcncpGaerwz+uDjMtUI1YjZ7RiLBgw52o47v5vsrnUSFINL90PG2AJfW+nzGXF9
cngRdBeNyGOtrHTzdxHM1NxJMoiLlCyKJsoP5OALQvhg6U14/9rEzVEnNRbgSJsbfwpgZOlnkCzC
cPS3ABadUC2FOFw1scnQNa8rmPsxNVUApx4S40bo8/E9K5DXeb1L/KTWjrZ9YQi9yBv9Sb//Y2DM
kde/IagGlT7ja8/kSS+RteNjvuJLkkckKPmoRtmGGx3TesKNz0BnEUJodlF/XcEQFfbs8Ho6gd4L
PrA12JllAVKjc6Nu4KRqEqEl0BLMgX2UNM4r8/nVIvjRsbJkjiTIQykCuOXPwU+B+1YCnanZqt5I
ktOl19zPGye4c4cdc3+YeCtMSvgR177pYVj5KtE76LHyCLvmB2Hkw2glhRFnSXoDtjrpJMgBSu+H
109gnZ7yWB3ucdTBXjQRp/hfzez8F8+FHF5TdVc7lxdpGEKK4S9h7lXDNCC/g0wp+rcB+Qbt0kdt
tjX7MRRXCZB7WBoNbcleB1eWvtGotwNGIiEArdI8t8AvDyBHAn/TMiP0GEOlsM0jEYXjdKhjsFlb
d9NFzvz+p6z9oS85QUzswU4WsbzwRt32hk5/9Yohqh8ZQZn6DyFP49b5ZnmxD63UhP0GnWUey6TG
b00jKU/mEyQ8BV29aa1zB//b/YQyHf5ReVnzSIyKwHpHy80vqpKc5Vo/FYSeEqX29kE2YqsGtMX5
99MIVa0Xs2dn7rRScVF4/xmYlOHnhD/esCAsKqGwJ4XgCE4WfbM0M8LCx9vvSOQpOxDfVOEi1BHH
c8Myr0+GivJ37l1W+xZX3xMMHhYeg2w0/KMcvxFgc99kVYJnL9+gl8tbJZXI2kCC1bbp0VGQwQn2
xN6vsKVi+b26N7oyKnosOs9VZMU+UCQGo4AL9oC0bSeJLdHseHVORFK2YPKn23S1ZFnRQxJo9aTm
a5DKtx2avzG59yJMEDA405834FJ804bBVvGUvtVaTWY+1j+nuKmPTJVjCSXclqUDSv0tjuoFntGz
qLrSan4pez9eS+UNoi6ZV+Uqe9azBVfnYe1+Zczz+NtZ11jSa0Lr4IHeOQevVcsRuH/0eK99y6gT
svCmIRA85/2kKDy9LqI167jnq7Nbn6ESs+N0YH8ocoZPmlmrFhlX08+5aaJnGJXArOFvee4r6h//
Ffft7bzXplYCK+cbYhm4j4ELkrDAoWxrh3LB+G5fWmq5MfyV33S0fgYpkNMyrgrm7CghKKH+ahgu
OjPviL/PkdTsoiZTb1wY9p+7nuyMKTbbnNzmm+y/v+S2E+g474kixEPUjW76QiiHbNVblqTDe7fX
MLXu/cN3ASleAuxhXgGlWhSGjd1P56ip91DCISmUIJgaswFbgFlzP/0i27EL9L0lnaeQcRi1JVG9
IxaHThXRMEuoLtwzbqDhpf2/NqB0InX1tnfjbdKKnJNM6JTJ4vSu0XmbVaWrtj3pniEzIgA21/61
/+S8syDLOn285KUfHTo/9iNCnja/e1D19Ow8Bf74W5YDx0Dc3XOGYbCKN6TRbzDW+a5acbefqUep
/KFTIuFa7P70DB73viCc0ckayLvVqgcY0BOP/GzQfimw+JuJRIQBB3WqMwMvPi/CeMMBg5PtyH3J
ftEZ+wxMY262MKBEc1Gzw+A+efux65QgjnhHVlePvDZPXUqsuF/HcH5vRn7EydB+w9I5IrvbMQDn
5dtEctA6ErqalOMyziLsyBxDwljDh2OGUZqsJPuR+qlleE99vRHrk1qqdwIvDoZx/uYxekS0Cn9p
2Iabc+qITWz4zU1JK5axLmdAL6sIuHI8FtFfIRRkSFoDxRDiY1083zt4tpgMVTvUlFxwWo+IbS2v
fjEmrsM94He5VAWI+26BLUsHwZd9/REifMP5/CCjFgelYVgONCLsLwXTa7obH1A9BsXvAzK3CVDi
nNWw+4Ki4byZWvZv0mKoKpNYyyBEoZmvsclfZoOw8YERaVmT9r3Ar/Vs1OG9s8nMCA3wE2oo5qvM
71x14Nao10BtHXPgKDQRIzZys+eKPufkJKvNVqOtGCoxNT3ZE7BXWfEJgohLRjPikpaWTUSA91wc
miMmiE8MxESTJ2D0jpgkkkwaYqb6LoVAEhamg67peAT+8OX4FTu3GOGHfWgZWgh48wy05PTiCqkA
TFUasMFOj8bPRQDlJfgngmgsqpWf1WQhbH1eG6bGCX6q5+xH8kvcTZno0YvNRN+Ju6Ws4lBJdCLj
Yc0Bdfr3AKSJu7ezWuLMnwZKbZO/ju1JkZ5jhhB4Iy6WhHdRgqNe7j/wNXlnjiEDOHD/Hlj+NH7y
BQaIJbI8q8JPuvEoB9NEUB2kBZkshAK1Lj/V6roMNJ6pDBdcw81ZuVZfb/97efC+pU3KN0j3GZgB
F8kurfNalmDMZNA/F8LNCUSQmNCCTPGVaOzvDiqLr7KS2LCajJ+wHxG54rYcrSEltC2iVZQRradO
rHJHgd1M5oTGtDRGgxSH7KAD6FfajIB4gD/U5meTExXOWq4guv/vSK2BmDdC8bVwtVdELizG+8se
V/nkRwBUrfOcuHE3KzztZ/xqDFv3iR4JLLVS8KZ5WpeUh+4NoKl4wf1LE3SXB4zl3R7HruI7T+gE
TQaSEPRU7ySO5k51NNPTU8BT6/n4cd+hQt30rclTjH6xE/Z6a15fhXohVvP5vc79HW7LSt17GQ6j
ntGv0AupxssRq7QEy3dKKdJxlWqQ45nH2lU0nykUe0YxlWnjIuE2koNz5IB+PAm31PDaQG3CjF5Q
QoEVdTSor+6nzDtNmEV5pHVfYY5RVA8zqJZAXrkUbDW2Iqgl/+cVLO1Qp8FSag1vIEfid/wAsJ58
xezqiZQMKNtKYxhbF1StHzFHoBo1gfy2JGFXLnLiB5hGwtEPNhYLgrQ/NSdAHV/M2cnV3YqjDQ8v
53mLUDcaJ7Pnj1nce85ei6c0U7lijywaAap4NWPOvffiFn/B/5C8nmCJ/ct3mnPIRnGLJJtxvM7a
rVFwpk8ZjE6YEyC2UH5OxuepfULTMkih+c4SxUiEPjK929dh0WCS6EhfsXTe67l+i2qsGCwHMc03
u8vD5nVIw1gD7tp5j//UzjKTqH4oZywLYB7Be5I5KRK0BrKiQD1ZxgaTgtzvgdkjMG07pxbQnTF1
DKz3vQ3cq6fUwLlLIJBSsnFba2mlRkf9AZSK1NQbkcOb9aJs/1e5iMU7ukGrbHIo2CAAFNr+PiDv
qbDMXX5rbafFE37P8df2jW2I6nIABWY3vqplcdY1R68LGSmq7RQI35oqJ0fSrR0bFmfq+2AfCKyk
6W2icOhOqhyKBZYDCm/cVEUBLLtkbnGNHaFfiWE9MWlPHXsnqP97ZDanxCxHAaZ0rWPgyn20aEMA
R4fYiIGNp8triJoo0hJeftjlKIDKuwk4prlITqmDMhEIKIE/kLnKImg/bMR2IpggNnI7JvU0QvBO
ANWYD1wB0lSlWP6DT7tB9nkuuL2CFNvB7OXhZBLsjtACJ0JkrzOTmikD5QvCJJ/wGNrxx6V+vp+P
b4H5HlUP3yRDd7/ATrnzlIAfuEX4JvhrxMXzL6ylIBRGiOQoTyyumyzixfHggPD833D/2OaTqL3Q
EVfjKSm89RYKFJJGxF1jFrv826amCJlqfXO/upRxkzHwEWxF7eaYtzkqGKZM4lrpAuIc0MeEm4Lt
cviLJg6O8TaCUA2vD4Idcmhnhv4TeH/TCf4GEVhksgTwpQSw2ZBLfNTTnxLhPMMXHB57qV9tObX5
VOp1zjia2fNZXq3IA94HR0OoT+J7Y5iQQ0WU3PQTm2HMP1lZ7HG38+IbZi5PwC9wJ7r8ucIHm7kI
CW/wwNAowAmvmy0UXrRoHzi3AIdfLESP1ryILPFWMBFoLyz1MRbNngp6TdBRZBCWS61ZmK5+BGLf
oKd7xy/lmeN/CX1muBiQyy+bIw9QdR7/XYQLgKiHihWHzSS1H9t99Wne91ZmEbfb5x0j2Bk1+bbR
jssWcIqjBX9NRNxBhsaKe/fheIdczjSz8tuvg9ndZ17onLv1Gx5RGuagLIEwVQAkUohoWccwEyhG
AgKOrgy9M+fBq4002Ph8rG2nN3tbolkc+c0o2GrMgSRFaMuiPA/PW9GG9FLQtBv8XqfTbx6C+tfh
ytFMLh0JaG2698HJGM88XG6/cT3geVaK2kmbR45n3en40b38FurLqbqzBYEA+GA7d+RtL6PbpyR/
0vo6W1ZMBCD9WjuaVa5X2ssXCVCH/fM/AZAOshgbZl4GUTiIW8OkPI6Ksr35jZW2rOkyn1iddEB2
DBO5aWk9tCyRq3A2XvCJkl/0JJCN7S3K3IS+n9rpMPHvLj6PV21yXjQ7xmlUxhSOKXmLUsOrEmS/
/BplvD2pqgHEsEiaF3YSkRI0EYV6woFSflSqOTRJzy3QEVpSJeEcMJjxWHiXT90XxQcynj+oXCZq
fVMJ305xyHDalAV7GQrllmOySFMeYMv6RgKDsEM6qyngVpCSnJr5CSsjHoZaaMHebSCwgUDLfZPh
1W7CJtLsk0bQzq8jKnejqpRs7+9UF4Adkzrp6tKsk8X/sYaolh7GWOrwIOcfyvzGVZHpI3DrJOqT
uFBWgi8Ak4AyHbFg0bgmjC71BVp4dhLu8Vy1SWb8QvVlLbITmIxoGE/tTh8D/8o3Ex436XDSPHr7
4liMYvRpN9/X0GmYfWE+fe/UEy6cMuop9PgY4vjiLxajfu+V1742Fky5gGO9lr/QL7V3fAhTXGF5
b05j/9SPw1VCIcFSpKwqGOtu6ZepWGuL/ZwrvMSt89JiXwZp8134P4S0h5FIejcEocsJn+iv3eEk
bCgy7F9VcsxmdlpiBJ7vNxWAdfmatJcF4tt+Gz9TKrBcffwHnWhr5kgHWzt9gzl4oPTBIyw+T/HT
aPkWHVM/XiLJ5flg4QlaPHD9OQbfnG8lLQ7/TRpO/02KyjsdmcH7k4MuP3bcEdybfI7o2LXISibK
stoFi93BN6SavpPlg7cpsOgXT/uhb43xErNVo917wg+tYOZP38Jhawgq5dfdoLWFPV35uAg2XovP
e0kZMD/llOUM1tHPCdmdD+QELIRJQZg02vmG5vGwIpCRyvC4Bl7ri6IzqCxXvi/YJ8cVwvxbYy5/
wMQOIKCg+Ht8jVOKxaWmdK3/Dzf+GFJk+sNE+tFS46jeFCzna91XFgQB+4Evx2SLICELTSaPF5Vq
rOQ2Jgtyr6DfRHD5dqrXFau2YVgETG3433MI6Hi1zxN98gvxAPkbtplBNqDgppjXeQQLYM19F4Jn
oDFBWGxuKuDDfVed+M1HvRDJcOIapYoQszACQS1cGURG+ESsvgWhGngips5iB83F+ywLzyoW0OzA
ajh31Auv0EJmkVqCUFYlCtzaV5C6qiJ2DtptzyubmgPILQFXgdJtLIqpFB1WECts+cTiYN+Alnnn
iyCdCYLepQMBvNHVf45OhwOyUOnjP3vvS0x/xbWxbH39O8owpU9PXxvMM6UobNgyxIFVIOA+JuRT
klp837M+D4VHTw6+Mi5atChZkiakSYA4cckR/zvJMCOrL6Ekdwtxu8bb561x4ASoLOwanpvakt9q
xRB28JEYtQ8utspux5+UmbI5zNNVw5pCyLwSCP7pgxf6riy5kCi3G89u6ECUc38prKTbc7IK8SXM
xDjU/hv1Z5RKrj+lX/sARRUNd4BJohqgKcERcEJce/f7clxedtj3szIo9TVbyHA1jXOtfYoOfwdP
8Gi8euR1qNaGPqy4QAPb020o8ovyWxA5mxn4mgPwVumCN9LqAazJdVMl7yQwwXli058hzCFJ47Cq
jaJ2gJeXzrY/8wrmoMYfR9EMzRYTBh2zavVd+GdxE+oWj+GGlmsimAuQHKDpcOoTH7xmsLD5WRN7
hapl5hsSxAXJSmfi/sxlTwVh45nEPnJWOhDcyywDiJGQEJCOrpU9wbPpVBwzRzlb3N0vQEzNDDhV
evysp1P+3bg1ELl9E5DO5g/OaQ8DLwF3XER6UOrPV1DwLQ/5Szt1q+H/lsBVHCOSv0JUN3daPQbf
YiwlqNwbbB1oqQcuoXzYQQWTp0MhZtVVaV8CWrM6bgHXwi5OtOXXrfa5jkJ+ODmFoUzQU70AKWhR
svgGPtrUCL5o49pJDyUXeDkJmzjo2K/viW5fCch/TX3CyJYml7hxNTXDpPBjog0A/F3ZDhB4PJpV
U9KYQusZcShj9Slj/Rde5ZXmWYX6nwMTKGsM+OaxKsWNDhHSMozXjCjQQqL/8MYVfQyRoauLnZoE
LX2ZMmEJZ1YD1XD10V5J8aVkr3YM/KdhTOGbjBeudTFo36iGUN20dkI/Xg1C5lU3Rxq9fRt8zLAf
b6UPTr2770tJsL+zL1riwWb8AKFQAq+kDIs+6FQQV7Wmz5bY4HKPGViNpCpVLFBW3ppHCOo3Snoa
1o1eud5pU4XHcA0CDpWgFZnxDkcjkjI2AE4UbSlMnF8KWFnQs1sZZdYqGtgPmMLXasibnGHYH42T
iyXseCuZwb4QekEcVBydrcRvWGJYeAd1N1Fx8cBRXZxLgZgOp/E5VYEhbRAeYqWZOz4jYQeR8bbl
VruT94wlD5Ml19XtOWipr1vi5HZLKau+gdaJte7gTyC2uKtfXP81sxDDwK0rlq2BG/h+0mX2HbB1
tVhyQdDSWyH+18dJsiLHMILYFB55qI4v4iJwPm1obpSNFtO10f1nkVRMPdrimOup9vDXxiNn/Cia
y5vNjgVBuTv++adUMFJ7ZZGsGGM3/x/VIZppB6Hq6CZBb0U5n+BcgG0D7j7oS9qYqwaKDW161ioW
gXD0oie3g66vfC2+2yox4WCnrhrCj55x+c6AEPV1MtgdsAPbgFJR6KeUTJLCiY1X5bIr1C/BYisF
2ldq3v5oUAvQQNAKJF8Ps9uia4IzJDJaQoYHNPbAaD8JHlwLIV0/R7KhiDbP7HDOB/hpZ42pl+IU
54ux84fk45KL/JqJMQRtehNS9cimEz3+0pfH0eRY9ZV4tS1eP0bJ8EoEpHuja5hsunmrXLkMe36m
anIaWoywrvnskR3ZPe7TNBFjI/y/UilRfXkStnmXQbKmkeN3TemKABKyOuP2hUWt6JL3d8GnXP35
0bLUwzbcDIosCPxzeBm5it9Fv16k+1YXZO3GH+UjNFch6VoNv6AC03NRudF/NFEAg3HOsxm9gM+I
jwY1aScE9YF9/2sbYn80U0J3jWLRw+i24ainam0UFKk2ObvD5BM72gFm8a2bZcs7eT509jJpAkx9
1PeCvsN9dIkwcpMgX7yt+4lAGIW6nDZ0sXcrmK6QdGxg0EWVTYU6LfYcoDblsQPegXPnjVfruzLS
FxEvyMSxWHhunJYUue0tOLz9Xo+KkZW0rKzHjirmeePqZdMajE8JuaO78PKlSY+8V1iA8DXCLwgU
BYEDNlOaVB/FYNOQ9xxdrgR8eqg1Mkj/xK0k1Wx5dhgIctRDvmcIRvfSItVyZ00vnM1bOXhWnhHu
9eM1+EJ7N0GAB9jjT91CtsuKB8QOFFD41Yhq5vpuBFQod6dkw2DmIEcvbkV20rDI5GwTQxqtEw11
JiiNAUCu+vwpIrwFgW8lNaSSCf065kA3Tlin1KTtUIIEsN+eAiqE70DGiTUIieK//XTC4v3lnqlo
9DpNDebsjf9mCqaciBdwWjHUSFGgG4wVvnIY72r9xNH6HtKj7BbtNxswkbPfY4rSQzZZm2feaFWs
iFSJ05kvWo+ask8SCm8Lq5uYUBVgyMtS5J0fZKMeyu80Auap12HE2+8fnttM1cTAL04ABjcItd3t
AeLj7PcctxufyMrw6roGotg5/EqE+QZ7hZ7OVudeyWOkDulR+VgE1a0OxlSA6pje4oa+0cJ2M3Mj
/OwLyjWsDH8WhbSc+hgqVHJ6YSH2gFe5X/KC+QvMiNeeOhytkhDe054Wxj797GQZnOaDyNoe7ULV
wIBhLT4eSLjdpQ0TohMhbhJysYcxJbPEMnXsSHInGS95GSsA5m6n9AX1wEiBUvcuNYJbeMvFPBmz
PP+6HLfkNqJ1KsZxkomMZPzYa3B7BMRASZX0Jbx9v86DIhTX9PX0fhVWmutrPSOZ6akgSzqWNHNh
1HLj22u5GnUI96zFInnvExJ1/nYNNlgEH7j9Mp4dMOCsO9Y4iar81xuk2F+PYIxjRG9VPFmAtXmM
vGz5Ha1uDwxJmcMOWR8KtwJFUOU2LVOexgawK2ykImAxREEEu267lYL4wK+hYkIEweZQdea7Mjf8
JxyuV68JyXrfTs0j2rJ2Mjez7z7igLHFB6wa5nKhrMApP7BPtDgDY/XR531aMCU3IQtVmQWBhPLk
l0dq7nfYCj4JG6+zy/6BFzQYRp2PMf9/WDRWO1ccYCrB9kdXeFVzMr8DYheE5fZ2UkWHmB40B2OV
lH4os4miETYJxkrgqEX2jC0v/tJcrsA4W/LZT2UKiyOrQaL/uaX93Bx5fKXjEQuHXMePVv6GnvNI
TabIO86EI1SbIOKYuVgg7PDhZTJ4Q6C8c3B9w8XB9I4n6thAhnLfGKiruOwJhab6qyBCo9L6cvw7
266KChaDzPX6WFYX9Psssvt3f4GW9bJKAZz5/7MXaZvHbzAe3MnXEBzlqquxKkpLyZpOv+g52W9x
n3Tk3oWRi8PycTjAXwxE57Nc3xIgxiwuRxKDau3MJyy+nt4SxzcfemgJrfXYHECTbjDaby2GxB30
wvSQHpzpS9k3qg8zV96TQvYrH9ZwSfI32LcixDLees/YfxYQW7GccHUgzuhwBbB0FjFRXhH0vn3A
ZTisyEYi+icEZxVt5c0q0EG1UX77ursnX0+QJU9ZQx7H8nOtRzfDx+LoqUOz5X6zEXav/DU/8+SP
669358QWyPqnELu63ZBI793bSMgpm/ho0LYMG/mPm3D0W0bEsfxKvV14Lrn0WIzR93vxZGrTcm6R
YtypZlIp+GjqbU/KYqZ+V0fkvqKbjb3ZL8TVuukc+fsIEP7fABX5NVGS3jnjudQ+SUw7uMDvXcEW
rt4twI0pyLCx7l2vKvl68b9dHPpRkRmJVlfhypwXkOQkBjGbKBvTnna1lZ/Am9eGdZjKqnk0bgw/
JShUnM4LM0jdZXmSdEMo7ZsvehNIqxN9L1iC3PGdduAfC2vtDSMgvsCd0rar1QYW5OxjP0aOXZYl
FyhYi/1JUsfqa1eF9H9uuU18viINWC7I+NRq6hfHmGuu2PeikTeBMlcRf1lOZUQxz+/OwziWJuhR
H3qqQWTQKdjZwdf0V9Ekdm4nOaHCD72MGgjfQR20CAzGq/lhyPyKG7i3UPjTTg3qECNncsbsEjC0
5EgkNiivqxNXzMjz5rJeyGYxFyN38qSIYHDXk2Xv398OTYYkTJYLnfJiaZIks9ZLsBkzAkRns9sS
4hmEmTa0cCSSRh5QZm1FGCpFfDmA73uGC0M+sS04edi7IjftZo0cR7Kd2jDnNDWoDCgtf1KzgwoQ
6u32oHGb33WafIF95Lub2KgmicK+boXWUI/i4IqoAKMQ7Gj0m/OyjukJu+o1rYKeDRJ832EZxsP3
hDlTS9V5oQznWq7mAVD8s0sinSC8Lrw15rlrxOLOzN6l1WemlO5jFoa9Vd7vQg8apZOKABupBKeg
YyilVa56traxR70GpV9bsaDGeQ6NMI5PokC7YWoMVXJBEcWtsPTOJmv5aPgyKcmfJDNAyt+lKN00
ue25IhItyJ3D5RMPoPzEnUZAca+T2OnbLQidygRhaAuaFHpmwAVFbvPjU3/kxaaf53CpzY9Fx7lY
o6G5d3TTXCGhbwDrfA7bhS56cV6dMawtINdoIz5l6QUkuX42y6btXcL7WaIUiAYpXArmF+Bp8/sc
Taj5LcrGvTwvQjSFxzVjV1oopVkwWaCpzEOQElxIsW8y+vAkxTMzKMInQyzSSaqE/3Rp/CGmaJ9u
36RMhZxsMLqGqRI5Q58X1y8KXn5jt6zLPgxBP7Yh53rahQP+lDvMg/V3G6O/UrohJEBU4YaTht5R
1R7axWuL0rHaH+lAsPb7Frtqs01Km9j4GmQzH5blNqi7g/lzun+sIjmIwqv7/4/9P3k+vM69XbUx
Pv0AT8amIc2TNcFZzOxE7ZU3fWmSFfeFvLMQh5LI43BcHrwq9YsEbcX6/DJgmqp5ThFfWzk88rQH
G3vvuPgr4ppCur2qfiTJva4d3RbR8oxmGkbMJ1tkDOFfy5+9rsraHy1h8XSCG3wxjAtRp9fGRd0Z
dT70Ps99hrT6JqijCxIyAzFgkD9BXt49yQbs8ofl24tvpm+6XAuJGfFhhZ9csaWwhWHfg8ES+4PJ
El+2CgrNbBlEKLpCC+scQsrw80Wg5++xPj99idXeWYpdNlHX1kk1cyspyRym+cGdcW2pV3AEdFJk
Z17wAeLPOfqsj3lp6BlaWBTnuQNTVtBN7WAi0KH27Kqi2N2/3Us+991hsmywA+rxcA84eY3DFRPA
nxX1ZtgNa78FuEYhaSXwWwhBrGzEOsZunQz1Fd5OZU9ejrzMOPhl4bogrLyZx0nCI91BEnVSPy4S
CGWkWVoyOt2KWn/q5MOmWHJP33pf+J8QrtyG/4i09kf9G9OMsnw4IYgUdZBUWZ82wwWZPvuouEkA
sfqP47Ef67dB/vko5Z5Sb4V7Or6oE0KS9HV3W6cj0iuGaC68wW549oC8n+2L2Rm4Bn2yajTxkiSp
3O+OSBAxwVtfiVROJzNWvvKSLrN57prUJHpKf+vY1LA8emrmdUIIMGnTJzwC42Itn+tn/1nVw/fw
PxxF0LJx+JfartbtAMy+7zcYtYyOud6vy3hhdQQeqQ91vmXIi/Wul+e5xnZo9F+cgGCY+bnHu7TU
cix/NpzuLNRl7XwRbWFgAbOG1eTpL9MZghNGedA2kdST5xfoxmFCYfWTeGFrz8Ziar9cmiCXjVNO
VAOq+1isEjikY52rHyxhsL8Z6xotPVBqGLB3uCIASvP/vTJOMou1/WcgGs8nUMIiqj11LjGtbf6O
KmxaDV+jmzgXtlL5gpf/bQ0pvlfrrevHqpdxSqLbuhmW30MkkoBJbC7Ew34y7UaLbt+lhofS1Mrz
zXHpLYgFSMo+ztprm6VjAOkn39yt+Xmkh6A0gT0bTQWD/GNJbEokhqhqVNMR24nbfSkZsnIMewt4
G090UiuSijHHDT8ZjNCAhjsffsFhTlFdPnsMfMfWk3fietYNCtkb5boYMBk4Se90Kd/jCsiicmcj
Je9m28Lnd+ktXwu0ewQmLhDxO1oDArIHyLUIaxxwqTggjwL7OxV25vDdCmoCAmxWc1qMhXMdHycf
OzvTg0o2fxSxIVHcjY/tJmf3kTFOzGJEeMXzej0k4rwrtft+1gh1Z+oDFTUdlsx5turh/TU1vWUo
cXTxoNSw14klRZpP5j0kUzLYioqXIB2kNd9/oploSpQ2DRYYdI8t82dWE74/ck2x5Ws4V1g/Vb+H
AlWqZ1v8NQClsoVr3Og1DBhcwdBFU4UWLqFNDhpRjkHv0ff9wx0kzhMBm1JDKA74pLhDJ8aTDApL
adtscYfQ13AKv9UDtIyFaKeoZNrIpqtN3CwHV04NgzF7/5qlBuBO6hd0djQXsXG24WVCe1cSe9RK
6D5F9r7y/fCgM8dBA5ehRzM1y3KaxRF8cyteRREfoJdg/mv76hS+ZFCUuVMSJQh8dEo+VGtB+sVX
8tY5pPlBfcyagRmLYhqch2Edwidedy7CNZWzYqBjnvQyz/jq6p8hQQ6ZYCazhCsT5Ty5VevBWglE
fs8XJVsAmEhX9jx3wDU2g5qVvZkvC5AlswpHtAewF//iOBKNcJyC1C16mAyNJMf0L81cui1KeJFK
ufVoSPgaIkK8/RQHKY2X//RD1oZg0hlcZDmub3AwcFH1FjZ/4B6hEgXTmj6G6lSRGUkcdLcl9ZTz
xn40IwW2FJ7sRgMzgaX8fyxyUkPVr2yuDteUTH9UvKqIxzevNebBMZLpuDM39FiPc6pH7j+kUfLg
gahzChheDdYuSEfdInoj6VKFTX8vkyiMQzFqg07eKp8bBJ19NMFLyVESl7RIf1jVdkPuzPGgSI8z
p+i0CVOTlpwUZ6hVPqPiHxrDI28qYX8161a+Hb26iHfv74SeriHLJKAkXJoOQ+zhL1cA8Fuite7m
6k19ghpY4ZoTvN3AcPglNT+3QjNSDdkBxYgaolElpSG5/RSvtNCW3++Uq3R9jQzROhrafDhevv6T
7ZF87MKZeeQGgCw/Nnup27mnK30uspPPj9s9nZzQJV8tRUcy6u2Cs3/iQLKpAhHhgflFxOeekPpj
Hzogphfm+7qkef2sUHmbnMzfv2ntnenWNKL7rh0mm7dG99+0R4MD9jPUoSF3Utw/dUsb7XpYsIZf
C7BPBYbSGF/YdRWPpOwAKGwddAxUOZyeOLXuxNyAhOevvxDr/OikAHvkqgodYLS4srmHyTpu9TEu
e3Ui6sDHF467u7A1uGeHhNiVaMHZdsuyxUaKQnjNToYO7El3BVRYmMFvzMwj5r4seIduZtc1kptW
1hkrRPHCztNsLet4pZypOs134FY435q77tCJxICYSgIeehNobPC/goXkXrCnW7CmFsa/8sRkmYDX
9RWMIQcOPfKWwwaJoL3sUqUnCPQZzXT+Mym4U0cJGcSg6LgSFVvl4vSmkem8CXVKE0SdCMQez89Z
EiMjCC7ghHpmW23MVwFWzJBQMn4H3Svh4UCi/q6gQlRMUFu9Unz2ynRnm/BVu+dqpX+3fSjslXQt
NOBQFF8tMBBCu8u0xi0LGZ0wGMNSMA08PTdFp2+w4+eGXCqNhyFBlk64rk3q6Q4UJWZALP4MMa/9
hM2FoPzCONg7G8dMpJ/XPkoR5iFJFpggJOGOB75yIiUuK8BB8R0yhIgJ/9z9aPTtKtenU3S0bxWD
ph5VypFwO8nim0966VrwrLfqpyDVzMrzXg5Q62mpPSN1FD381Lis2TIjYSCyL9lDcOKugUwn+kuf
AKZQVQWM3DkRiEsDDgWLfit1z1SRK3c+8+KyJLjjlWUSvPnlGwKDa9lBep5SyG6WI72J8UYYP8iO
FN9zLehzfBgBVnKpl/jZUiPpwmp3imkn2cQbTISLuS0sA0qfye9gFJRnj1L4v8nGBK6x0QSG1uNx
5HT1TskYUSDWHGir2k8EXmFQvacwcVpWwqtu5l9+r2foP5F3eOYfx5WOhAQgMnPuLGMCKxqiapCe
eKWIW2U7AVXgBZeyueu/iBzveFrq4RuapZjCTC8Z4oNRI8TReCe2LdmRIqFr0QbKgYRYmkzlmIwj
9OsZP1KiyFtCLtvkJCRxfxdRQoqTxBtyId65CaspdPTowcIKzm+xI+KM5de1Yc9jO4NMB+CsJmpN
/GjjMyVygl4gvNXBoY/exd1b5T5Q3k7ByAZIVGjdt7eiW6mOsWLpp+QZBhw5if6Ngp2qLpMuZsG7
9zLz8rye/sbicBKDhJz2LYQ+4qe1fcGBb4/pA0ZJdhmiqetuMX+5Ghgy+VmEfne5I9UA4TfHeL5V
nqCFio7cxnSiJtZEGcuzZD7KgnxQLYVzf5g+TmJDw0VI3MLrb5MWIajvyoUjvDF/x8t+ZgeBrinz
FXrWr19HxooOV2vZ3DrURk3oWkp8mUz3t9tKDX/UucBLis8usaGQgnoHdtmK0XnFrzU/ImtusnxD
//kziwEJTQNcyLtOj1gaa/fMuPa9WFcTRTGO6MGLv8FkzTNh8zGw6PbH6/ZYx9GIT8z6JqwrLT/R
plM+JJ4thdf0cJbpNJUT9w6STMMp4LoGu+pJuMQozx+gvSH2REAiKEGrYD+Fk1iatv37T1G1GK5K
dlivDQXFtOlFzSOZc6nNZaqfIHUvOzVRvU8DJB5N3XLbgOUszBIuLm+CkG2P5ul/dJ/JXdMpXaJQ
cdOjBn/glXK3T2Qte3NlBJ0e/TXTii5M1BuJo1KIovPtdoaef7+nac+IO2vIvLBPV+2q7zt6HAMU
YvIldLRlDYvrhLHR6QuHAhnJHtEHWfiOSHE7wYBAquyiCNzniEtwWZvvqACOuMiWXluuA7AABnl8
4yzMnOKyWbcIGVkaRBymEPilt0D+sBMpjCkWw04U1TIBbdyONhm5bUBWtCo1p5Rd4F6j0UoBcuyd
B7G3+xwd0kn/gG8Yd592PToubPxCjE0WKjjSocDc/Fy+kvZXUxuJWUNPpQz9rTRJtxkZEzUOqU1d
j0czqCKQZf1XftTKTZ0bdOKc4ZNRknLCxVde8ymF1VCHxTqVrzfR3TMfnPL7i0D4+Ci6rJkk5xuV
Of9+aS7VleaM6zwnrHjIhAUryBkkLTuRddxljkwGj+5oFkFCQGXY0AyBscXzZg8kBB5sQEJhj81o
ROr1eB7xSL/2beN0TYviZNPoUBd8xMTpMZzYUKjLUubXq3PomH6leP4Uem7snD5cvwXMRUNO4T8Z
ReZYs9tOql2A7xQCjetx1RL+Gzkt2pOFQbVgOC67QSe5jv9oMei70Bh5dRvL7k0Y7rfM+F0MTQcW
TiHBQMqG55Rqetup4JczlzBIqN9HMo/Rz8jJkJELgEANGyMgok5M3/N/hBb6wh5SOuGYz+nTnjEL
rwUvaneAg0ozsPt5GznM18IRJ/4RDFHpcb5QiKq42iS+l+A/abXRCuI6nrxkXFB7aRsju3apXnjW
6BYSgXI/En07+rZMOrtqpTkzzx/PdOwl3G+BCCWcXP16ZyHFm20bHzIOxO3ag929q98Px+mnKGYq
8kJBMyvabrv41zE3qi8lsiyoIjBDypUegEFO/c/2V09LKl571bqACuWfIj1YmfPolEMwZ4FhWN9w
iCLwyNR/qOxxr/iu/6f0yyCuvxQSnxnXCqSB1lCEyvNjOAAJWTp2omN5qFc56oDFYLyvB6gfE1t/
4oiO80h6bLepem/xQxYjritePPLxpRSrUYCG1Qzzks6qg5bcc6ytlO2naSfcsRKNSsPp5PcYYoxB
UP9Z17XPlWmrBEvEmHu/iwdTeiTUrxFB3kpzNIWsx/tsdyTohXYIFHvomiWfr0pLdim6qxCdcP0l
IyiEe5ZoddYOzVr4Ch+sndPj5sFbnKknDaF3QCutGXZ9++ZIHGqU1EzohQZZwIOuJxX6mAU+4VBZ
4EUfsy84dt1MKXUJsvArBDcm6bi4AUmOvjjVYtgkOV7Obd0yoduMXN4sUmevZqaxrZ0BmlXyqGcz
ACuzB/wCsVRL4JkmItedMhlGn8yI2DHrwuryv27YBz8irhipx4mAByiFj5quuLAm8XO8Zbp2kbsR
58wxggxUsHvUjZv1cDmYCHNkMT5lHHPJbgwgA2stVPoOxD23YYJeAUtc1FcYceONYkCLcKr7y/B5
47SsLXG0P5yq2W/FnWx9ukGpVraV+AEgQF2pW0ujKwrmlgSpgoT/fjdEnisE/c2rNNVjkNJNS1HW
aKvjzZ3c19fTg2GSwQpUOYtyIpkJfrgUWBkkDdZHGxZBrgiDx2iS43xTd7AaeSYQgA2KM/NaFQyA
r7GQAxkvsvIhRp4eI9gyzKIyC+UzIa07P3nC4MTslm4OkPBoF3n1TFQL44VcdV9VXsAXeMdCM/0o
q3pZ+JaYr3AzvZMYE6ZymK1Guijjrwa4nqeXThRsbt0rhqg9XPxV3+zHpXC7kmwHtRw7+WyQfGzw
ig5mIvdl4YKJWT0cM6mDXBmUze8oozlkg8LDstso/URnJbBQAs+CWEzixCYj6n+lN7U0QP3bNxoN
eAnW/HkoMl/dDBQBymxzNxS8N/zbC+j3lSpeH5memo3/XLZBGwNO3LrHvGWEipqr/m8VXTvhTtfF
TaOsZONmrla/ndblNFTL3jW4HSe14n5f1i6vsNoaTjkaycSqZit8wMQULifkz4Ekak2kSOD55VoW
WVuJoQdTO3PzpCGUWKWafPtmko8Ec1TWhulKfi4MIoTKgk0uCW3Q8H4hvlxEAadG5oOhow+JNT5+
YnlS10PXK//0AYW8m4HzCjQB5WIewmwEMyFcVOnXgfxsBHJAPEiCFI+IQueQNkIY4iw2G2yKklcQ
6Ri7beIWpMTfYaZAhchVxyR6dYg1BDlmMckNFqDhWEWdapog1ZSUQMR3kB+mE3YriBVwdBHeFlgb
bjait0tW+kVoHR+s3woSU9M3/cFTZupL61/yedWgL8yk/ugbppJMYrJHp4k7ZksyP5imegrZehV0
c0/YUsCU/qi8k9nOItecFFk5F26KRX/Md2X3X6Rp6ZVCM3uFIDwwItlkLhLFCfXN1t7SgFCFyYEu
x5G63yOmIL0AtoXxZjqfsoKGBuOfqXipeEkkf1rs14FyfTBYyfEQo2J+pGoMUgM1Dzb4yX3JHipG
mSequGhGqwMHP4StKp7C3TOi2q5nGD8MQ22eEkaZVtcI6pZj/LjPgT6LiRoYliUBUvSgmPD2Gu8z
/VfIH5uCtcJ4T15u6UR0c+F/8LRSToNllmMzLR+lp4fpy5ZB6oz+t/pjUa/e9EmYUO7Tmv9FYuCD
q6E+IMBpjsbdusOfobGxcaPiWMVHEBK96w6g81a/FRQC6ODbUPrSpKE46uziuwyz8qLyUoAFy8El
pDtFsbywtQQneJQ14pfNe7MY1M32pPTKYJ8Mwwl3FiuEY5k5GGkiHoARTjNpEnceQuYTTP3j2tHz
XB9JlTD8hDS71pAYj/jLLw6C1UMYjM7WW3NfbaZVN02J73khKd3NNZqFCZ2KbzYNxok6nGqP1IGA
9auVJPhXl74EkxhVshfW2H+WTqxTYJCCYql146/3QwhMefxrUi2CQqH5sBs77mDhL559i7p9DlIz
Upqk4n2SlovuVFzw9tp/l9kRzMwvvDLLAZApX+zOLnDhVxzc8HlyRTVmBsF20iFqCXiyTkmbKpuc
Wyu4MV6rti7GQnONfcAoJw1tqXfqpD3nWUYFQOPpy0RyeFK9PXbkD6lLStEFDQvoDeSoYLTUqexu
5wOBXe4WVC3NZmm+gQVcti6wYZGxxS5pCsLxW0X9E83da7PCGmtQXka9100KpB7jnpNDHrYPnF9j
nQHmtOMluUKaxpcDFwdpWlKsb+LXvD8UTWlRgQ1kWCA6lUSLH6/Rgn85N4j/0NX1fMntPXIk1OnX
ms32JR3nLW8r7H1blnkOkPX0R/YKPZYgHv759cZZqwYESh5EZ7tX/XYHJBjwlLy/stMOD5uFsgbG
0cseYkcuhgC8Fy/vghcxVvn1BcfV8yO9keMc0PYxwPF+opTe9jGgnP9WcYLgV9r14+r3djCvmjYu
+XZ/BASJb/9xrotNZzorvuQwK074RoMTtUaYoaa/v2RM8MIo4+h3f6IfTr0LjGXz46PEXKCxAfAG
EJ093Vn72Tm0BNUKa4ycKW4Jg0YOcnfYe2TIZiH10Bx7K6r9Ulc9VZ7JW1ZYSOt7uaAFJ0hwwp6h
lG5wontqALLTKKn0cG+HY6NVV0kqrELKWJSyLEbWTw0GSiCIyBCPpxUQr08iuodkzlu68c8l1k/9
WlCY/eX+scGSmbNPs9jhVnc7NagnClO56qA/NH7HFu3NgtG2h+qP3CD3UBEkYtVSER7voAbMVeJJ
CzpKn4yxOVf11K9GqvsAso15Eq978sO4fuKQ3La52VgLc+xB8kio+ni3OafCCQY21CpuLbzVi27X
P9EV9SsDoMl9BZiT21NMLO1rhOBv+HJguk8fFl/AkWlfb31G42rsT+eWqYWXcWwYy2rb2OSiEur9
jyYok8nmE2v7IEiX9iVvLmcorUum32TCV6VbaOVyWeWixQCG+YRkdmxOOpxJAU0jV0sV9Z09ZUwK
fPvc0CY6eynXhBb1SRm1G7jSudXgGZ3/Hxmo8sLIaPFy0KMEsX3jIlEQ0XQZvUABi8Yd0r6Cj/a5
aYwKoICOUV4D05M+nkvF6/YKhRj3DH68OqvlZFOHKh1XjpyW0ZjK1ugWSsl4+/PI8USA5oJ7mTdu
7q8RSh/LOzKMj4r87IBRv82Zdh5kE/iDzSiWnWmrEKplzdSqoCCSPj++k8lWcfvvJWJ75XLKN/It
Dzdtul1Au588NuE2gn9KDwJXm1RjAs1A7ORuYjr6NckTl7QoZgYWS7nlExrHqTuYujDKbW+96Mbf
Wk7AI3M/8C9DIdAH8L1NVpT9G1pnkQ4zcJaqto4NkoCTnkDWzmpD4j+exgY2V9DayXL1jaFllOS0
Ytkk9Lk4KE8Q3T4RbxaAf3ebo0MbrvXQXAPYZQSt89cDSdBac8uIOyu17Wg10Py2NerFfbWI74mD
yn6xa+N5l3BcwngNoaOdlHh6aUaal6GcE37u1i41Y4oT3k9TEsfyIuADCrO4zkk06utEJY5zc3St
T2dOzyxad1SeefMkC0i9XnBjR6t/n+5kHC9ukd1wuI1KXFoZtmuxsVHiQCkn1gl/5YIEiSqdR3nc
9iZVUs4O0McNXMyaq2hug/0SdvOmc02E/ukLsgGLQTkBinnH3pa3oN4jlCoOHRPUDZLe6RH32HdY
rOzDHp2pEiWmxhiLve2XN5xX/yKJc92Qr88T+VBNeVxW2LlARfLC7tN7fN38T0Tx/raMguymd4px
zKhLe+YuDjlxhmNk0f49XGf7qJA7z33JKc4zviGaxJBQ8HS4C+mVaDJdKuyHW4HgHd6m6j05Hg8A
dsgD2UOxwpCVmwHow/lxA0V0XHVygwKtaU7YUTXsRkLyRSGKWnXVrQE3m77a2vEUc2ZXuTQ3SyfF
OT9Zk/s79YjjMkWKJo+U5mZ0hG7PDK5/d1kKqdiZwofX5LErVRPQl8yo7d2R4PyvNakhz6YS4zOk
BxAgNOx1Q0YyHBOdW78gOdH6Zc1c+xpTqJyKZ0msBe9RQieKdoREnalQN5DIHH/+ReoaVnkZUCPN
zz48G7HV0kpCbrgIkt8RWtgkNaGpqkfqOB/7l48b5EDiFs6ksJlgFV88RXsVCLbbswFU8yqHj7o3
Gk/JVqOgRHFkCX1aUkUlmP0+qYPIVoxq+i8hNbKbFFX95SZDu1FCNaCDh0xWLsuaQvrm4FM8o91Z
kg0EQ9InbxANYhgdQmcLqUOvFTNA5Z6+p3gKyixN5HLPj6h0OagdeofaeLm3iwf3L7fvntf4bIZh
WntZVbGo4UtfBnMWs/QLBNZaodTi1s+8yuleIWzfZ2KSwhQU5gwRsWP5/QCPwiadzWFd5WbNdqIJ
vqTZ6Fak8ES8QROsjtyPVBUDaYnFl9PWULg6ULiDpfY8d29mXwwSSsrAicOTldfWeW44fI/M+U2C
pXQod6GWsKSFD4oZnmQP9aXVeeNAYqnI0kt7fNL445TOa6wNFWy0Ukiyv8gtY8RYt7pGOF0xNdCV
qrOKwbugkz+rvzdhOBNO4/sOqmyW9+15YWqL2nLRNz1y+CE4RvJLp5PfYOlvTt7NLSBkO85IL0DI
HpJfapM5bBnxVWz+a/0HtiIIm69e2LKQgnl+5iaxwKBtC/bllwD3bNvq5JfjIvUwIPFxvNrrsECS
92JX5qEPK7n6M5HbLsxfTsk9azjfBAQhal1L1SQ1+GPeOtm0s2TBTiOUSKjHp5l7VrH6Gs0opWpI
1by88EYBLIJNqVB7zOS89sbRNalZa7j50YRtBYOAjipXTAh5gRwdJFOv1O0SPPhKd03ms1uFHz1f
2yycyinoOvZTAunWWbTzhB1WfxqAoz921AADOL9+w5pC6E54yR0GtwY87Q9TZmMNo4XmQQRGiu/l
8CyQeTuVGayA9YmsFiGRYQmq9Lgjn+PIdmf3jIPZ62hA6IjwtMdzJDDlvuWeK6TA1XDExhths0Xl
Ho6NO9nshvHaxI1XwFprCFV9jUoN0kPmMRUNoYpxEC1v3tDrqDq+6aEmgEOFquMF7nmtqf6tI3lP
z2K+zaprjaIWiz8PomsdNstixj9X+oy3M+WjFFYd31h9FNJ+OD2cQCFuiWaDyDvcTvakS+gWnWrb
6nTg+IQXcehyB1Y1OlbvxF7We7suCx1/7m6MVQONFBeBXdZ8Iypl2kojtQmdmsMWDexzNZ6yHwfZ
RgL7ARhZ1VbgZrXkxA1K4K9RAqcKmREcExyC3mxyzXudesd0uengEwfP/cRJ28cyPbagduVvKHyB
/50oszyK4PrtNqZMBgL0//tVExGdl5OsCeyb6ANkipHkg+wrFfiUxGoUtChQrKQAqAx7AVqZGvZ1
f3PLG4K18um+3IHZBgG1dsszskuxhh91iKTXoX7I24Dj54XigTWE1mHwlakyDAK/O1ucIQfEjyew
8fwkPl7V8hweYOnOeZkybZxgonvnAkSxxB0GXucP24M32GgBTuJrQJ11H5huH/tLkYveQfR7VU56
ZHxh/K0wlLeWOuBjx8xMju/MTubfHsliL0qp1nGEtyUXjoOlSL0kp3HWCoHuhcfyXKnmAS0Nu+aO
TODXhatAUePeIj+4xhfuMtfA/pkFIaDGxYuJCgRI9HHYowOA0SNhqLWjhivYnRzMnBIkU2/tV+3+
1l84o2dhSYd4QocNKpaYc2ETXwMN5hYOHosLVDS0Ha8xpmzxQ1PuUbZXe9ZK1HV5Ae21QLsuG6gr
MnZTuWIj3pkG3k4TYl2YdvDeGGyGEEQwNhetMmhDYFC/fO+xm+ZAz+GrwtnIKVQuUJchTzubonHC
HFDrEuHNJWrHryxqy7PpmgNnkUMZTyTjpJF9G+60VkwrHr0f8ldcQnImR2+G/t4I+HVQtfzkp2w6
cOVmjDfJAaKmUOWYBRZJ0v+j2tEt+tSn0FjOMqJ6RkRY25VtEnTcV88/Pwr3iH7gUCOkL4pUjLFi
RMXTgezoF1XU901uq4oiRx0q7O/P4Go3TYmN2CcWCgdIG5o8P0Mu+83x3Iijkq5TOuNjZ/XakhRH
Foryw6OBBxJ227Z2m7z+aDEGZC4Ad9Rxuiiv+pyBMwD8yVu3j1e46dG4aQBGD2kfNlT8YbYaSCcs
DnzAXq7TDF5gpAsmwGmXJLWwcp2cD36m392Gx8PjWK4aNnYhtO/33/bTqM7ewyOKB2QPWbATOaHd
FrFzpfmwoc0O+Q9LiEEvIdOonyf++C+juBIYtnFrp/nEkEDTjCSmiHIxe23C2ql6JVe7TczP/9sF
6j4DCncRHTMGr8pLmliSno5aShVEa7Q/rm04mNimPV5MQxLdSOFXhWViTexLS1+jS568/UKOA4cB
lB8hiFt4y4wIT+6nuk+Sg3k9VrvNepUSPycWlzHyKYByxg26Md51JsO9rwH/QbCJj/z5KFm217AU
qA7aePECZEjVPidFmfw1hPCvrVNn3DtBjim2Z31biV+1WOZ4yk9QbdGg5zSAGnsrN/0E/HJDVIAs
Ii73CE4lmYiQ7294HO8D/v1LAhkxacE5X5mlXDnpljYbmpc1sbYwFsUuz4ICLntYXwPzeavI+A3B
xh7aUuvR887qZQefazwlC9PyUIzXlvZ7gmn+dGwjRx9jDKwCIZzWdn3d2sjiDwZ1rlWotAzCeZ8V
8t/nwiHdn1qi0XAtLdoLAreYb1a/vVZ5xUROX49crxFPyOsYRtaCmKUDCvU4m0TLPAFb7gQCqjn3
/0s1terjA8lgKEjZCnD8CpdXyP/GNUceDHFzWMaLcnxsHGXbDUn5lTTMkpKt/gDet6dHX4UefdvV
tZqjsKcgSRXVQA8Btjoc/2Xa9IPxsxbYrXqATyy8F1+wgt51Bos/D3SIkxRhQZWQF9Fyl46LFdKd
GBlqlZkCbQbMKV9oyNVOnwBZx1/Hvn+iqNLwaEJz7Pd71ys3HBmYBdgQHz7Or20HNxMRDr/UH6Zm
AiiCrF0g76HDF3eGJiqew3Qm3SpfvYPBQxZxhkVDbWPaKtiy87sYwAGfp0vxAotE/sV0YrtFdnxl
ZPlrZNK/VmFDCm9+7sEjPVce1USM4VQyMMlpMVlbspCaNj5STUduXYHtMsN1T0aU/vlgQY0X0yQL
rIRh3k5TDUNJwrS0FI66et7Ie95rYlRfSXzscYKc7wshJLiGICdHFPfQveKbdigDkcpHvmAELXxG
VWmC38/ZRNXxyos/iwTBuwq5NSjZczh0ATJj68h/KSTSX4+6iGrtVL4uDjRBirGGS3iokBtIcetp
0ahMXR8Q0czIX+3ISPHN90b70WWDlALuIW/aJ6PhY5y2Mqob7XuBdJH6un8VcDpowCBDobaYXsye
urxxMCnDEAezy5iIUk3gt0k8lfEfJsBI88HGi48qqSlPfHDyKYMnJIHnLW2JShk5+vW+wJZeIJzz
c8fOZsFYejIIEQaOW5QiQe7zlF0I0M7UpLVMeqlHBZAHb+UNrqhMwVbrW9pJcdhn9akEcJIKZQTn
5bG3jsi8j3R4S7+HBTL+qD9gvE2hSmI1yLdpDDxCkYC3xccz81DnhS/XdMDikDDQNl7qISxakS69
wEdgDJltsZHMvolj6fhjH884YIgkA6mCyCnCZUKL9h23pchKnk/q5kqAS/oSbmkkVwjoLry0LQhN
FeUzFB0ljfSiXQ4SAD3upuvNlMFOVNtw6Mvq3A0yf5HCAlS5kSk9bty86KfScBzteleaP4IvQ4Ow
EGYeiN4VgXNLVI2u1m6TlSh5052uCO/5yQXR/DlHqaw6L/3gGnHqfFi25D5afOUQXPa45M7wJAoH
k0GVD5JCzZJhWiY4y3u9kgZDQbWMX8UPQ0GnkpRd3/4TcdsB6BpsW0hdcT8CrsT4qO3s8MG5tzKD
4+bIa78AfT5PZl/Uh8ZYqYNM/Ldbaj20cdiO8RB+LgW4BIzWLKIAZBL6qg0kXNe8ycrLZttxWJ6y
AOTxVR/edR0DD6EFW4j77QXB5GH4T8O7AEtLEFLNI3wrAskITRIIhtEF/dYnqxMVt4Nq42fnE8QK
k16YEPxY+CrFW5c99xbgbpLRIJXCbENBWre6uhKGXDgrrIQO11AJoTWfH2X52WVb5+FLmpYaM0aU
rvX8VQKtPdV2lpRhC8O/ddhJ3EVrdkWSPrdogqX+nStCY6g6KL72vOhFvI0abfHogisPUZdBgY7A
IE3J9Oqi5r12ZuE8+leMTlTJRbBeB+oDxqT5A/HNNv6dazdDnIWzS9zjyb+khAie0yFOMB7R6f65
XhuuZbY1860c0WnvNyYHp8PXAToGELu3L6amgggfKEX8LcMCErTsCYtrn42oBBwvbAGbrPGXQ4Xe
sHtRxlSVd6QOePHH7LDASYDsp+tZhhOU8LQ9Ku/Jb0hPBR+ZVr/Qc1Etg1Ezd+Nvl0w2B+RfdGov
ZSwDfO1f3IZaZjvfuLC5WwZrJOGFshMdisDI4TdnxRpVQG1NiaK2yqmDUQtlz/MvHXQC31nEXqqh
cKck5Vw5IInRymA5/A4ZqxgpYdQE4a18RD+LMenAh6PUMz/XV0CeC9TMRlBPOU1jt2UDhHVh+8c4
s/AF3oFRoL+fX9qDhZcyM7Ke4LwmzVQLGEsGoY+k9yPAS7ofyUZNS2MyeRh0hAKewijNGmRuOEkv
BF8eYBFt86DsYL6/k907esGYEj6CSUiHlrfvj4mnoUiwmjbhaBwMgvHxMO76ADLVonZhd/v2HViY
O9/oe0auAvxtCDUopuCp4bFpXTnfIon6GPudRD1aWsC/fy0bs2vwVyirtiku6qX4NIVvKYqPJj2Y
ZFq6nx/GKxD8zYQln27aLsz78dyfvHrggTADf+QweowqDmhEkDAmL4kY2Uyg7VXpwHxKkHiu/ZTl
CyjOoZq/YJv4sniC4cjtp2HtZ3vQa1az5IqVT94Bxu1+tjRdp/txfX0raP99fretYF8uk84XAfyC
4j766wkzOa5FLnuJ9RKiIyo6vNJr5u/9DaewH+f83gYRhBwbp0lxsMbwKrbU76FxMNzJCcRfnXpP
IJ3fokEfDjvXWMesky7eruTfh1iK4aS6dHPLkCL1a00rMsS/b8KZT72HPbH2r7xH++4S6DO5qG9v
87hGq2IO56YsoSulO//hbtZWpSKP4VT1YHKQTyFdBVkLisQUlO8YvvlnSqhANDfNQRffUKyM2qan
hCncHZeofaMvynpRQWSKWnnJThdwRKThtFoiEaKqCAw7xhIpPoaRET0QmevoZe71M1Gvs+DX+dBm
VtFlE9jA10y4waDcVPaifCiA125kM9bgLtLp8V3smL3pvLuutKR6FpbubeQx9/UFrK/b8TVIvdxG
wnmJhlj93WdinEyv9vnYUJ5+2TE+DjBsFpR//03wRVVjyNencBtUb/qkYZKd0Rn9evKabsyCDkzw
VEv66IfUUYRg/JB8MQQgVBBLoP1nA/zkCZeDmlIzUyDDKdwqrJanx16JJrDVtclvKRuNUL+fQ/+T
QUh3A263Wukbssvmlv4Hq4ESjjfAO1a/sLJMWhGIHAak4mIkKHLxZb9QCgjUozFmTjD3KPyOR7WH
/bGKy2NB3G4OM88vkMAeuWGU06mScUZWx5a1fulM5jgUVCz0tGBC1EfWHsc0AjsSE7FNzPB5g0jR
V3XOl05Yw1WFP7oQUER9Z601zcEhAiBjxvc94CTe9qU3beIwBVpwTZ+K7IR0dLKIvtWLunRpSATo
uGAfcBb5tLWCLlAZvGQqxHtg6xMj86nL3W1HcNX4FnGhl55OkMSWiLQeC0ro2Ll+s3v6eOEnjFnF
FEV5XtR43danMZMsQ4ZzK0EdG6bQt6XTvrKtkW2eZuC3RolT980TBW4Z0MptSXsKzBQgdC+pNcxe
prP0OHNG3jiO2m9Aqtw0VRCEmKZ1csmpXROGFWYFz5S0iiiFbHi/Hepfd9R2mRSYNtaqnXpwSun2
s3f7vvhGdloFcP/S057jzDFWk6b8PDkRgkbNcTJ6iT5ek94wDU3/lRiCvB5aZXu23ehJsVuvoUVw
q1tQvQywVfW1MFT+RohlTn9YFwdh85yuyruRUNOMQWoViUSrWfyE0SZ5Cv3Vtd1Fh7w3vPzHRB99
CBhsm359vWQKhh+x+QkcGHn4fG27ztXjqE5B/+X9ZDh8cVjaXDIDjKcB3KlrL8ugMiVs0xQtcJ3v
RpfeDCTDltyig1FmllFUXXqtM7sNq/ZVGZAGsG2kichiAiRXvJkR0bSL/+K0GuXeANaJKSvxuwHK
nTK9lEEWv08LnBuzZzLnIOUX+yg/FEVZLGz4XWMxzEirKTRCaNwvEAkKkqRHWmSzzV57/q/cTjTL
eEoe7b97ZkskyzetTL9toU0vSVXXpStFraMUFvgi/J/UHUEybbueIjb7XsYwkLk0qCNMIteZ9fFb
dchAcmwGhHGht0eKQymBe2duGE8BjiVIVD2DIvO18swAdJntfWANjyCMrng9QLARatwiSE0O/1f2
x242iuBxOI71vvMmVnG4k5YE6UHQYFPiLO0G/P4jGs0X7e9fhfDhfaiihkngfnZScBZo6eiA+A47
mBQub1W2iYaq29lLVkfiPJCspZf1aevl3WT1YvRr2lgUcAvxLWZLmyaBR1wr/PaNn5ULUNCHVg2m
MnUeiZuJBChNwCZod5NWb0fCc4m9GFMWrgXghaXf5JsPguNAfi7cjOxoHF1lSdX+T+XWkNGYJFxm
OmXdNcnbt5gDxSrddPANJey3K5FjYiudaT3PkNVVIEVbWMmnbQfKysDC4slgXATPyb04V5ZiLu+X
MU6SDXpZhilPAZNpxZrPXYoym4hsHKl0uqBsyKAZ1XP7wX/AB0NQ3UU89E1kAKddun6iALvoT0+A
7+GV6Z6qswp98Fl3xLzbkiqTuaebyozIbmKSuHTc9pKzRJaArmh8WfQ88uwOAfU2fMdafGo7+TOo
xuzbDdcQZJ9/S5KsgDhUZiQ00XstXlzDZvhB0rQ+BV2xcsDDPt1kapkRSXUumRJq8+hSE6Y1ARif
Xoq2X7mJJ5NKLS5EH4PHwcQE9K70yXPeWA3dZXQkZAvjhNBfEs8Fu+XXRRSwlBmR5DJKFhWm+TWW
Fr8H1NKgSGeniwgue3K+vxiyp+z8G8uq+YC1MNtutrvi1H7GvWqc6kSky/ZY5cn13MaQg0BapxzD
JK7A2vH7K1hGq5kFxhQAJuRfE2egwd0tXeMZtt9NUVYPxoYfKrw9S/c1pk+kiOSmRH0+wA+m8pOJ
ojMv22q5RPrblctu4wZ46UhrDceh2t0VFRZpLogdNwS9B39rFXgBVJztnMxsvO+qTQOJN8pXtEZ9
TAE2Owjnec0xm6dbYcT2epUAeVFKh/jMrumjs/5X83qaavGDh1fFkhHcJh8x0Xczt6cj+GShJSzw
9PzXvirU02aPYemz1UpPNT//D8ij1pFfIoOY/b3q20cYsXQf8HI5WjB0fzXUxSLx5mOceWy74tjJ
5q9iZDLdjoD7QMfz8KujgGkFnHe4VdwISodNRFIUPnsDHowE6THMQAfGTnb6M8Kgx6L2NkkdN5Sw
lNj21eawjdNbPnFxrLkWOssG6xPUc9kpnOPVomG+cSXcB8uRmDIMsLE/P9gLbQrVwFDL5EgyLaZ7
oq3Hu/wgP4t1d45Oizs62qMjwOXIys3T0nHbfpYZwosCa4OtMpn9+KiSNHNiCwyNeche3JoUotUl
OAXGM131cTwihkqo/6A8Nt1mlj7EV9DUQ65+0r+s4aQLTr5oK+XHUgcGCe2baEx9FWJzq9QlsKQu
mhs2owesnKmACEC8Aom6qzY2blKU1La1gGi5l9asocLfMk9K99CvZQo1qhCzxAxDHOFTdIb8zaJx
Eu837/yzkSnEZlynbBUGYAdRcYXLqNejzim/PcNbdzRVgqP7Z9834ghJzMVk0kdU+Ngo+ZWd093B
zransASxl9zW3mSwBQnp/rZESiRHtXHwbuaGoqX0Ws9dcgkQn7d2dIH3qQZb7xFCwaeG+qDbwXtc
StcZnhQ9hyRaXIsOJtvmSb2HSjwtuaReZucLufhfBI8WvNQkfcli7zQVPePJYyqQmcefHn+/Wlsd
gsVA7aZxf6gFk3dxwOvCJVV1ekq8f0duheqWDLpFnijkr/N9uETRCxALvtyz0LCYEl5ZlqYk8ot9
feMNdo9V+5cDN+pH+x1fX441+9Rw6ooMIU9FkUXkWsH10AsVpGLf8LRiJFh3Bm38VSX3q5M97QAA
T6DaXndj7LjNnGKd7poVC7XqlIjI5YtfI3ZV8HeMe6SVjYqMP7N20bstv4COqdrMGxuPac/hds00
k/swue3m5iuu2WDHHxW7Sw6n5abQc228deqoUp5QDv5VuEsZy8VxZnLOmJniTxImICjaOZGS+TFT
93NLtCTI8JnM0ou5ksfFOBrDU/lx/Sh+IujnLqeYu6d1NYv4T6ntWQGiwzrFn0q/w91NartVTdAl
yt4tkrNsBrrLzY8x5qsnTi0jEOgAvGMKBWmxyUcBSKIqeLMiDuLEK4kyY6JYrabILGxGxzdqGggJ
3aKTnrhLmrex0iyAVcWKeq3y4y6Z9GMn7yr2bUvk/xGPkXPGzuQ1gUbOK6JhEsF7WDvoIbrth/zC
tRCYdOujZOABfRLtJQnWX3yD///JBIC5oG+IQyId2gsUP6R79KbOtAC6I0D2Xr9bjGflSlQ2iCcA
D9EicHchkOhEby9i9XylwubeNK3E2z0JZNFC0YtHTkLFMaM7dwbzPSGhVgdG2FMNGhDVtj/2RU2q
ImcZgj/GSqBrTzYz37c20x6OuoAq1MJKVNpVo9b7GUlHz36F+aQI82Qwqjur7z2aa+H5tWbl4SYF
Xym+MOBhYsuthcEp/yel8naAo9Moc9JrHR7Nx2E4hv6yGBGtnBi22cPCLlDrJJyXoSg7d4lXe2Ru
a74keeQRgk/2ywk/2Zb/6mewRrNUy2nf4E7ChEbSVEAXh9xC6z5WutsEEwSMK5Q59pMaxjD9s2Cd
sbCworEyDVppnsO/XGdUiRK/Wy9H1SvSS3m4x36hhecTR3MvUBVeRds0v/ZSww1dy3YlYp7l6jq0
r8/I86ueU8PxkZbci2pb/s8zjTPGT2/sRDKr2KpzliFFjsDxpNdLQaD2Il1/ru3vYc7dX/cN6MJa
Xzsq6qfarNGCRVugPMp7OUA0X/Lq7RD9XBsMm3CFjVVYU48e/aocTfSHPz1Ez4O7mi/eiPNYRTz+
YA+b92oFKGqkU6LHrSTCxxaEXwsRJeFyEa0QZ72J8XuLODVbRpV6J+qiGP86ONrOZXv8C5ZeTgPh
RwA++XLDvyKTEx+2gOCrmsy0HqlKfVGt8tXDmWUI4NNE3/Agbq+21umumuHqTgHQqVSxzNJLtobH
ijnTdKc21nFVMnpdJ5Ho9bnTux1Ec/A9WYCZV9YalNMOGocBoDoMBVIuNglnon5h3JOx+56tVVVy
Wm+hMoOCHhLza5qS2z+vUTEfcYde4yMyeiEy/0vVj9RCFGHe4++Ba3RFNwAUemSUYVyYuLRrebCB
JRK580sdf+lX0K7bQ8kV0LMZ5ZCm5yyiq4C+WAM9DHri7OVvQBGNpfA0a1fgwhe4IioLNBVxP2ex
hU7wTFtgjIPZqF7EHRtAP8wFxPzOS1qWCwiJ4FKZu3eEozklBqh/q5X2L6wMtiRECO8wtJdWG6Gv
tiaXuhCfnkoh0uHd3Pgjb2acHIQAIobdJG7SNgawXEJ653sq2cPhiIZ1j/tUN0utaQzQCNAxqIYq
AzbQErSXrk8nDh6oCbF/VG71t8x+ZTAwMB1RDkSq0X3kOSQ2bMj2YTdlTsLPwQPHv11roWRNSU1y
8jUWBADIU2w1lqxI1uz68vdczv0jBN4PYUXOwkF4NdpGIBrw8nsLb2jay2wzIopoeTwIwYt5Vnz5
dZ9JHAJH66k1MhWG1RBNBIxAZhUg35PrI33KrSf2bWu8KtHsVuuJ/HpJu7VjlrYcfY/dCWx81U0P
89vWBxTz2V66W2gDPELgSWfr24u/IJvQp6rkm+Px5EL1PQOpyHnTbbyVlVLEbim3JcW3rrGUKbBf
HOqvhKbBZEebRKwIlZlWEVJuePM/TDSONEoV0xIRbmfgm4bamu04wQBH1CfK9az6ls67OpGTvcY8
dOXEHDq+FR2JQwn8xz+4kxIuc/FXyVFPTLI+LxOzAnqOfq5Nmh4zpxCgg50xhqohmHzYze0mpNWe
RN8qLKz2uWUDF7bzzwDzR0JVYSIQXyAx5X7zG1+K2Chp2PJxAXD4yGF6NKsvFpRSb7pC8Dcz83jb
eOc7boww4fPM/SYKUHoFBq/fLgcds5pnKmcc/7TG5ueLRQjEH6acM1HpMaLFclfBDSZyUJLu5fTO
BihnOyR6qBH4SNKbJ27LzD0FCUakFlO5xFm1PXjgtQO85KCVIlTApuSU2WohmON7DGVwpl7//pmJ
NgX/6YWPJfi77vSasEd2qjkNujAXdxvHIL/J1lx4rtozy93r3kmwmbJIRS8BAZQ1Y+PH1SjaHBo+
7Fz2lsHt0UNz1j2hH3jKaQIsFtCv3YbmiGiD2vBI+GvHAwAuml9qg21Gfy7tVMNUtGHA7kv+rj+d
SFo7an60mZEcfxyGpv4CuFA/abp7E4yqqoGek0k4g23F1KDql7FApezqApoS55j5GxfXLeXx5o8W
mLlPrmI68aiPuM4v5oluC5DMvUIZAvg04FgkcIqGM6zj/TPo60DBzMTMiWqu7fTP2J0fqGX1ESfA
TvI4qGCkSa0drSjjG1Ds10PAiyIND3PVBTGWire+qOzTaItUDEOOhM4zeUGzW6cCHK3bW/acwWPg
tAEl4rXXYcdI1WF33gkI5odFXXGQeDjFKgNZFFFyennVyKBknuxA8NPyT1BNDQX/Uibcy5Bj52tz
ohM0y65GSsI+cFB9nfEIhZAzwZNNAXXVskMluNdb6lSdRjOLhQMxZC04O4tvBCmoihFpm9deL8a/
YG9MsT/xYmR+lZ2gniR9h2Yr3I7x7Ys8Azx2VZC5rrbStGUZk7MaGr9YoQ6I7BBHCYuvDeO1Nyvl
3DwvGfyrw3zD/JrGhp5EKr3cqOLp+Nz1qz32fVF1d7abRSr0mXBU4HOIQAwWp5dNMFWq9et4UrsT
U5X6smJcwZFOe51RrNME5SDpg2hC0yh7PCFaSVWzq2JSR9q4TB/qqBbpuVTsccjytSKaVXnqy8Bz
2+YBPfEuG5YUrYNvYTOH2c6CwbD5+iWRKHBiUCpT15X0H2k5CCb/7m4uHTNN15v+449jF6kNp1eH
kC9mowKI0njceS6BIyZnYVuZwr+riF6RthTTBW+CvTe6C0XMWfqxxWp++tlbXb3YfT8gfsnU4xXD
C7/QiLH6Xt7NqhY7tPxD9mVhD6AvDYgo5BZw/Wul/smGXykBQUqPKC3hz7ECOA7ARLACBZrs4VJF
ltDNcdthSqy+PhLULabGmsmKUeZ9MHRmLuEMchvyB1BEXlnKipmwPuI8YTDfiSeQO+EtmfaWl7QK
ZFy+HQrlOwjtM/0tp9TqRFDFazEfyDMt83QAsvRFduk97uM/Ih+qvsWBzu9ViR5DUIVWN7oOMZym
10SisgHyQOT2olnqoShSkejPfThbrew7KpFPOeMZ+tZcDGshPxaEZ0QU+J0lm4CTYS4GYtbxXEbh
Xp/oPsJUwGbJSv69B5895xReEC0AMx9nixTjoqOvpvbCpTXCZPe8IcQMHuNvSPaDsiZeXmIe1YX0
PqfeU2KRZjree6XuNkYaZyMJzT6K+uFyuvRW0Hs9erWGzQrG7gWKjXZ73Q8/QqSGLgWOM1K65vV5
rocavaUMxdn0XIUNMng+leYwIhOQsrLon80kFe3kzNmOSLChUU/BVdasAe4S7byfYILOz+9hTQ2p
61mlMhJA9HXGsXcsKHphFsd321hGFr49bvOy5a2D4kJvTUGl6XQdPOdBsmIaGEtPE+4jRyKhD1m5
i2FAVNqj61O5gSVvTKQT/AhHyJzgqDwFsbzguEAeCzxaK5DSuJL1gvfyBES5aWhljJkAeNa+63eI
S04qg4MaqCsvhIl8Q8O01EBtcQcVtzjkAH4DqvTl1m2VjNX5HDHgIQ3tTuQB0q6/OHG3mszSI3A0
GXZJ4dmFCop7S7RpSXF4Kvumws6vmaHSUfcRoht7Pa80GooeCrBeWueyq/SwD3/lHI/PDY72+SI7
A+2PqM5y03Z7AUfHBsPPbTJewx9VbwsXNeXO6OU0qCEOcyG5u/GojfYQQDzzdBFFI/DyQbLfGGbv
JfpBJ65GNGPYUZven5g43NRnV4rZGmcx7DG6olQqPyPP4gTdnS5Qvzgpe/kqmAotp7fsMvJ+ZRyd
XbpgPTohL4h7lMZ1smRUGo1gMR5SzPGPhU3NMSDO+uzLyAcJ2IC5r2QiHMFTUDmrT3v5o3W2njyi
mHxB9UPGDmMHbM4pStvT9qKlOvbIey3q8S9ugEdN2aG6Ylx1fDa2DQMh/Opl7+gC+9VqJaH+Wt59
hC4gkGU+RjrFUgeGUdk3srKrOvGd5FrU4jDCuK9XWzsC3PrvBpbPLvG61pXRbMXxHsLyt7+i9gle
E/YA6PJV73C8zcukg9RB8yVgZYrHC/K/EOB6JgOEiLxvowWgWdmF9zm4f2DszMRGyjGXlb+SM6sX
ildDK66tWb6nNflUJ41dRWWarB6Iwu+s14KCZXn1F+JnLzLauvMwRokjV0Yg7FuSNsn4iKVqyccl
sY8GfEKe2kxJE4lHKx9flOefFjHTAZ4CqHAJz3wjcqAq2kJytebvpPXJQlZKGHVMmmWmyE02qrte
XeK3kS7T1tlo7YhMC3Z14WjEMLat55L/QgI5IMrwPz2GrNOWJywO4Uu7I4Wez/R6gsCCWihNgnOD
8ILjCNsyT+/Xi9fqXSNe2Ij49mTHwVR1RiGTBpePDm1IvaFxIo7pkXsd7xJNcZ+MrP3rYjS3Ktve
ObH5A2AN5nYhi0DxNNDBwhsbnRdChLuIVagXCQGYpWsxzzpkxGWDtHgb0OKN7+K2TZEsaBeelVjz
l81Zb3tZ5Hmy78FI9VWNxjjEj3VZiYV4I6gW0neDIU3pWLflkuDL99tUgSDpa5s0A6Em5/Czh0pu
t2Xqv5bTFIOBIjruxLLJkaE6CqY4mW/pd0DdAEiZKuZGFk8u5IS3V0CrqmWfGJJkW0ogFESx/JBE
qDdJ0KXEr3q57rEtfgCB0LFgQk4AXB8A5dAGos75FrhGi6F1XAX54sUKand9PmuLRQKAhiLKOLGt
6mS3pa2oZ5bZsvKyc9p4qgM0JmZ/ETxQpgN9QtAP6rSrP/3luazSqERKZtEeFGgqN7kLInwxnjLq
FyGc0CKVuXuEWWE/9qCX6wPSnVZ9UsKQ7DapKEtrynbduRopCIqReYLxH/XnP675KjC+m3S7mbwo
+h0buxOwFzQUfFQo91bBP9AiiznwU/l1P9CNjgc4SQWgq4DZRGRNxyKS5Vo8qU5MGTgmTULVgfPz
qa+JgXENJXurGwA42ZiJ1k+niOYGxZ8hAJ0WpbcbymJYBngb3pUgl7dsTcSjXNp+JD3/OMlJDAfn
WmSFyCBNtgTOyZaUkUFXZ6HnA/cNBmByyVukzZTNGicqSkVxJiOtmgkkvecX/BZa2fwopY0cr5Qr
96oUtzmbH6zP7kf0HY/BI9ethsfj+GlN93/lXoMX5QXYRg5WJaYaoN3ii8SQYevcrjicOs1sfObM
9c1D6H39Ez0kPT8XbAy+qN56PIjg23ywADheXAn0+oDOQERlwGi0b0D5/BPZYv6ZzLEqNEDx4wrR
kTxabYlqrMAxylK0gpGRKin91frW+Q2yfNFE8wip8Paao9pr+UPIdpwEGZIxpwMxJGioV9eXIVOa
ziOI91IKmF8iVDXuWcd/k5XatiYUQ8k1d94Ufa/NNj/wFR4DkZiKqmTlzDz7gcub6gNMhVdA7Qaq
H6kQ9AW0/GsQ7hOF5GxFbcBjBOwryE8UCaHY4R/DJak8HxQN7OrWC36TRHJYhF0MACwXtzOp1XTx
FjrHm9MnocBH7GmEyVUvwBfCYddfw67vmF36Qq9U75gT1l8qlcu9vNBVTxk8KwvAxQEt2E8tOgii
0ZRN/+WzDQNSiGv9Y31zhKdLJjsth+xi30Xf5vnqn1FvGiA6sJFYkyFVWLkj0kLs6FbGQQCa79J3
L7psorQhoza+Rsw1y2VEd1F1mBuucLnP4ZXyiNYJblvAdyeHRCKlApKPG1CpoPxYG4K17JUVeynb
0gDBeg/W8FC6SWza3fpW7auW2McTW5o7Lr18THt3fh0RvQnfRbqkAOCbG00gAGaw0DnS+kD1WYYO
G0HjPTKt0EnRiZ7dFPegDki6dot4OKZGIinXT/v/JuyR9nicEcW07KfEO9Qe77f15AzNs7g4k/dW
G83Ii2VmP4I1mr8psi58CKpGq/rHDuUNwBs6Kx6RixymZPb5Dlk1HEdeHkKSQxRlwt2bcHfaR0CM
ME41KMkX9rsihmJO3K/SRKiVKg9EDgjrnkR2VlcYQO8IS2aJaD+xrdsDMoEK0lLO1kwz4hp9KzyA
8/ySBZqj1ATy4r2+zUN4cBmj5eKZqN7HHJPDyG1EeptwIMlTEVQW+0uYSAfA9FOy0yUCdnmNS7XW
xq7+dYqAe1fB0+YjjE78leUmLVzd2wIsBQxJKfEk+6MsF1UF53Eb7e5FB75Mo+EvQnV0hoF49TTZ
dlGBFxnKsyxS0PbqmOm8WWEknbI+CEIzs2vSfOyEahy0ApOT43fhQCt40Cn20WiaywWf8v/zhVI+
4RDCisk7R/cHWrxP3VOEfeG6KE2FmgGUK3OZQ/g7fHMqdIDVaC7k8p6KY5tbP1Y3D3zUsw5wyZkj
ADJmjbtl3cc4HatvtrCuwHR6gLjppDxVtXs+qBNZSQZZkc50LiXxpi+aYddIkU68jjVtyw8KlrpJ
egcdGMncAGo6HGF86zV2B1k60qJgYIAhrKXlePHPKLEbHKDGcypzu8fvLGuCFsTjN4VlRZhXSsaM
bJntBSrv8MAJPgRAcOfe/lrz/ldiLEpTAMS4Z3ryz7zzyDb0G2z5smWkNVhlX+jPQ8M9/kly5SPD
OsG90rXVpJY8/njKzgAH/bsQlJ3IopCDfo/kjdYXeLA7WU9VUL8tOv1gDzr4x95GDBQ+8Gu20fa0
DviqCy0kZ9Z6Z3d4RtNoaPPwc+So77R7F42TXnrzgfdbMywmU+FQQq1aMtzbQfOyd3FEHhzX0q5F
xLxWRvbGjeJW4GVqIbvMg9mSTdXSghXJH3HMEwFD47ftkG8R/9lOep2g8FHZJn0jEJdgeVF2K8vJ
IcmZfPrfvU3xhYdxrtQApwxa8JgXJflvP8GyDwQJznu6ZuG2iCv4H4K+lW+oz38CYucsX+ey8EYi
aj+feNsvfpGk1RtYdFFsIwXA0V0DbLElvf5d3Gm4II+STh7HwFhezTPA9pFrO6T2NDaouMEEl+wp
o6Nej5rXe3KpaA55VV1lpR5WuglDBhMi9epZizdeX98k5QinZN24Y1W2MX3Ew/SJpeTCzxf+Wxon
A/M/Gfs+BjLmGUzPDndX4ozZ1Ie+yaG3hGfb64NRuzT8RxaDsABWLDUzt0koPygHEFt1RCVkWkSA
5osPQno6kFVr6qgsSTTm34kEDxr/a6UQVn09aPnUox2W8tZFik0dgG3IA4YZRFrKMGoG4lGbvg2T
cesNIFPuefpOkjSpYzY6b2xd2l2PSJoBsoYnRySCyfttTFO1dOdXAJKagoV4NAdP+LG3lUA2zWPm
p9ImsKqlU9GQ5+29vsarrCiIOwpItDIO5A+3SUuljMboWKz/J4xTsZ3fYDNqZ/RWH961p7n1DhQP
goWdctWFCp1E34Z+RICyhBI6hU2ei6N5T7apYY7uVXKciA1I6oVs2Dyof8/KcZvcTxPNL9JTf94U
MgRDgCFv6VG6U7K7KaJpscoyvCDC7zEp7+u7DJYRaXcJoLy3OEoiPyeDOHt/b6ktnpv8kEDEj6UE
j/m0dBcQf92fOZSyWNV5CoU916dxvF7d1Mq/obW7io9OomIAf86I4VTbsz7KCRTsNtW9sWUcgv+b
XwDwCysIAkC32UTEdFw6iMb4R3+YWhq/vS5fgIxD8eiaWWX4OhxEjGcFSuVH/bmuiXh1Zb/bBeOk
STAz2lUlvi4no7u0yHitX7tw4gEhTaCAbjhJFVTnQ6hbgY23EbvMy01Ow0NYFZVsbjVGdcDPBb4A
KqCvvQczX9iWlxQ8/iSXk4/bWI7UXUxgYyPMWt3GU0EiytKuF3GxpkxBwQYc0A+D1IdpoymbSlIe
Jsy0Mv5q6N8MHMj40r+OvsPnVqH6CovsYjj7V+PKnyRDdfnL+FmDOsy3jjxI5aZfxewrQYDX1On5
o8zntu4oFgxzOELpzNtEXXoN9NYHwQQUTL1vWZRosIt4IS+TNzidkZsYaSmlchS2EZhjohdleT6k
CwetQe/kE3WQpjUlfd4DuZmrs5E4Lil5KPRaaN0NAEX++CuDEozmoS8SioteJSZZLYLg6H/5vA4x
vaxzcwbSPERlUfVQE9C17E2lIp8uSorzL7igy3ns7VIc9YkiAG4wBA/SkCw/CwD00UNvZrA6pOQ6
zkIIQQcNvlsV8X+2QOWzjTtIbSINl74QAPOzz+FirfemS174stnFpOXVgrR/NI0Ss/snp6Upi65i
DMqXnpVk42XUiVTwWXsi2l2APh6q0SRIgC3hGwageEPRbfSs/7fXJCGJRTAIf2N7yEbYL5i5tbNB
L/N2JlQkOkQEhXe04lb+dfsNB2ABUT5crAdSCtalpv1+wq6in27icJw4PtHvcqXRfOnkxIeEPWx7
Q6no4div/+Iprut4MMSp99g4IppkHpAouwHoljNsCcBgRGuXeEgFip5BnAcMZkMnUmK3OwPW+RTf
xaHP19txbY9iv2DN0ohT2/9q8KOLFOiE0Qo8AJkeThY3iHUV7OmpLYtcVBm1/fkvCqoBcpUBm7oV
/YxP7WiJZ2iJU+ns+9KlMrUaqxdUCau0OSzSCmIcxtJ1gA8yZJaUiUMs0AroZoShn9BTcosu3wYb
btxEGSzE5Cg3AhgeXBs/gmaGiXGCQrSL0+lVDvAXC0eKeokM2cmUK+IA8FPIJ2qhtnDKxhU+Gb/e
md7xXgrkQbYgkEFaGHK6+uNqSjkKPt/ELePbFcKDIK//EONDY1PCPZmzvMfWypTVYr6TpoH/ZtQ8
cFkCB5e/s6NN6y1F3R4PyRYMbQ6uFdNtuCsqtUGydDh5zYOV4m0TtxR7qYOdjgpVTBXWjCJKPNb7
CbpsIsSmQ8oJZcqm9NM2WKdCxdK4GSVNUJTl4pIfnsvNQmezgzS2O/nduLsGBZyP1Fw16pwUS8cB
ngYWs9TaE6QSUZXmuDSSqailpFLpfBqHV1iOH2uA3JehXA2af/nQb4/cHl4m5tijqOAwBh44t98c
oCzGDNuN1j+H1RUdqQyQbBluddcUMiDf+g/GL7B4upDP+HS0FL1nOnfd9CV+OZJrakjPCb7nn3W+
7cmzOkdhUEFJyLq66FaqFs89RXU2ggUglAgrzGilwaBBBikJEWMSzvYULmCj95aqRx+4yoc0TVTJ
MEDumtI+ApFGjGmMI/4I/H2MXUMsxDSqxYZDcGYboIeTaV8aeJMqSrhcJJe/sw3ifV+8iIs3G2IY
9Em105XwJ7yqhP0UNi6/e9U59rLW+A/bPk1MydcYNACTHilbAp8vFK3I4KqJ+6vY4vr24GbHVPwv
5Kx5JeY7myJg2N+nUseoeDklx2JdGmIuXUMxNRfce3N9KbPo8cK+8FkNMKsoPLUj3KVC+ArK/qyu
850svZYIjqjxKb6DjppNEDti8Hk5zZkvR9WN6Kp69/YIPRiJKoun+Ya8NOHCs6thmX+2gHz86jGO
OJCv6wDTF/neCR+HpluBV0Zvv/x79fZna7lZPFGe/gDPuzuRNmaZ7NCH2W+4KD0H/PqgLNEDJuyD
MMb4cK43pAS0A4OMdcrc76puHaAqigHWWTwuh0QPcbShs/Zt5EPtrxtwDYXoyxL68ITVUfdawlYQ
pswxji2i0N+b4YKD/Ot/GdIqZZF294cPNTApIGABL4rNzihrvwqRA6IW6VbM6hATRmgAPWCfRjLg
hSAlBYJGDFP0jrzUaieHk6S6s1TnxP5Pkks5Yzk7gj8etEc1ok/HWhuhQZ8k6ke5RXtWB8ER1YH2
sqT4cy7ySekAtyNYPwpYzf6Mi+JjXsE0tmxp9YzXFc5mDGA1mVCGCqjZlLR91sONXFmonM3FjG+/
KTZfkwuOnCL6TDpe88vh1U1KZtTaqgT5LrXKA0oEtFAPADkSq3zpm9FYusDlpy9EoAKNuglQPN86
tI5PKJWw4jVr5MHhLJADjJ414Vw4Es7WUxS7et91f9UE8GyY/JY5/JxTpmP6G0+gJvlnvo//Ca5H
2hzbLHNe3MiZ4g5wcqklEB0Cu2PZ6/XLxR2OUt46IuQKy9UXuUWycuzh1HKDQ0HppWKymOs5Ncu5
xJ/qgTtEJd21EpqlUwG3jAS+YaonCP0LEY2myvwjlOytzeM+Vvx1tyjZKQH/TRThPtino9+LmS18
q+sGrXCU3c+mBYl33d7FFYLtNIbcqpQHJiGBY0MszWG6hHvXH5n9CFpOa5XaK+tiNahIDky8ItXs
znj8l6i+qTlscEeqJVAxpFEntBnIp2k00o+g71H6em6DQ0P4wauSGZmQXGZIBhOxN9INZfYHxz4a
JJ1mpCp05bIwobbt4lFw9k/z0VyWezFhJ1BepeeBc83JStOAx0SkBPtocUAE7rp5npI0LQab3FzR
OnLp3Z+NmyVdBIzUD8g6/pNQCWY4dPlsjFxO2eIVOspR0L8KNzPCoqM5dhPvg8BKDK69NlCEhJ9z
3Eafg++ajhwxZJyETNOiMUZiTseK5IzegM0KnqSv/M5iJFp9kLqaKkj8aVeVS7PNx0BspjORaG/P
A8wK2tAIGrr/xoDAAIhsZJ1vroJLt4lZ6e9i2d1RZ86rl092S9XYx8O7iGQSV8m05ezWZKPvJKIT
rpXPqJQu2SldvDPIl9weqiLDLrRC2/ujV3IwmLVWFlQpngdnsN/excNqmOnehfm1/HWPxseskD0m
HSA6HZMaUDodzV5b4HaK83EWYYwLHYIxWeIg4Z7zC2kmxRwwob/aFwzWFRsQjb90R9lsdYlRim4O
w2A2VK5pdIEObvxWA4fsHd2hraxwMm437bogotZ8UElEhhjMpS5TY4IBwecXzVph7IazkwTLDCuA
H95CDoUKeIiyPwrR55ACIVqL72pcswhm01oYEeVB6AV2l32OVVRWYbcjkR54Me3JQ6zrTftCMRAM
4E1c32bwiNpka6kIs8OMqZdoW6WSTfAhK/bT+45snHizpFO3j1lBZ0i6wXzV5yo/0grYvXG0cqi1
s+XhVW47STNxb6NRpjUbsrxJIiTWGtl1cI9a7rJ1VDSnsJPosZ8JkHZ7jxyKsicYaTE0BSX4i96u
2VeQII5UzQS/YyDYMOrMQVVulcwGbmIAlIHJl6fSj4AmMcOUNV0fDueOdGdG0RM4VmBMe9JiVzA0
N0blN5y5AyvZCROoR6KZDKOLWxqxzaN3zKIQ96bESSSMw7E14ZW1iK9+J4QrJbNW766kKQj8oS6C
FQHV9klVAhH8aO1a3/2UorLVVJX9Z+HGFinJTeZ/sH5wUamDDmx2oJ98cFcHu729CxtUzqj3lH+b
Ttr2GgAyRcvj0qpKcwSv2vYMCxlPfJRWIyUDUZopWB/mo2qNdmH95qju8zGE/1e35KBTIuepopFM
HerJwJb1rtStXWOR1H+lm5U1yOc71F7Y2kVFjcEXOr/OKKGbOpsYJS/ntqLM/dLiwBgegCojcluC
BwnDlfjk7bvn+dAjSGyggG/nFGHWYu3ChlehJW3oQFEIKpPJ9/KmIUj8pMT3Tq8RXoGNcWfDdt8u
2ts3si/72BkFU4tUiCSzpMtlV8pZqGXakyn1LGngYdaq0ticaFdBcbRvK008XIcc2yoOZtOaUijk
935OHsTszSSJpKiTouK6Q5G1rdmcgnI0kYs6rfOFTes6fwjKMdbFQSOHDzb071zQ8NQ6Bc6YuSPx
xcv0kOnJEEBfxJa9Qk3AvpGgnbTiM7kGBYSVsR2Z/eGj1tJzJE9m5KK0zQWhST5iqkomRzmiKKzA
b8gpZCTaIra/Id+zAIfqD89eKdSAP34q9HM8PTPCDLU8PP/+UtUARYtG87wKAhiZlvGnwwrw9/ri
XJLfKdJGF4nTlyQBQNobOSBUVSA9iPZT7yeUUeogkpimREGrlHnLebrQh/bHzXnJ7EFLh9zZcBD/
aUxrhFpNeSjf8mKeQnjFM2c5WgpPjuRZV7yNrXmHbP7qUFX12JO/0jAD8dv7MgPlG2Y1h1sYN1cN
a1cWGPUt1yb2Z/SiMa1nOma/FXLcnbDHPV0l5aXYMCvPOv4QIR0EEU128kHIYwqCNrPaAFbSF0fn
cn/4H90xxG/MbEXd8RxTnYXxi3JEj05HjFXIuswAU+wGKh8wEKukf2n45CyUzoget1EJ/ecvPOt7
btnnCdy5eJX4SSZ8W643yW54p2kY7oAMmwDUIAl6OThRBRYykIGQ0LEpbRw8iSNetA6c27oFm/at
4iFBNDcjKz5EyFQp1LYmQt0nxXEQCij3fu2JekRZE759x13DBurJi0Zbr+/jYYPyrTYLdLyNrJHw
No2x+2fN4Ve+8xsnb8LV1gc4UmJpme11rJo0/XMXVbDW9qGCQnFl/ZuO8+ZH8qTltEXkekEYZ8J9
l6iypfd48S5nXzeHq0yYcNRdPlOdrQitK0Gf70wlIKCuUz1v48Hpb4fTOY4yJawAAfDJtN0R/fod
B5kc9vM3gGVmo+e7CrJDPUdlICC+RmQQ98dBVP+FGeB7tFx1frxZ2oKIg6VExZW1JXKW5jqh45tS
6TtPLY9hSfrBsKSSXxj7eXPc6v0mTmnD4N/NwX/GWqPiIkSE2QM+A5lh3iR4GbfXaSWXduCFWS9A
Uw+gFQsVlHFt9qTvx+fV70s/NKq48G9eWvJMgChouhczCBswcB3eXXi1VSaiZ0E5w+dCL6JINJ9+
luXejvg4aC7ICZrrS4NV63J8Kic8AznlrUJmlBtnx86VNCvDnmJTJAo+CLq7HTHooaMSuuDfuf30
JcF5vNPOjvFUeFf+f4QzPZUmZakrUjjIMMfrNvaCkP8+hV2bQDXrnCx5R0hc85KXpQUhJg9ySJ7f
nBmU6eHEqwITXqaA8bjbRhFt4HYjbkb0+Kyc0dP6Fxdbn6K/0pbWoE8unjcLid3oqRbuhcVTocfy
86b/mcOJnHLIXg/ZVFhvqDDc5p+v8eLylue7kAs9z7t7VDaHjBm1e2voD5YYzW/bRcvJKooRDKMZ
4VGKFXrFp1i6gHn/o+3ZMQQLM6V675hFBZspefe38zspSRAYjC3uAbg7DBzGCOa4AtGRQbW15vaT
yb2meMOFE1vaIPfa3hlmlbZv1eO9+aM0dSkWrwYKR/mE/oj+4YMbOZqKQXhS3Mo6D3meTDpb5tX2
P86iHsm0vKS6I+jiMDTsyuE36eAqarGY904pH28+L/5WBtP8Nbgb7KSAbujDjdvtE4ACRh+HphFj
qttNMG1Eji9fdYKEHunjm2PhHxmiO3smGbJ55F4r5PgnAAcWkZ2hGlImyZxOYicRLgysYSgSQA2d
h2GqflVfLzyscJ+j1fFu/E4jcZMOUuNi2+FDvHHHsgzKnRzGVakEkwzgorWvYlO3g83xsOxssvBn
Y2DWeZJPDjQnvoP07r8GQgSgE6iLhIsEyHrvmwlcGvtdFi/q2v1SRrgKv6dyTL86fm3n8Cc1fsXY
K8CSnCeHXqbHhvdu2oSwouFPZN0sCkfhKjMf3FptcpFs6N9fCOQNw1Ral/UjI9Ytp5F3klLyigND
67/w/OZ8Ijw+gm6FpCnBRIeOODtYE3VjsVNzDwZIyIhxU0nMh4UfeE1o6HZv6ppqz+GvMpG2ZxR3
SvuBaQT/0aP1+GqrXxI/7L92cLkAiuv5l7UAHjLHbCxw8I7xRXwW0JxJYa+w5Rf+4cRjAM0+3/ll
NNWfypDQfe5BlTGTTtAloJgBI2bwjbPai/dSmWhQpg9oYvqRSj1WmDGJ8Bx+nWTERbC3CrnvjxuX
1zkMj24ZgyRmXHPVB5M2qj+RpSbAfLPmavvG/kuuOM292SGsB9EkCvGVsnEk6+Su0XIWxEvinRTT
gTDEb+FE2uy4HvJ0nwErR2Y5ivOvlqWgblRpCLK9U3x+2qjUEjcVEWV7QQKoJd+iE+cjLprDr5II
t25noLoTQMSu+IiKiEEuoZ8r84VK0v1PnzeONjhUKHiiEks5ruuneTILqCJw/p094bJHccicWkPt
0GsdPiVXlpyrXKrZpM4zzoBe0leor3u69bA0uKlV5F798HpWRZuUE4eboCsmnLWAAS7IMcMRodMI
zlJuSCUBmnmHJHNUrxR2IuwWZOD+f3Y4mKUyfz/dVjmauUTtdLOYHRtvSTv+o8VVdhy5r6no23xv
bXEkxV3fpom4f3USi5WALJfGh1Zx+yTrG5ZKSBAfPFyKiM+RvTOI5skatRNFfEegb75Ea3PPGlZr
vJUJpczusw6KCt+5GXYr067CMLvjIBiaHqlAsvn/rI+drv5AvnXOEIZytvBbDVgeOJCWVIpi5K8S
fZG9uosgosKULBbu7gDE8WvdRp6JPslK3h5zJ1J0Ln3dU3OsAOk95vt5g67SMKudqYnPsRmcG0ym
cL+T7dYMMgDpP475wp+YcTXiSWoiLIzpfcFI8/B78Tl91nWivnen248qFHacR1HV9/OEQIbCYFg5
pt9B4FlgMkucdoma/1x6rc7qfobRofrMRekRAmIc1g6VEAOhRhXoGG6gn9XwP/CI28wnO1J6BJpy
qgSa7HAQizmmcgR6UNOVs8cmYhvwsDBkK0p4j1ZLkuPnHVu8yahm0ZvfWbdOUF/5kYJhlcOXdQKv
rTdCPVHbLoyWVbtQYjPm9bUyBjvniz+5yEFZYTnl90aCGAtVSqTgP/CjyWbdtldjMWSyTSpcSBP2
7JQudrQ57OFi5Z9zugBzFIybFAXoVPbbKsZSwjQZqO7WyvhDOJFRz7WL6+Otizx8fvxjraYDc+Nx
vpGqRUFo+rtJF9IYNKlhf7Q5BkKVopQu4XsdocXVz/on1GGka/f5/f12CKbJRtL6MO/JrWBHRU2g
rqtuQXZKRCkZTH8p0kHpeZ0Rd+lqBjEX5wnu3eaZAx3Nw0/iNLAoo1oSj4USIvkSODfdYRaw3Dtx
JWnkutKUxjmnBVM22KFYHs2MqVb7K9n0obhTNbI5XyK+T1Ccp2WAPKur6YzU/+eDf9eBN2+3QFMt
fh4k6mOHWJTggfR4+CFxvV+kFyKhM6fpw1rIhzcUMwl4UnSZlbYstHh8pCAVu4+nBwdC2LB63Hrb
+5McnWLwRRQMeHiWkPuZRt9oCrAsKWMq00Uvz243zcp5cU+Uw/D4eFGujZ6IKzP3qT1yt8Y3eP9v
vBwGaWkmd3MH0NSshBvGct1PjeJvJOpF7qAPSvTzVyYtGRC4mibqUeVs7HwePpQM/9WeExQPv9WP
a+4qs5FkqCikWlJ6ncN2ln3aRirz3zmn8x29sya2hlKOOO9uXgUmv8cJ8HW4jnQcxIFZNj0X2+uA
05bHG0fkfIkroAhgrRfEyayOivul0Rz0bx8bsUEG9MsU05ZnaiFwzL2O45jQi1HgV3AeOKy4uAhu
XmqtfA1RyrEUcqIuicPEjR3pKPlAMTiOk4cyafBm+vLZBNJe7YDWc8oz7QSjRZ+S8L8/37KOhX9e
h6BmQbiou0iURou9AH9M2HbhzgeEK+8x61h6Spgi84vRRhngg6Uix2jGlrosY1Az4t2EUFLq/S7s
y5C1e4/m49lao6k8S6L4eMUJ19322fihDBqYq8T4wof56CHTvM/0P9E982NWj4W8MN8HAv6AKHvd
8TQXbAjjLxEkVQ1cqIxbiQn8cT8axdciG0Gk7STnAQns9yWsxloblazsX9gRWnSDC3MwddWk5db5
Xt3kPCpbHTzlZxl26xGNupue0DBWTdmZrov3IUxU+P8CqtOp3Au6hysI1rkPdpPENYPcW+zruPC8
4N5xs9vEiQr/qUO6AtQEK4bIMNOWcOGw9ISYFQB56rytgGpE4xgbjCRNuRG0AJ/LxRfzrNPyAPNB
u8L1MkbITMh7neiWn/klAdIZuRdkHud5I6nBgSW2vy1wIs39D03a+GlnbVBREI/Vw9p8fNI9S5AW
R+YkPDKCTl5QIyxJmyogPtyaa26008itWsXWqO3EB6LdpKwhlVoKy0atQvTO1f6OHFXiRpvoK031
t0Ed/an6ml88Meymjm+s/J6D7uI5h4ALEjYITysGVSfncPKQ+s7vePzRkXZIYJU7MlBBwlBgcOD5
mvU3tx2sPlYht3b6FDAJy4TugkeQMh9B236qFGqdezvq7WoQ/itsaMc7pVi6Sa9ThObeHd17lna4
phxv64mzrdVTwIlW5UuZwchSm0qsoOyY5ss5RH+r9QGJN7m8rqSeX/i4yN/fAC8eyM2JfvQ8mHJN
JxX9reEnUQ1L90qbAiDBzsZupPd4m1URrwIyIiT0TuUk4d+fFX/VkZ7AKSjrosL+std5Td/gyTHS
F0NpDCp/WlQR6ErCX7i1nu53N9P4nb0cim2uvUuF+cam7e/NbqKFWaYbAERrfuX15wc9GKVXA6Pp
Tt7VFr6zZLNgkIdHg0bnKo506Chpx25lMNlI91wiqBJ13G/k6s6yPezdGOr9bbK1w3dXxWwolkz7
bqcGLl3A25vAE6RO6D4cFoBR8vxNYVmInUebejq5DHnWb5ns/uiyErkqgkVhC4wsouM9TiELSQkY
d+miXkK/RNSpmgCVdv194etlrhLx2WNv2kNix1ciLPLsy0KFKDwoFI4YhXxnJPAJAkdorsSI/g/C
jrsi7xCUbHAFGQt0oFxP5YRc/vGqT+JdsyWGii4x98M/glUodc62hc504j1gyuYxGid8HM8Kw6R3
AVoXqKHtrSkBkP712CY3QuQ1MjtF7GvbFDqcYU37dd9Hd8r5/Rl2ixIxuXlwQQOp4Hhd5cH4elab
KGZOHlLkjhJbcgIWt7XuSgZAY1l78cr544sx/tfo9SmkNwkThHS4QB74P4DIBxmoe3khZmTJf75S
krBs3AbooJOQtAr8qMY8aYx041q7CoeWVD/d8zXivk2C39mPxotOX/AudbaTqrjH1tdjnjjBcI5K
yrVqwoC1aDPLJHbZT3HrwNS11F74fdbdJDnbi/o9YeSGwfAnXAVQaGjzJtHHY3JLqZ3o2M+MTvhk
JYYhZPNrPnIsgSSRA1Q9hJ9Bz64LyVB9n+rJ2wi0PvYPMVDX9ZyEcBQHHMYoZCcq8GVPbF1JTKUG
0mQ9thOppyLjmvvPX0ldzugfBaRhHsHh2FI6AA6112493p+m7HHqLKyuZrg01aQ3FVTQTcodDkc4
JMayjVOxpvsbAbCcrnxEBN3pp9CXWY+bPerS5M5dJghHiYWNLPSawKIGiRuKl/5RzLW7cQSBVTlA
HfM2tG7dAgTOSV4oe0A1Fr2eMgqQxoN4Kaaa4tPVR2fBQAGCs+TZXKDzQCloBIztWUb7uMwVY8+0
01/aGSgEsQQPECzHGKwPiaJ+o9fVMfzlUEtjMtrPRHJ7gWWNOhpdWzFZ9vefpLiljS172t8jF0sK
btwGa9ImXvvshvKFJAEKJpAOM29ITLRhKMZ4A0iFwwLxWi0RcLV9sq30LQEf6BTSegSXSEfGgxKV
gDDbkBpUxuI84JPauJhw2n4uR+wQs3bpRYQObK0vbWpG3lpk9P8oPfG3Woq3o62NaivIc9yFBLXb
TP8z1YX3/k/AB8Dn10VoGg9iGjQsvP7u0/j+J/SR6D4iMbhBmcHLIbeMVAjNUGKDZ9YsrVEG3B2W
Gk50D66msb0LoISxu5JgwhuD+Q6QzRigz3TakO7ulhCUD/5EDKezlG6SHuAiMXahr380+5CeO+lo
MHIUS7lCPq8BpR1h9nPc+4rRu1EaQmXIH/gxEYwtj4+ZEP6yzSvbGmuYWAXf63UYoBD7AzIfYyc7
Ha4u4OXaJz4EVHzcUCd33xsJE6LCl3WdTIhRdzHHGnMW4BmwR5fnwKdA2rv2saBp+rKyrpkVbQA6
79VOxJ7xmqkgx9KXKWGdDaGkldBN5mEG+GkuI0SvJwfh1NPCsDg4Wy1G2U25ZNNPJF2tyYwp4RHk
lWTq4KXZYOBF4/u9BOICUXO97TSIfz9FoqR0ccv4A49JXOv8ePdMqI0MgnZxUL8b8whLfB6+kAvh
BFlPZcCS4WhBKqkwKDtWiNR12iWSbQqeYanYVqZE/K73rtqYQGnt2w6h+svN6NdoZv1CoUuppgOK
eYobuYJGZgrsxNR+eyMdB/SAq7B5+ztE8FGBnwA5HPyFHxJJ3dCAK+26aMBWLPIHM1/Etrsofn2h
JjVh23ZMedmJW47IVqGMNsvpZhgFX8A23kmVEnvU+ELVBadkXz1nNE3K4o9v22bwZcjGS6508Y8n
jtdSVoX8bRIR7G1YNfOKGVcDFjieFmX44rtvLAoky6Lg7em8uHP6Xib2jsIUmLOKAaFd62VvuVjO
yTvg+6AZkAYMstbKH5G7IZQEvs2toKfUTafd2aB8KKo5zky0e8vd87tHLyDyYxlU5IGaFb3ROsIN
i9FKIW+mf7rZJ7IBfXqKdi8K96qf7QY9hpA1D4QBeK4kyBSzNFRudS4w45uGWZ33dNiK6MxJ3C39
Vu334foQ4LKsuSSQJGnDabfilx90yS34otAy+1C56tPbp6GwqCWAfA79e/CYm+NgwIoN0U+PjU7y
1pm/oBvJ0+RVu0pC88u2xIv/uaVIuoiUjmK6X6H9aTVP1cbPfm0YXEv2Br454ylv9vSsWmtyHtHC
7ZiVP9TZI/DAxrXI6TroihkOKB5wHOuUOB07xYvFKsY5PyxR4KhfbLrBf+nKM892to/lAZ3P7A5A
sfOJVFmQuQDkG6GlV9YDNhxbX9Dwe7SFBoWyt0/a0eQyBRfRsV86TTVdlNg0mjJ05ymGQj8AHFc/
dkpCpHXJruk5Zn3TPar71oR4sOnR5N6pr7AsAjHsKvBu/xgSt6jeo2ykB88CRSprWnxZ8xso/UDQ
oPQ6fsUCeNTmcds8x4p45oorv87O6mdWEex6yNkq/8EV1zktevT3Lf7OuxhhvIivNwxAW4fZdhvN
3Dgp/BeaCPr3l84obJHuRyHh7AD3umRHr6usoDuHH9J5BEouvNXsJgzsiuCGSMzgoF/lLXm6bzkk
qCq62oNzeS9BLuWC/PQUmUeLUShEVhoGVAZmPfEH8x55DToZTzZhm1LsGDCJxOqaO9NV8vtd+fIS
Zq7Y5ITzoMl9WzN/9iWbXyKHz8ABtB9cg/OaB0yRdgZ7Ts3CnFu0cYi8JMjNnc6PkCaWrqzbUCSu
5A7r6TqEYj5fzVSuVpRbIRPgTN5JBeodu7Wkb2lzuU7I/Noo48ONETPerAEHTOc/T0dFRqK893ST
RfM0bIxpl7nyxCj9xkPpc5CRgKEylEsmqNm6JzlQ4ACcZMN/8IZdxA9PVfee73jhC5mmZUD8Gsgc
roQ2aRraHTVM37VddQYHZfWbKBuMO9Q8Z72nOFtQiDLhGkiDBWJ/TADeTQUKYzGqANLcD5oENQGT
lf04YJxKewL1kHt3KK3R124PBYwMxWqgC/r6Fm2xUuz83bOdqrSIdsqJ8MiN2mqDL8tJB6R9pm1k
BqUcKEFiM2AcKHpvoUCRpMMpPr256uawawtBiGisZIXG1t64iVq7GRd3PwXvMtTvgTNlgCJ0xobb
5rvA+d5t+m2JzONPxIPDmibMJSlFHXljfTHDfXzKdgXHJoDCG/nVlLpUnnhOL45A4myl7uoQz6Pt
Axi8DDxEads6sKwXAiPaEzyVS1XRFcvJh6jRGMxoxka0kWQSMSIHKUYNheWLgeeNUui8FbHkHYYG
WzQCOH02HVswDMM/EsGKClZ87AemX14rv3l2/LhiYZOAKaSIupiQFUGHfOOKSeRVPdhZKz/r8SlC
Dfhjq5d5TUm5zIg/VTAtsA9rbtWZ0xZHkvOJhe23LWlpQedHop3uqK6UwREaRhTu/0k5oxz/3fwV
6Vy+nbURhf7Y9nUOxcJu9d2JZftzMehQrcZc9qHr6iJenB3+gw61WfDB2rNP8sc4mvcI0XzSTHvf
Y2YLf+irUhe9fOxpvPBXwyGacWuUfw1yCXrT1foqaDkcdmd41C+HvnbZZRgWJLJegiN3drBVuTOf
sBCkPHiS8nytIr54FQwRhJUvLWrDSvrEULh0kPbod0tmsFLeJv2YmC1wtQYz8nPB5pVciB8DGY1n
cswkqDsfJpy90FJsXCRsRGJbGo9JsbCu46yM5yTT6aTRtJFASa9xy3eDybZCzwcnPFNPaoLU2HUi
Shv9KwTqc9Zxri+lMXQFf2HGVTvTbBykZS8ABIMVHJAwpfudyqGUWX7BoHS6CWqVJy5I+wLYKI6/
9Zw7YM1AdmsRcluvOo+2DYc1irDASB3e+xMMCBWdX9XclZT73osJ3m0xHUznVN1yf+n3/8F/Awhx
cdVhQI8HBtUQh2HdlCACEIVjQ6mjmJ4KnyGU1XkM1KUSGXUoX4ISfOQKbXutPjcC9TQC7j2zEXG8
zfc1c89NUQyz/45zTLuA+C9BB0iLtqVuK+LPiCMgyKA7GQEJOpnTGe5lG7lk6lK02G5yP5CP+rp3
KDjalc9W2yfYXChmwB/5rK5Fhiklo/LYhdPTrhwrOJOQe3aGg8ZnlvhHfWx1FBghEzsRxzXnNKIP
ST/eRk1wqnKM2GK7wd5sKI6PXaNYJTMFG8SeGpNkTZS4LD55QRblb/YguogovpRCfWFmEw0UqTQk
9jcGdcFZm8VwxZRrCkvjNasiiBIK34SuviUACHHXh4tgl3e9Uj4uIZ9jE+di4lWWcaZ8ssANMW4Z
ekvkeBXQEFnUbit0tC1N9tJy/9pkvghXDlcNnBfUIAryiaGq6Wj8ok8Rp9luJ/zh/B+sIyHNLxX8
Zm4dAOHJQrVT8PT9Alh/25KTwHmqrosQfifzrpMwgo62Ol9Im96tVcrpfI8XP/MhASHcEk9lKVwG
lOAQZnyYbi0k5pxlBzC64HJhbZjxROYoVCxWEEH0DryeW5tOXd31nq+1bGw4SyCBv0IySt4BZxqa
1xeCK03QoojZmvgUW7SzOnFqevq7A7LSXiYmLSY3eT1j1BUhzImVMMLCQtNgkE15EO3OIwre7jtb
Sv+PEWmkOXCPrpA2awM751gYambk/r7DI68PgPUmiUkabHXfyK7dzkLx2DmggE8bYQvp7Ca/e+Uh
yDJAw6JDUoUwhabLlb3lnRachddZ16NGxNQx4T+5Uvh+vdA+3s9vwmO/9/ys4bI/gH1IAFYOju9l
lJfOd+IE5PlOlt3hlygH/wH39lzy8ZWq+awynnLmulSEZyp0tx/rOyu8MzwMhCUISXW0x50RtIjc
+CXXey8zj66x5t5b6oBONX+R30uX/s6HmtX5ZbkWBbqHmw7OXK0+s6axZLTxndn4YJMIB43rUsPj
m/o7s7u00teVimE1kmsgMLP/pZPeBP8lFLE416aOKKBCvOulYuNy2Bckgk2QRAIzsaxEtzrCklNb
sNbX/pC+OR3PeAEDMaecp5Mdq9vyn9oDeOki1Ga8AYxZ1aqdn2+12GE6BQa5ni5BT+OxugW3/SVn
gGpew/qOERNjV6h7ZYTHk+K/FZOOLStvfwGOYIdvxFY8LGdtPY+SiBcDWrb/pFDBQdOEoow2B8VE
E94zHay+IOos06Q/7C+TqythyAMjQhU0VzXxlwhHQoh+Gdaw36WdbVnbrQUNwVl1fwqEEj0iUfJj
6Jk8e09bOFIHEGfy1k4itdFCrbFvynbO++GkCsL7UBU8b8bCBiD8StMYavelT9z45mJ0TPMY0r/T
Fdfta6B1qUAR0afCUWdfgdF2RuSrJA0UZjy4PA+EYxUnThx2BiD8C4Zds9HKyp8entMUg6iFGqhG
b/BAazdV3FSTaDstPL0F0LAHTi7ZJ0WxsgAAlAikhE9CtIMnfg500LiR3PF5C+8UjNxqMhumNcyR
VJP/gv7ZXZPQLQL36vh0eV8Go7wZNJrwkHj4euTLQXdLHS3cMtChOFqNPFNJICMxrnTmiEAlSsRZ
S2LVejdWQnQgQ+bVf00VUJ1QrSPyGbQOj1flJbSeNk/VM24UJFxfJbb4ODq4pz5y1Ujma0+KJ37O
sXBJE0H1T8HJewUgh+Kg4qKf1JBTo2zjraejpFoHK2qMj6KFfekhEbhWJQPNNrzVjZ2IVhSYLcJL
pDWgJhQ6U6jSqp2E6xJkPrjqTHpUJaCxdmJ/B+idHHUnPpFB00ooST3xUwe0yLdJ6fwsyBb+QmZ6
3XixWb55kJW7v0TafBSvmt3YRUgq13AqWSkWwhWPNQUfzU/oCjJ/nUKgWKnzHxQ+qxtNUjjdfGTZ
zw7Bpa3wvIJ/1b2Y0G7Fl4ZDVud2cLOmyNUNpMUnqnTcSvvBAUz9/iItJCDEtzPnL+O5muLTU/Br
UQd52JNLK4JCyGiCwVKUha44KmekAGDCqBmQULVyawtWQB5ResjUgFSxszK3amY0ueuqk+A6frUY
ilIViIqtL3R3ZYsLpXU5DMkO2pLAABMXlXKdB2hsKANinoavGt9PQsz3kQ/1GMY0kw6sXtlzA5+f
5iBXEysqpiHBx/eluRooTMFHKdO82R/ROqgjJfyKkY4lfBkqTYXx63ko24xA0g1aNjUNvICKlCKW
IpsIY081p3yECQFI9E7ZkpeS6XPzk6pf3DW0SZntpcflSaUTyZDwxN9+rzTdp+Uuqf9pLl9IJ10B
bPEk1Y05bAEcbm9scSW9FG6Bz/UyL3HPMyhJplj3si87FnfzfHY7sssTfvzBVdj1WPB/A04Tgpsp
idqZ6f8t7/c3mUQHSJxMqstDkku72Hcop6eYLUrvSLWbXEYlSaF321vLbnT52uSrdStBpw9OT2pS
rUPxoi/94VWHeggGMtFAdgXOFBOAHJKa5KQJl98O1FL/JNvOkseLRvPxZeOo2Q5T7Sr3iYAlrO5y
+xJ2if2Y9sqxr/0595FH8n8uc+ZO+tYRrQCwWMPX/ymkM9D8GsR5qG9mArQE4076bz5AKxIFqXfl
TfIArz1oiGdffZ2Oo5ACbFCikiUl+QuK0qJSg+7yqQiSAQ96vxeFTZLlDDW9RuDTbuncoj2+VdaP
ze56duIQw9CmGkNenSz5Sr0ArGqYQfzpOyR6h0dgnmKICAJb9pVCCAyViCwmVjdwigPse0cXcgyK
mqkmDpmcfSs53/1aPbJoO0hTJLir+gM9owncTCZGtYkbadmYbYB7sVrJdVOu9Bzv95wdIn7a7MTR
PYx5sj6TSLTAGb1et2Xkn5oCroh5VMQ+RE/QxRwx9BtFxLOAUdhN0U0/m2CV2ztf4QybhuuK14jV
4Iids+dP9vQjDMul4fWasfmhoizxPCm3iS69EqmUiEeB82CT/m7aFP/eG58xBddN+0D3KGGVgenx
xSN57/T5o7Fefigg4PsFW9qpAakv0BddJyQ/73GZT8O6DOj+Gt5cFBzNgStxmh08nDIdk7nJJ5XK
CRfq81RjmpnGUf91TzNSBXnWL/ctfWhqL+w/hU7Po0AUWePEWPVWnzE7mYmt7JJSxu9qS0BxLTEX
9/f4d8xw8LPrZvBkvhAs30gr7bmx/ZDo7Zph3PJFrJhgoVw+Ah+ajMpyH4V0OevzPVMPGvO+YIfB
PjaK0TbAa7xf3OIDRrBRlV4+3k35MfBaEIH6oE0Xmk1ygepGC1w6NXBzLqbEyXXSAjCzm2bKWt/J
7QvfJvp+1jZdY7VXEwh5Y3DzpBiERrIxLi2VLGGdtBRFdTEcks7oY9SUPcofZ8n5x/ZsVTrekJud
LETBV3Ta8TIq6CcnHVDuOieA0A2/NHIJ0F9TvHJ/viuRWrgBdfXxBMGhHdKVqE73ov/Eo9HCNPby
xpLsdPPAhd+dkrLz6apkhITFeSwSjgdRsZVk0Ko2hM/bDeVnhDn2gd+cIR2yffaHkQ9uCxYMGgmw
q2B2GdDJ1kuv3PmfEWeZ5zAoAI6j26R4+HoPDZ6gXDG+7q6/HaHmmPbNvZWiBG9vwZWeHRc1In2B
qxZipgO/wZwXH35uwEMBWjd0c962+3OMmuCjWA1p2OIFAXOfAovnW1rB8re2whQVxCHmfvs/uzfR
HF60BzUzpcGDZs1FEARW+FfCiVyV4ADt3we1ZQ9rhXsIbYHRcyaW2fPqekBkr1HFioXwALq0AnFq
fgrjtt3bOCmhcvVqd4O+BdJErhidPV0yEhbMey8zBIPLyTLwBE7eBYT698ZckexPSh8tXL8luXgj
CSPVrZHJ91/EIGHGAHkjivx2m1nv/JPXXHWAVI6WBdg1bfLUXgpZ5nAHkkpsnGCpEc15jykDqFp9
G5QhlWxk5hKpHDyWS/3kQb6YK7okJjykavu36tj3r08cTKdFd2totMjNrxiWkuawSX2ZwtoMCTd5
zHZIZ49oYSGwrUBwvtSO5nE3dCNXAARbz0IKyU4Lh7MdgeF/Gbinw7silRCzGcH8diojyfRWjQ+W
p3NKG7aWgux73sx/RuNajcJI6QijkD3cTVQ4Kd3pkAPmVBXBAjomPtZR60BY9zdn0escTaHUYzwD
zH0a8CZdbEmstWWqQQfiSBh5/7CVokz+y+9KYJpYDEWvF0HCfbQaWuq/exsrv4/AnN2S1ZTta/70
oIeLA6Qf0BgPyUrazg3hEt3tQWHLw1nrrxjsgp1A7iK+4pDg0z795lYsYskIrpTufJWSQ5JFdiPC
FiaDjsn3k6i7jtzvcDqy4go1XJba0Tb55N0RVUczXQlc8wVZM3kjwh0KFyZSl1gJPy5AuxOwQ6cI
X6HXiXNuJ5Y+QXtmRbizISySaOyROTZXvakCRy+oTzempoBCErMZBmiyLxYw41Bip4LVKA4s65Gf
g6u8SXNZN7okiJAyImm1VqcDrjj2lMpvRWb7cSEWGS/6L7XHo4R8c8FqMDSgPijaRuMvch4hw4j+
jQULGSdy/rm0Lygkx3q5U+jV2deWgC4qH5V5seOyJn+lj47xErWsRqwtaqkAtKNSo8xqKUpeKAmi
w2fVCWL+bAGRZR5gq0lDHuSygMmWoBI1lFe7AkuNRudT/A1w85Zi09T2hIJNgbOL7bAF7ANqlJd2
bfVyyRFcu1Y2Z6HETjyvykrq9/C9c51JK/xNWOJTNbuQgMVC4RBxfNqOIpWwHo0OQSHJ8a+GkFOP
/xP0dayTXFsQbE4tsHwuG+X0HE9jg8+m5k5ixeI5/iT7Hq2HkerGtqXZeJGce8gP1zvgLhzaH0km
SBOzXqYkEgpm9LahB169DaYOzXS3O0NnVryRdSCuq9xoP6PARnaMcEDyhqlPaA211bIS7rGhVZ8+
rO4QwtdEnFc8vEWZFMzWUaJ9JsmpJPvHhqL+T851u3K4hiygqrz/qe5UnIvyUrTZb2OuNwBubhCI
3LhHahAoe1ECNum6HSMjYwdozcmXXRuWtjd0CMb8KDxN+qmMBaB6WRQcEx9gJ6kARZ5EKq+KC1W7
mADBG2KLDTlBw/JsjKVaCF9qrqbR2OV7jKBf/FkwzCpN96pUrUWWd2Tr26VNpdHxs198x5Ye1KRl
+3lXu2w8QQUnu9pIJdSat0FOk0JeHJxxhx5ygdP0l8XXX6UWKbZM3VkZJ+LxbggRsBp9sWTKJQff
lwzWyAMlu3XOb7K2rJ9Vi+Y8KRFEJRp4SobzgAMfrJJMA0ciMW0G/SWoz6S+Amy+8GBuebXJnXaB
GGA1e2/ZeQE7yMhR/1hAL0PhxJS1Hoo8IRcHUfeV839bAae88kTo2aEei026qDF0DFoZofvkOKd0
EsEJNksXhW7X6fEyjl63NGKeXYdB4HgEMZ0eOTU1cpun7jCWH1sSlfzlglDpqyL4slJXBc7r0qDx
XvAW3BIVwEjht+ClfQ5caurCD1L9qZrAG3rJl+rumiSb4a/rhnXusPZlHPMV2NAoTVZtE+8GSv2/
/mk3VYkuS1WU/8LhlStjqMzwX3aDz1qlqCsoAtnSDcJpulebQMDnioRY0CnUpiq2J7lcg96CHZEw
F2Jv/vHpNN9BZEQEMcj3Yud0ksJB6nI7eI4UL0FMi+zPXzuPRpjJL63mGR4wPujNeok/8Om3Myom
ORhEqhXelAiY5MzfczAKKhTOfcWrmIeq7f1Y4P7ix5gkxenNbPVzxl7taimBGKr3Ok2o257xJYfE
EvfY1/CsfWjyYf8s7ZLz4lWbXM8W90Mbi/nlL63wiajvtVR6u8kC5Qtt1U8rBs705bZj438SHCq9
hxqNP11JOUD76xwdq4JWMG7CQZJCCCxWDneHErA/MRZjOULS7y+8tvDBy7Yu1gHFyOIOtHeXt8lA
iXnjjW9OecibJiLIgPkFqi6BK6iNG42u3800ZLj+ro+uR0Tqp3X7Vjb111H9aoYFO0E86TfNxFrs
WiPqjmlLQPCVc2r+q/40MXG2IPaMskQMjQp0zvo9rmejMfscFVJ6zIcNTUfd0iLYLCu7NTqotaoX
3G2Wrly819Kxdsma4QxJcJlyNaEdfnIeOax9GXRxgbf22xZajy5xYmWf6oVMW+/vK5lC6ICd/9MS
orzWf4jG1CGYJz9vk2OJwMAk1q/Pd4GQWX9TZnWil/aueH7kCB4113WqoxNOvsZY93XgbeL33yiR
tuzpneEH2Hx/+3Yik5I7im2v695eUNRsxDTuNDqFqkL34Yg6AuphATkJcHRUpWXo8jGSlw17uEp9
zFj5E5TT5xSKoMKlChZKaQGJQlUTPE3URB5M2Wkr9TQG5bRn4/dRFSnOGi3pBfPahAzDN3Wicaun
MRXtu14SEmqPTPzFI/4ISU61sSJqWJl/e2A1xfE88HDP05Cnem5zHRuidCRXJme10/1CvVycsbjT
2t328qJfCTBtbqEDWGBsHlCqAIUaSCtzriJw11ZvgjZ6Rp3/tLSHPODaJBMXh4sSRpvG9UDguxDt
+oizaQ2OC4KnZi7bI2AMgPTBSyINNJT78dmIASOZZCQHibcFm0P3Y74XMBdodMWtkGMbMlovXXNS
GD77aJxp6ev/5/70Z7W61+bNwvZuFGsmFtEsDdycZ/jcBdpS8/F9cNjLxiIi7ZM1G9RyknDs1eSB
3GX2NA1X0QQC14byy3uZAt5i81pHIEQ2pYFRY6l+E7yOPnTeiMhpXIlD1SIC30Ir/ZGvwwX7DR5+
Lc1L2By1dhg3JPiyOBURXBABH27np/y1QgxaKHpObAYSmbME21CWjzuFdk5J7lLL0mlHwP9SVJW2
XSsjKq18UyP8Au1oR9yfAMWQUxKB6nI58Z3WFSlNx7wCsy7LoNOFMz340WDUpaMvYbksdan7Ee6E
EK+UIFoT4ljg1g3vhSbyRrIUBZm6rFxVmn6JWLJgmXUqkasPKeos7F2i3mF+mr4cLrCJ6XPeEk61
n40wAYLAg4ANqc68jRNs7uOP5lvUJlmFT1SqxGDXhhx7RBd9eGLFmkdszbGUDGP0UBrvqHA5p5ZC
PAcmwkGto7cp4jq8BwLpKhK7zdd/8LwxS74p1AbcGT2foFfMtYMbSNwgAhswKn3kI0cgmnA3Up2S
W4W77VghTIznSOXoSqaT3c9rvvuVd569XouETfvCT71LjdHFTRXf4HHeee8UXtwEk3HEwq9VSKUW
OacMqmVYy5hH+ht9gpbEadI/xghrbUyXag2HnJgeXzh0h4fccOcOloQeWTkij/j8KIkF6EvgxMZP
Cgw942oDsA6J9gryd6Q9x9DG2U1JjglgvOr0HyI550vd5qmiTnEvY0qHq8KqfensjmhENHP9IDkh
TzE7eVSKFL7Fxar0dKpw+plWd+qvyjop57xu/lNsy5d00uY3aF3MOGlas271+TuQTzZy/8rQsayH
ZMcpvEjKJ5fxUQGToz+wR0HOmBMnfbFKkPPfC6uXWwF5GMNAqZG3cW8KUX2WI2y32WqKHXpujGTa
VE57W23vBAdXq+tWCG9H+Ln4MohDLiQ29yprL79qhu68x0gw48GKWfVBnjW6/2IwezZXovzvRZHK
1GQDQdN6ZwwRemveXlwILVtyA1YKhUaENY5o7/NHYzKdjQNjVKO05jin19wRwRTinywTYZvOdxry
z68u9qAsHPO4U5eh3ePEGjD+0eTXQpyr/QnfqmkLUW2DcqVkipxP5vy7XJltEW63Bi+M+h8JT+Rl
9okzJMqG373Z0SxFtB4U8iryI50lQ5DRDPH7nmW7TX+uKetEuhzgC0RcjQknUpR5abb2a7XFwKBR
1kJQvyyfIMRUTC0382Fs3U4EEKbOPaQYl8W5gsWsqq+Dt3vus8Rje40NiekKhCWW97HrTDO08SFv
2OLlw/v7kyEoCBxLA6JhP6jJPvIac+Oxo7GmuMrlH3dOalWKrStfxUe7LiwMqVfPYLHPt9CiWWhf
RkrJ8Xe5H9NiqZvL3nEcZk4lMjmAqNGECe6vzZFlyKzH9T2bsEWGKAtR6hE+rSCcn7Uv3Y/62+F+
Po5jO4hKKmWmYRBFR6yiRlfX7VeVnzpwAToaUELEJ3+HaNkv0G6DLy/g1rpcJ3LdPXjiqpEgN6w5
Udq/mU3oVvGN2b810iVWa9cJeS7m+Xr0yFSYHJydvfZxqY7B1g8dah1b4BQFAw+MzwFkAa0yCvlJ
G52YrKln+frQXV5gs7hhvVNAEnEggvUDChf6rifVq1FLHFdYE2/3RGhYXVb6M/LpONzBxg43hyR9
i1DcXvVs+n+aSDkFqHLFLlr2sK907NUq7WXBgNoU9xTLQC78jnuyk/e+g4dhy8+QUnXgSWD5y0zQ
AWKPj4S8iOPles8La2bDmHaW08EDlCfB/iYdKkSP8wYG5GAsKMCZA6KlGrKy6FHAn9ye1iCW7qP3
2v4Zbw94JITAVTWbP8z/g23fPRcequWHWz0C4QcMFQXb3luXfgqr0qstFJim7fbvi5daOpt/3zn3
r844MnfT0PmhnQUgL2/hkM0QC0m+O5xwYKUIMB4R+oZmhbGhNmZs2T/LNGUbC19blH3DsHA0BYVu
i2rIZRWahZqb7+4J7Jqg4YhvknbO+AW5lsuhfIKQiavTcR+eCLliZOZXr5Vlp29pQUtrtubKcBfo
mCQqJ4zsHAgcBYMiSGrOo9bKupK/4g++1zuO43S/f6ZNflLpm+b5dwxPC2Wwml5CvU5p7AcKE501
5v5itcjtq8C6+J+Y4sla566OLOzzlPhhABLVOs+GzcyCd4FGwWviV7UrAtVp19wUY2/O1AjubwqG
E62O11hWjfAK1InEwJq3eIWmk0sFLXwlrAnkAo0p73sPLJPn1un+1JfzyURJh8TNQcd8FJRZWOza
FbRnaS+o5C+NzMz7IbZX4jlD4cc4dGf9HNMw3vzFWHuThIA1M2DS5oJmDimenWifF8+Hb9QsUkPL
QJKB6zmS+eNptuY9p22R+wNBe6JOMzX7rzQ2i1hr9xT6ihRvSqqe3+vc6+ILiu8cp+8gokxx2YIp
LKPUN53eFkf+0fn/rkP+jOewh4453EKis1cA6YMInayjzTaiW9kvQq0C5Ns65uVGVxKANPPMwbYu
fanodH2pAsJsxieKyS+jvYlCfSyaabyJqBW0QsibV2rjvcwA9sDbQRLayQO1tpfrmtc/Jpz+kH4Y
6DMmJfBsbN2Cg0SMQP7v+Ud7Z17eaLzsrdAVKIxoM9m2WqTJsz1/Db2kF46kwdL7jF/s0FOYOtlw
V0FRJ88jOD1Q5Gnl/5zd6eJ2CJQgZGKKX4QpOAz7Y0TtKaIK04Y0SwhgX99fkQI6P2BxzaK3JPo+
ZN0I0Z3yeUZ7MoCmF4hmIlPYuiYAJt8iODG1CdnXX1DNhDpsosX4fXfEOa60b7HRYrxknDNTWnhM
F1Wb898KtsYHqlqXi7OIl4BILT0NRpCECrIZtFf++n1t0iU3xEds1oaB0i1H+wWn+2AnDJXfVkCY
/u0G62pLgx/va2c1/V+B8ieXT6J0eMAMLIcAeFCYBgp8vqJlgTEKsMCQxBVH5R6MyZO7S0cpCfhd
phJMQDn3hmLeE175kSS9scBxyganfO6bTgBijEow06YeP/pA0mfEFIFVUwrxe6EdDCtPImM8BCBJ
FmG5CM2KFGTWdIKjO27osD+6qBDob5fFrDr5b6Pcw6T9rbIGqbmOIz6qWlz85Qxgtz8Eqw9JgzUz
UBNM5Py2g0vGEGGdJhoTxmaqLQxMw3yzDVsga6kznPoiI5mxXRCrbo2DnOo0/4XGlM45c1hq9zol
p0DZrmikhXOAV1EnPoENlJajRWLmBP6Ae/vv2tRGRAfaPrH22ksAuSCwlULC0TszH50Y/kcJl8dL
QFzof+VJs8Lwcrcx4IBF5MUU7PBBN33uphjiD+A4gJJFtziuC9WQBDelyTUHuKPpAFMGkGomiUIG
gwqwTUvLKxTOfME9jzaWy/4ImFRzPcvwqAvlzWnk1vtmvXt9EuD6S4uw9ZFwKJd2NcdCPkYGwFjL
HunLe7mwc0nY+eywJHFY77SlqTtQaWniDNmIhebUn5d15tkhMO6Sn/IxylwrTSpQAISSjnguRX0P
a1wZkOQ2DQiNBvUZPuR6zM/YR4R6AvoXbDnGuonT3LzIJ+WIGW8P7ZTcK05ersa939gyWTw81Pu1
VVgVw5zE7KMwX3mAIbsf1Oykq++39RTcQ6791IeR+++7NMJ21qB2qcpQFiy4nJ6KqCMok8pM9bCr
i0kS4CfUuHOadQkQPAHxeZqGFIz5cWypL6B5W3QC9RTB4r4ZAcaFfLQQJkBs3UEM8CSRtMKrSz2U
HCCSVhIu4rNo4pPAp5F6JYrbe+2/GuvHMh/Rm31hc/sVtqHYc0sAewzX+ulfs8PWYpsBi906eho6
vUh9xKDKrRzZceBfIOyXaa7IMDJYaquphjhFZIFPeuu1Jm4vTaPEOi9I7YdGQBAwUGJc3KFwysoW
n6m0+VoKCwU9exbcLKqjoduS5K9OmTVy95DQx5sgO22UBjQvSsWISPni0uRFp6Xr4bUtjl+3Cb8J
UW7cJVLc/lUjNoc9tobxSTUaP9UgN0UmxoleHNBSuXjP7j6B//JHtndMJR/8JXjvw1AAw9qsG/sD
WAE8Icg5IAyMqijYglTa12SVcVBWUZmG1sFLQe0qnx/Ku9qrbIkRJIdAoLsBAiT7ZvRRCCMPiSYO
aMCVQLMzdEKytg6VWq8GRY3M7oBZHpIisPDHA+i1xuU+WTQWRYdg+aayFM7Cu0jfp8LnlIIgoc6U
b/RNe/wffoNU1dqz0LJWopnFHfvs0NUkKzwJ1lRqB0PhqIs0lLFG3073i3DwMWNuMYIYF3XknctN
GriQlzuj7Y1PdWKLno0cekULZractqFmD+k8wNbM0YVyh456Nj+Fe/Ukt2qMQXUwmycuXcl2k412
qQWO5Owd7RMnfhVnzi5tOx3xi3QORfujDDMrrzxKmljGz9hWbxBn4o5qE3Bb4QuMoX5lwj/omt16
Y14ME7JnrRomXzY6koARGGQDV7VJvD6zu43VygbovUy7C+ALaMJDzIbM8Bnkun/vuM+QiahMnv0M
JJP9ol/PMJgg56g5bwevFr1uKVDrYWjxda5ywzTejRfl/5m0NTB6bts5Fj1Dj4I7DkXxNnH9b40i
zk2721wsodvFuWu7t9TvLloVS7WolQJ2dy2JsDG38BJ4gqnGfT0C0suAeqfgLMpFptxd2c4JgNf0
myS+54l53+AzwlTvFs/LMkoMPOBqDBBmbk97tbVUaw5UxHIzNyeTruAUZlp35pmnTnnUEqFL1WvA
xji0xnUM14RTxLmOqqOvpoqJectxVaeICSvutP8zKRQlnrwdqzRhXsW+4Fc30pQ07/jGJiWbR76+
maS78RnzWWovGv9sOoiImXAZwP6jHmVjTAWrDF3gJtK80CddV8dymnyfGr+bJBZZLg5ctVEHuSHe
YhKvorOf3KigF7+rt+fBnVX2T0zHkUWPBSOeJCRW6o55PVZt3cdSmV1h8Xr0yOOvS8L+B/VzuW34
qPK40J+BFBDSuaLk+GAsl7CJOG36UlC71wAkyzFWoKkr3KNidBalvsS8gxZj5BY+jQLXI71K7F/j
8Dccbytq68xP6CnWXPW2IICeQvZUhs5zs+zYjgTlZS0GMbTSSCXW/L9XQz+R2pQ23RhiQAaBTwBD
Qwviz07b2GIFKoLp0vEhXSMyQRPzy5C3OBb6ma2HH9yOgp5hbEX/GqO39peALLDIVvjgVLJM+GTq
2c64Y6sRtCMd1KsSUu6eG6TzeVMsLACS8S4+sungRlAhQfxib9xAki2+1NPkWRWau6V3obekuwc9
z3UrlcxZm0x2/7WUfqpPPSvCRrK5QlJW6VId9EjeIbkR0wWbukz6sRDcMMSYJjRxJYEnOpmh6YqY
6I9gQFyPZ60DHAiry1jT1cV92kh8RzIb6C/9HSXfumtdc0NeAZRmS6+1qZNQDllAfYp3PXn2SS45
CEBCGO2HumiXfbtEFTqARHgvkEaQI9pGFh3jIHl2EFZZvTC6bJ8nht4r52o2YH378aVnI1js5ikT
Jehmi64DCiPkyEjVvQaXdeNlhoelssLKBtm4GWQAeY+KpTabweFW/7wXeG8xqveY77OAKjvjGByE
E1PTpxGq1WjagbcMNKXoyKnSVM2tpT0W4gOjXVf7tnKf9kOaoFlnHtT0pVD07bzvPDrxc/q6uTMO
kiFwpaKJJkS+15Ygf7cZrmu7uxGxk+8809GZjyqQJ2LHInpk4KGLHGMj8XMRvUBFeVgpbcxI/gSD
5/P2Lps3r4GOUpTZgDmeHL83TbAIbOZmyQZ0QA+qALP1KEF1nSWIOdy+LW+r4+XvJtLflds8vO6p
wliDtDcZEsv2EKe5we4tRPH8z/e5WYneekhzmMn4j32YoAuSchsIKTrcPBCP12qtoBXx9SOSzp6F
dbFC6TACEhrB3XCEDbF6tJTJQ7mWow5PE3aS8a7Pgv+whVtiexGIrCwxah3WHIjDHESNIo06XrsM
62ibU1mE+ZLZm8FZLpG6GaZUMRcGNtUXImfnco6+KY7o4vdkqOSXEd5efjZTHZeuvm4YRoce4RFN
L/3OjbJcQVnBcGu9rNGjMsqUUOzw4rzg6xKjX5QqsiLh6mRUdhxsi3GW0GMROet/4qFKD8aPS5Gg
M2fsmTIYSvYCHr+/SqouWtB5OL0otEzysY/IsLcNANprtz9CZhD/yVNlzoS5EkGuh8BEoaB6aL0A
rsHu3SQmfV7d/sbAmQA53PaiLIFkuugLvVMXlKuEkmKRDIjc3YIKOs0JwRcnU75x75qffkM0x6Na
vRezPRxpuRBaxi6CLfwUjQH4L1n2iQ8fMpreef150WeOtrzUVJezkJUv4/kJmZ9wKksHDNyXHKdt
g5473ra/tkgrghpm3qGekDgzcLuYhlmdtolu1lgMe2LFJyWquTEgtjqZMVlYAbpxbt/dCpTv/xNe
oPiCGU2RAHsg+5a2kguoIb5n8TPbSEhHxWwQGLsSPB0E0CDcUobKm7NhWTx/yXG2uCP8ugvj2RQG
u1YwtHU3Cl2pIjd/hpaJZeepXAX6zyGRM4klqqfZt2CXGZKx7pCR8V/RJ+wzwdA3GO9Fh7KaC1iZ
9uMykBD2k3eYNEbQcMBv4gCNmzz5ivLokvj5Yvnf8ykiPsfbC+cU8RgO9vjbqHq7hAEAPFlvfwip
xuxotV0MPdgcxvGqv+/JVgE044Qes4a0pDZEsUGK50Luf5V6laG32SZ7FAJfEQsYbbhwB2iN6Xnd
BRce8g/DzbY3r8NUshEC8JPUnArV3RnNiiCG0KdClNW5QgM4FnE4nuygwszf9ZQTGvG5fetVaVOi
UOwzDqaw7gwMH0Uzg4ReUCSG2+O2tioNiUb+JQdMrsqE8NceWIhspVPvA0Ft6k0MFzfGRrCrMOUz
pu8C/fd2lKjk2ETklm0LfeEaMds/k7FbFvCcB2GK0CW2MNWi1LtKVBU6VjM5bC59z8cLpxF8bK+O
Z79QHRZU8A/Mp6SL+XCeC+RvHXpcoCKEWMpjkZqzoe0/4XszzWR4RJjnmDnD1kEYBk3srVdNlCBI
08Dx2puJHj6eV7OnwnvMYkynkWfhkF1fFskEPUBlaIjDUb2NLyssjvvfuiyA73BUN4DKOOSiRfk2
7D/Fv4eSxowGuSeIGm5xMbugQeYPsZlsS4l7QexX3Ui2KhHzWP3DvDFyTLbaE4X0cjRDDZV52dbK
DK+W4jNSMsjevysoJi0s4NvTZ++qj5DS8P7JQfINqVtWVOopVd5MmvNw44gwri4SzudP7sJPGVZv
Ij8ywGNIXIf3ks2fVe4KVx6nRQkgXbjxCfZ+9YhemzKS/v/q+ivE9GXRzHINJmDcOBx9h5g+yTw+
9Hdm3xsWp7QgNNI6fSWQhRAAnbQ/WjshaLukwRIpEdLCfeJdxVT9uRaxmunwuI4qqvYH0WJvxt/g
4w0CTgN3bJI8JNhfaWaHIiDdr+s1EdfyJFOUJmcYkDtSh1culUCxXvWDgmW8aBKwNRsOA84usgt3
vysqkzfPtTl1rExVZfWd0W5OW722NDZGYmzscgG8NZulSQo+uR5cwy1VfGbGrS4GEYlqSg0PnEPN
QkjzFyqn3dGVLBayJCEWih7unanTOFShlAC7uLbiQXk1d4l19kafd3jJ3v8SIoj/hx0sc3WO/UFR
R/7bv3U+9tJ46drgjg0hIu+fbMtiFYC527EUo88M92qoEDPKam2deGFjgRVySFV2Whq+Ff6TjAIr
1YOSUzqKOb+iYcjrxk5quGamjeOlZecWv/dyqGF7Zg8j5HULqXHA9bheV/UHG7vC1N70SeSVGZqW
1ubS6CMdWErrzE+SW18AcmNiWkBVvhG83T1DJPXkwnDDtnokq7z/snB3EBpD0EZwueDZkcaEEoN4
x2XISW/SMekG1/QCrYU87mYUP3sW7/OO3ZqcvmwgHE8l/AUf7uUgTeCcMp77QhOEE3PfPMJI2UYy
Ooz25cJz8hH/MBHYjEVxZ0LgauOccreKRopqaee9lp01b/PAtd2ymw6SXgnJqEExepTzsXYiRIT9
LJQBxebHcudJl6eGzD6eJQoXEUYjjrWNsGPo2TB2/HKX+W/L0ZwX/z8eYUB5M6L+dJBeC0hc+jL4
44mkzCH5Ogeyakyaejr1gvcvYvK2hqZNJKEfNdChojLNcxfdMhSW9cYGKiFSGHHV4q8D17sc58gl
jfXKxKvNOhpHF3983tVk3qG0uynCkYnta6M8Vw+mxPheSVNKCLEJQGRWyw25+W6HEabcwxIybOMJ
9XXTJVRdlhtE+s/LZqO2xc0/T2rkE7rSTSAbSK9WQlwZul5VTTJB4WbkCFXgLSH7Np2+JqVpCROf
IRz9Dnk94lcCbx2y6WwvPQhPXnhOajfdL0vUBgkPlWaAfL7+ZcX49UQZ86nEO6peMlHsgIE96jv5
AG4Xj77BxqTCqTatPbT6IbPQIqRtVbPzwEI/NTfYLQw/0wXRa12hyE80WlpKdFH4oDs4GR3OgG4B
72ge+9xRXRVtcCJ5mSD92uBSB9NIePT+AtaccQnRc7osIr4HQDvTqR8FwYdMNwKkzUBcyXaNLZUk
5tNSVmnjAeaftp4lu2BwYTjmn5rZOOfZtfvECjijc8iduIZopjfvxGb/yFMl/T41vaZFsmRmhy/X
BqjzvAOV/Ns1ND3YA00Ww/h9WNqy7HrejGmv3rzOOMBTKk9j2KMKXfDwYUkdXQo/Ffw0+aLWtVzh
ddlZQSGbghckajoYUS0Pftpwq4zKLm9fYtEPosSeHT//ijI54GXBsfnO3S/4gUmswW/mBtQjkuuA
0ag+WwciGRTLkMuTp2yp4gN/0PNHZVhmVOv77XRwtts8iHPPyANlyGEZ39nxXH4GBCAzTO71N8qQ
idKWdQ/vDslWXVlZj7ikMPWufVgd3JpgQVwuz4yhu8jcVwfG06ldpDbluL7KctndqpKFdGok8x07
avaDhLZ9mgbZ291y134AUsWsPujuovk9oM9lqPfs1z9AJo2q+wB20OSDmKyAzn1l8LnCr7tGUAQN
pkdsabFr9RbpHlQQfsJm4MqXzdihCiY0G7mHOj52ZR0tVWK9UsPiWyUBTCynsQ4S33hviABu0JpN
WttnihQcZ4URXaar6pMtTiG5HyHXWWJDDEdsbpnWQTFFZ2IbcCNQ6go74kvdP7ySbOOI1pKfrynT
hDODqGcuzxmdDS74x/HtT05yjNfDcHruHm4gSka08AgtBvcbTHrJgcP4pplkq4FysUFz80DCtTI5
JMem9e3E06GFP1R6N4hyZSLvRjByMxPAeAkin4dj9fl0JHT969C2Lr/+K7B0jetxBHth/5382UAl
mR1QStZcBH6UaJa0IDHnA2hmO1HHfFV9K9wRf3O1BXzMIMIeIhXeDKNeWGVY2W7phRVO8IFOUw2c
DcAx+LTfYkdR0z5gNM1r0w7pAuylOF0SxQXJLEGJ3VSmrlZFjkxB7US1jmYV5+v0p3/QqTFkwpak
NdAyJfpq20Af7q+fJzhf/AvIw/M8ZqSHxR3EhenroP3pUuk1oRcZAz2WH6ALQAySGdllW0iCW2NS
AZ9sydnAEGpxrFg0uyvsfgT2fBbXgw8tRatrlNMFyP4XhKfE/HLdW8AAfEJRsjAdinI5jks59f1+
3+uneY1E8DiyBVvyTxFVACuyYamPzpLeW8YIxCz1rGnUaza0W8FqAvoVqY1Ep32Cfc4vT+mAZkTa
6Ewoq8VWgN96mDytNUDQ8TmmX5E3HT2mQo2rcGjr1cHjkIefw4xkuWZ7kU3Kr8NIgOtkffNcvY+O
OEbAGbGCrtNJjTILAsIhOSsjk09yhQGOr9R6xDN9YcGmymhdRZPzUGzxzogNcDRIQ19icjYGzWAH
tEexRNNCL6Zw/NqwaxOO/xu1hrCO1wtsUVuES+BNGYP7TuQ0bKPE/PrIzGLLreupQoOxdwtqIEdX
bELGvxwwxhQa9rqbnTLWja81QjSR8is+bPcoBfsJBlnvrHMRd21emVZQSv6C2BF0aBvLGvaPTqaM
mWXMysHxCwGzqPvyiJ9S6hmlzzrVFztY2zaWlZeV/kl7iuSicy4bUNK/8bZdx2FWDfrkkUwCuF67
rqV772IHSdz8cMP/gmt3a/cqy1bbDr4unOnPhCdB7Zj38D62vqEnT21YFyDkX4e82kT2xGJK0m4+
sK/ial1WLckgLvZKy6WYw8SQSaClh5onXKdVtJXbA34fEM70gf9XK8JedDeyzKUW3/ib96W5zvHs
YFRIc383uiSNGis2sFVWqDTEfa/XaEqcnOa1bnGu5sccBB92QsdbaK/jqbD1Q5DeP+HG6vxkoNYM
8zqDguik4SBnYSHaoljVJ5XQ3Hxk/fNug/h/xQhyL9xtOJ29WY5X8qlubvVcH/2HdaIF9Z9tLnK5
x4s9ycfv0tqDig4wShs4naxF+rz9gbhkFjA0y33h2MerBk/sO7eehCTXoNVT2GiIINCsgWFRsegS
6AQDykIYkhrBW3o21QDQTYxHF4sc4IOpHKWCi2XB4mowYAUayAEDC03YHjBkMAgExiqP3EPgZ5nS
5pBDF/ILDshcBVnVE6DqrR9IMGjus3k+RCYdpEVyxULc2M4F7nhVdynRn2DLW/iw8ZG9RclXhQjl
rGXLEZT2FxjFoVidOPnLmUCwrwKPY7YgmmAcD8UUdU9tVv2xdqnCHISEHKXLaRRDmVfiZGPlbKxT
neIuuuvqswIm+8tA5OXiHJ7KQ+KxRHJOvIHWMyuZghQW1CuqK3fkabO8XAuiu+UXqyFnZ7VQ/5bf
IyapWwjdCSYbujvj2UA8GqsAT/XsvQpK2XAtyLmSRYBcr7ecyZDvXwi6d3SX4poAvGshwxWmFRTR
HWhRF4N+siv3whCETZhjljNnTBxsybm5bYla1ZUOGVnSDTGGHZWwBftlcsuymY6RywXtunfRGsWZ
D/IDxwvhuurnrta4+R4ykQCy6jxJuy4rhQDuzM8ZrBybeUJ/GkWXjyFwZEnrGu+smllivYTNmofi
zy2uu9uCkwCVgeEEN4XHVuJo27/QXs2RMM0gbgpHZm3afYzKyIft5H48He2Z2C/WSxjHQQBjvpVE
smqT8NJs50P2goNWERbQPvSrobbz1JBX2NhwEELefd884sRMM8S/Z3e/eBC6ldkQ98UcIljwzaKT
5vXvQ08WD15qpnzG8dXYxFM05fpFTQDkGWsENWx/EHWCA1DT16HyUzcoOhsXGijz/O2q/c8OgMXB
gsucNKI7+qzyghot2nRZZYqCzH/TSR/91K3EakfL7o5LKniQ+liFdaE89z6Mdat4Zk/jS9TQxI46
jivhTeuMLkWz4yZZXvHkfHd1nEtjt2WtkF3BVhUhwvJ6bv+33w8mk/90oWigPuZ4QKTrIzz+AoQt
cbFKy5IfHjSt9xZzES+xYEv/UQlLPZuhRYkc6yADvjBWC5isgXYhuJP9UPDCwxkOVFR7oKrLOfRQ
tkh79vOiyzgybvWNY1wCpkbSCZlDHvKxPdnVunIVSTSqk6+4Ucj9QIO02E1+UEq8Ft+wzvuM8MEF
TlpdZgr3nJWsGKJyUxOWHoOJh+rm+29yDTZ9XAUjIDL02W8Scq03QkYVATpGptcXeAI02TUNQ/To
qwlL8H/ZkFvCFmEyuHB/caIzfMj3Bzagn1F8pex5OSYyKNrdk3hALuMrLg6sRyGJqKfs6/dhoVhS
vJL4OqJ3bVuWj9PyrJDX6sptlPhlUsunm5EwPOeCruwtB4Ko4y+394KCet2LH479tkwTqagClxU5
BMTvSd4iZg38CDKmqd9CdqhQxSul3ZNEqM0jpExc8WPyJZ2TX9FNNTZNbGTpl5Hs4//WtZDk6QGr
/RoTB6ukC2046NAcJJZmfALqo+27p7d6BuOLeDNkDjNwCR5ft7ByaHFkHy0YRam64owF1Dl+tNuY
wDcTeJOgOgUTTDkXv/gjbgbuw/bkxRlwttrsJjspU2KZy6xCn6h07x3ClL1QBW08JK6BqzUtogbA
KfrC2JzSd2oOgSNW6bDsZm+mRI4+mg0zKqGxUaoo5uc2B/o8ldPiN236K3VAc9KcT0nKT3RPMhD9
b0WJ1qL462GwNb4jBYSg0gvLhyXvQyKhji/YG8+l0n0qolFC0NB52AzTrS1JI+UTZht+NjlVK51N
DvZZ2rFQAc77uCX74lJCf9BUoCaCVU+Dbb1LHefyJa3s09ItZUzo/ib5m4fwFJKsQAUmIiwf6HVc
JsrWBRhZeYubi9p3n4oAFZ06iu8jNnYczxOQbIsCt7ipMdBn1kK0seRrZDs5TaO396lWkelFtsNb
trvSPzY3SR5lGcJIF9wHXANp250jv8h4Dk80tA1k+OjCL4Jx/tfOMNrfH6SkV09Ekvij3a0HiIwz
tR8Htj5qoFTvpCVybbrvb5wQ1M2/Wx9bA4u0Ta07OUiqGGPAKAczVQh1e4nYdPPpZnmloLgy8oSk
Qy53hyeJ8kiqhP6PNrAJx7J6hsn6Cor2yDPmUQ/Oiib0yElDInsqEU7CtfSZdQxuQESvKqizwW8b
Z91wQQJBw13cR3Eebo3BdDBZFJEmhnGJxe+SYz/Z3MpuYXzy28rC3De2n2t00ZpVRED/fL0MURdz
J1NyOHkTGcSJ4jXv3l6f3GZdFPTQbyVZKRNgj7FVyX6lffrpS108oOVdJgeZw2GY7i4MehyO7xMv
dYmnqu15a8+VThG0rys90ljwYalODauwjJDStKVstv+F2Zpn6fXfFU6tqpvtKIJ3r1trOkvlqgRs
Htg9cUejn+YK+Jrjwmw6C8Ehg1ebFjiRj80+/weQF0R+ZEDd7aLyW+y/uOEZqapGK+PowpE44Ypr
KKBeks0up8+ysLtt3uC7NHvdK4dE3SjlVDPEt3JduQKjS0hsqhVzpgHERRIKdM3+G2LODawDDNTL
MivyXkQt5nKowsCHOe89vRccLe8qWabwbrrIxEeScQ6Tbco2G3tjx4yKLvtChBKAPsR9B9CiTNgp
wspEjBnzLfEcCMjFORklsd+7TOF/5mxIWgZ0CMqJivDMGEVjwIHubYnMYpLjlhv1gZz5cHHDKDDJ
eJCYGeaA0FK1k6tG4jmbB3ys99bT1THrZy2PqRjdcdQ12bhHt0De9Vq/xbH04cCT2NcI0ESK0xYZ
LOKJBCCjwP/mYqHF7zr3PILQlFeD6M8NWndmUTWc+/CIEhYnszkllyIQMPg7/hNmqwp+hA/RyoFO
2WM/n0oLE9oCbVTMMXwOwTrcvcMTFzDoDjdxaf2Q9mzjGtwlo9vqAKCLg7t9Bm2I2P8XYCiUCwjw
sN66y/LW6/fubMQzJ0QyJrJIN4f/4qH839mM90EhhB1oY7jxfzV5Ie/Ig6DNUEzdOFrYd2N/nflB
ALVfIBoSU+xInu1wovcSVi0t/ckQM6BKScuxPVqoizBIzVnPfU9AKfI1IXPmAi9TTrR4DXqz1gTz
6KWby2rgMuKpNcp8t7PH2agttxMpmSY2rdCmaNxuAOVm88mRiL9BH9SOPUNcp/SQwIpWkRDWNqRV
CX0HpJJqWfbOtvIsBnabQB3Qx1SyjbELo5p1yPvuB1OEvxkJwVME1R9vNumwQ7qHqBaRylYQMY7Q
boXmxW9od8ZqT4QikN0kq1ZDd1VmeznWX/oxqZpXqjS/TJVqsIZQKeWF7D+CckOGJi7sRAzjNEvw
D1PCtn/Vq7c7LSkqxuZIMlBiA44W/aQZquSSNl9GTrcmXpCeJmfLoGOfT1UaCaZrb73AAnA0ORLA
PpAGyb4KmVpoPm1NBXIeRw0Rc30m7uyrvfAgnqKLpNqqRsI/1O04bKUb0UsA9LWlYh8Qp7D5a1Jj
9FIVVJSeWgcs7DfsIUkoLgSaIRwCP1KlcGj1cNY1c8k2JOJXQYaAiGqL+CPOdJqXlSLwS7x78hG1
6bxhWgDe9miylwn8b4y0qEMHzm6hUzGrlpqu1dozvX9aIKHNSDWasRbqezjNoWnQ46xCjQZjNkv5
FdGHCIhP0XXM5dczTWbVyupnKinMfrLs/HRdgKCPGpEVfrGM0C9IU/LwkRyFsFnYH2GlG7lsLimG
kg6H0ZbEMVRaeQvzJVJho4h4yWdpWA7RsjSjmpfa8tbuileOx22aaV6GC7/dnVC/Ns5AMw7bF+Dh
qs9aBaypiKsG09/NgIX9t8NMuBcaVPOBTI3rLCTqVkambgJTy/v2Lk5g2SFnbP1nqydnJlm92+ri
07h4Dc4Kx5V26TCF3FeJsXxIf3Hg295QuYcajiJO6VLBg5aZgCFJBo/RLusu2J/5OsWbD8M8b6PH
e/eDzemUAg5sprLYVkhJl12uYwGtVQyVvxiIN//fS96B02pKaFpcZ9xsx9jT8QBB1u6wEzv/s6sH
9jN95NYs+htqDDj5yuYqH/4vBdgYIlo0YWMUY6+U+lC1oCro5RdhvOhRwgLmdv3aMKSxNjjODirV
njE03Rz4qwiPu77Hhwc8KXE7LW3Q2WPtLmz3YJ8NRQgDsrgpyeMimjeLckstkhKDEhQk5fr5eIX1
eFqJgPwd/Qt43StNV5hTSOMoSVrLW2exUT2HustSMOtMJauHZLoaDPHtFoModwH+bn0PL+++6BoI
vyZssp/Tj9I2B9i+B++gn/35pQGlc6G2kN1gvfyzglR56ABMtCPBQAq7vZZbOLLCISjzf8qfn3CY
RQajB5SbwGhip+kDLDmQ80gf9lX8r3LYNos8YpSJcBls63iS8TwPBctT+x7A6hdZyfnMIOO1EoCR
gSA63001xY3qTRn/DbuyEzquBFTcNmCkSTcb2VR2tvn+AkkV+HL9TcjsBzKv77MmFeP3vcECCVnc
R2pzubfe1R/1rdVmTcBfkCgeyBWhTD6sL4ZWGPkZYDHu+x8R6PC/STVAMz+7nz/qcDxZlmMTwM2R
FdsGgk5xL6bZB9B3jrkHTHGnkNW5bq7zCbY9dwHoRllGtjj+8HKp546jYYVyFvGTB2W/02ClobX9
yfWHpHQIgn+sq3kWtxhSKjHA7z8mk2VaurvyJVZvRFpjO/q820eEz2+ML8oa9KvGeYCKrOwS2ctS
3pPUZsVteSjTY5D5OrYN7Hc4mrvzDX4CHPxbhs1vyG118uwT0XGkp0ZW6ztqNxd/IV5TpZMFXjCc
AgmPte9SXX95VRNvu8FtoogCpeu8SHgHajJuPXRcU5ypTP171vOhZbphsWF7oR/KfxBDh4qXPf17
avkdwC5LKeMYcXAUq6mm94Z5Bc3GCxdz4zAcM8OGxOocViplB+E/iaJza/qvypqRxWKH/X2f9dfg
7Y1NL7S6llE9WvH8V5ogqwCsLR2bWtidbWOL1YeGxIsYz46K0vc1lXALTEtE52j3MZ36t7AMAyhv
shlSDSkT9Ifvimfu7d/HnHVu+iWbr9/p1doTkNkqNyn9zYptj3A7FeygLRa6/wsi3XiIiHyVXorN
T/3ib4ovJ+sBL0Y+L8pesi3tXZT4bLKbpZpjGMdIwWR+AC6Szek+RUGuqouFoC5Bx4tekChWEbK5
Gz7RTCI5typM31BX7SJdDIMZDrFpN3b1TWWnITyq76OhpHeg7KoeDiKXVexpGOMU7LczAgEFWGzu
W4AtNAnOlf++aXJ9wR4Jpn8REIX24mBMZzHnVhNyXcJN8RHf1txE8rATlif7HDb05zz6cGQoTC3N
ck+lRRKETVYLW/qx9Cw0UDP3IyGkbOm1lbmw0+KGiF3ogKSEId2b3LDYE492YO4j6Yu0ZQRsmAMS
GYOGo5eNayBiqM190N1qEw3LpKTEt/gxPG48+WoGCA/w41hD1sYYvW+IFFGmdU53+rFuDbPPUV47
iX0uV7ufKDEzSfKSVP5oPfOfmjuUlpOgr31Xq6/oga1ufHbwztuVMhYgDzyNNSn8nh1VFFMEU2X/
D3KsomDejAOvHj8bDcOeaBpeo6yGhEZUVPl24EafTY3ww382RLuy3jxajVN3ckZ/0A+eXWxAZ4K2
GL3/mSFQCDswvSsJlwMeNTRIgvXoL8pvcVVw2vJpUdf3CcjiJ/mJtSANWGdJkoXKzLcM+waaA/mU
yBRaBDMpuI4r9ruRZ8qNUh4g8p7KG1/9AbkcbWFFhf02C84KZwPimvRCq9+hPrhEnmvaxuqNhdKK
doAo4ryIp1chtzGQxs21rfOWNfrQuLuFwXlT0HiHmLReMyeb4WqgJ+tawY8pJXP33Mysc4VPoDEi
khgmA97KaYrfemf9rq8AUOagnh+5oFWUmaG/xON0NhiA8Ge7bilLZOUGGlk5hJdWE/paeHA1ZFht
fDahmy/pOIdM7qwerPdnqf5icfg3Sq3byXw12hqi34XQASy546Zci/t0fagD9GIM7sRLjnFXSXwa
DdNLrVP3hTAiGmEFpii2sKfRf+plE4EptZ0qda4Vp08xfsMKwhr1Ob1uc0vT1HsXuGWYMHtN0ZuQ
3+ybSMuOSpormY3l7pXrN28z6+e+4tPjx5Py22gh9PwdGHjQ6C82RIrpp7OIie+Qnl2OCGjehrFs
Llr1hY/KOxEZY5qzqrMbgo4ThzqeArMy3FPi58zR2L4nejtak/bcPc5oZudh1PN6m7SznUURXPls
fBG/Gi/VybvVF5i27wRVi+SXD4n610/+UIU+1O+hQSy6Gy5743YGCP+DXeGtPVOmcBcGesRMj+vr
/3qtJoyVZybeNpZb8Aho7g4YtcW3Mip8rb/43Fc20jzKhquaOITbl2bCClYFV15x6xiu5vTQ0Lcu
8FqoTeGvdWGuq/ZyKvGNV+u3+7HywYpTEJZcFAcBBBP429mWxynhlVoR68Ctnk38TVhaVMV5uuO4
TvDNTBiGjYJw00sJyLc0F1jGZ+wxY1eo15924Q+dp/3PseKLvsZWfX6PPSeV8xOmQdMhKRnY648T
Dct6n3FhFm3Xw8DEELyxYY9CxKzvkMH7yv7eiDqtk/Mt+dQ1UeYDU13+FN2evdy9Ee7OFAYwXpLh
vWn2EgNEz5LGBu6HQ9SlzwZsECz/4SV3YaX34feo6GYNe+XuMYZwWbvAvhCe61fzglyvPLekszOt
Sbhpqx7HcrFZFwybtZ39WZhCnf1g9BYNNqIo6CEBoQMuTiAnncLtC9wFjyYo5VzFtDrvvi5go8df
sC/wQUXOy22TxFmseq8mxaW0jdk/UClkwc3RZlBDoEXSa9veVo35s1eOOE4g3+SERrfA2ghvbaqo
qX+Z/Z886ZBCfZsZNSVmBrQleV+XnPeCPlGB5XG+Y/KjgONBnKL8zHxEvUZvnf3H7Lc6IWkwuUBO
ODbpyk5RLdYuu4axozKp1dhC43kuYT6aXMI91lVkt/M787xkJIousr5X1yF85lnMI95fSFaV3cDo
C/YV3Nq0AgeRbPZerCG/nVJChCn1XR9qyvcIfbXju+RJnV2FgrCvgAHcawAkwl6CniWcCSPazjvA
I1Wpsn6NSqIAmLAFdX/Qt80La1D1Ftupp1qLFgm/RlL669BXJLvsF64W6f5XW+XrAYvqRxn+w007
Bu/2oWG6DDn7EKjyd3ZW4iBRU5bCE6KcZE2jwjg2PJaLpqz80L+5DoHgGq+PgRBE7Blv93C/fmFd
Xwj2cfBsJzoSp0qh6Sftf1+K5V8VklqJrrPLghalub2HS/LpHe/Fay9gMd5lfOlrVMaUhTGnDokf
heHSajNM9wttPKoSV8ls+aKX0m/6/Mmyqdl10qbwtr557aKPYgn8oO/moh97OHrsulIV1d59qe0k
bKsCAyWuwUzSMmm+8tjvso4pAcMU85RWP9LMOiKgR5wPTuCqdnuytKTW2StRwQP0gano8W8lyiC4
ymUl1566EyETHy/y9nIh9sGFxIHodqcHrKTtrFqkdtrLRlxtkg697RoT/NGLqqEbf3YB0FjTJf3X
XOErA2dC+kAw5XEoCaqcOMQfUKPX1QpK/pp6WDjrkOfZ4LIeghJhHUlKuoWcmC466q2A5TjzwVSN
GSg0P24ioVZ1QEDxSfsj2FUXm4Pw50KRvg+AXWBDh1xyshg57Yh2NEePorNeooWyDlrqvf6h5sWG
K/YWxzS7lbG8CK3yGNs5b0Vd3/0Fhbwbhda1dbDPzT3kUGgt27V7ux6llkSUew+fSxigGtu0A0qr
Qbr+ni7hS/ma9aCvULfuoy02Xna6iQHbACoZFyDpehDz2BP0kuLWf20qsDNesehq2jx4Swp0r5T8
rioliJO/D+4ndWeqRHfjDpzGZOXCyCAoPclUmFSjRh/B2vkD4Jizl94ncF/YwHFod96qvNgI8XHz
Sa5Aybaiy7LD2xy7zmIT5BGFsxDTFhoM2M1QShKyOos3UKGXHgOzX/2Z39ia/tnObbw8EK3XjBMF
9DDrPKUHzNgyD/UWTGCiy5GqJ9jO19b+mrU0dDjgdzirlX2HmGPCZdUaWGfGHN0sgbNDWxSHL7AJ
ACRWsi44yIiuSfV93KtK89gBbiNwQ7Do/bnezaHJofyZ0bWKt9tNQfXZXk8yV13EwCgn+BEP28Oe
okYx43g31vPMyEevgkgxR226A++3a9zdr4/BmIq7GNcR+dfv3lJj6fZjKGRi3jyKEgfQ0lWAkg3Z
Syx2OGnX4lJlZrIgZwut3TsjZGOYf609bCZAZHY79yjM47vFURGmwSFfmRkRowklgHoxUhOp87NI
5Fs5wBOBRdZgWMiL6eYpVpUT7j83JVGrYnvtxX7Lvswz87C15OGHNAfMc9Rn1t5ojyhoBUwa7Lrs
k98xW8J0DvXBZ8Sw0InKNBzesVYWJGOIwju7Lo8lI3aXLpxsxpYC/QHvn0T7D+SDtJq1SKR1mGL9
IEa/X2gG8dxrUwnBGTac3IezpOZaVHLwRMy5ps+m7lEBldx8PiaAnZKvWdiHj/TskhMsuPBIqbbE
84FX9G1OZHYfdBtkXw2NaGdPmkPxBUUYu2a/ZSrZM7fv23L8Xpeusr5SVDe8edwuZRj+v9TYAhpO
8Ur8j3LZVur5bwEBz8qTGt1fmYPwf/lYdJ/QsI/OKlFlAeFayno/xpu9M0rDGWBpbio6wmEPm32E
1wVRDDDVE+3Dqf0LVkAJwDPEp224EUw5/l9ozDkNAEa8okSQPOhBCuEb1NPDS2qIDjK9DF0V31K7
qEk6OkxLTpkbzvUESufPG+FOrVKXzBkxaiDkJM67TLP834hAjVig6pp7xH3Rzk6K6FUC+LlQjM5K
u9Zbwz9YOlRQfqO3s9ydo4Oc0ptnn5RqYV4L00qULtF6WZfbDY8SCl7RTVXSM2gM7XsWra8mynM7
jzar2LWObJGtOrJzL/kut7jkBEg9kqE8ePsyvsbsTuWlA5xaFrPzi8tvWvQ4NTlZmXTE+pN1MDg3
s875GQznIeIUDVLZTq+jbd6hjdiE6nsGuLPBx5fjZZv1juXh5WziEXHOzJiVUDKFMExfAfpOWl+u
O6/H4FS8fgb7aIY3vWL4rYG/9ItYZAttHtn5s3tJpLeciXd5NkGS3kpMJ0JOiV90XMRCtksxOOqF
t8+/AJdAT5gax771CNHuRsJqXsU4OgadZ13G5U57CDJanNWFoqbvYUvEAxYyey2SBiYBsFqUJnOK
4tHdG/jjSfEsstlvtjjzx7GEqdYLR3yChwVTyhFG1DNSe87I2a7llThxwnBpwOG42656L6Jb+etp
3QtBZgjGSv+4Q6nmgrxtHUcp/3ZxwTRnKxey8d/NjyGw4hiPfL+AiDKquway4nwSF8DeEeWlNvOO
xiYBgMoTLqRhDWYTpRvz0wuL2CYZpgtjlkC8ka4W0AUMzi25YbvejsjuUp2mlBAQ/DgiEnZt4b0D
QrAn5h1qRnhTlldG9IHcBZB0P7QCYfnwhzUGchYxtYayQJU+ZAvmY07tGjX/kmE0/ZSLpF5zfpP0
BLPVSwROnv/9uH7xQokuDAo9S7/22lyTH4tkPWlUMTf+UfeqfdG31kaqrFORIwyaLbjamymgPhXY
4hyIGGprZdv+BntdIq4j2y9wnC5jST4HHDbvLeXOO68614s89FtHkVHYIzWG8B7LobKJaJADCAdS
gleDiUjtmrvocJdxTYAymfK5NQ+iqJiku4JWG12rwlWBqiXiEE8WhUfHkSLNCDMUmgDIhR6ONets
Mz+b2IdPdehDutZ1RrCa9Uv4mZU2z0Sz7IMljQICEmyD1m7wOwIulqziwLTs5e1bqqL0XKmzCugD
LFvwSPXxodcv9tUIvMVH90cp7RuJGND6SWz8dxGDB5ODV2udYqlbgkRh3PZeaDXsVaTRvnWPBvsk
m5gT6Lcijk209x+YMNufUEbU5xAFVSOhnZfByBennjX0E3xKYchUIeEUD3hKTqA91Q5y/clY1eX+
TvZ+dPYZQMoGnVA54qG7qhoa1pBQV7Gm5FDgmcD1M+/0IV9ejUEyZaAgRiJ7Fe6Vb5iPZNxuf6Y1
rJrZLec1NwilIKPPtUKnUB+fBLHEXQt2sOqmTaj/GO8xjAFsNuTckmp8ZS6FzWIkyym7YTOBp1Z/
BP5PUk9j/1IA0pQYvHbVjRgLhKCXWeYvdWuO5Wx7eo6w4AUI+M8XC4Agnucz2pPFuOW9yXlwv6TE
bBDWMWd+wgWK+tpA93Yge92E2ZsQqrInsjkNAny5thLf9NxCJFUwRMGJ+VUtLT9f8j3tzk9VwWEt
WkTyjGOXT4d495NFP4xBSxkb3iTBYN1j7aBZ4lEHbE71BdxX9ITkBjIln2VLQbNy7Iq7gJzGn/Dw
Giuoc7m8irAEsSTKKDBWdUa3hw0ON4UTHC5WFme0iIkAzy1pmu1YIjPI4wQRpKTB4Y4QaVToyLH3
NyF3U/d9xBp7s4VRFAfxagF/b2Us8hbTMOQqXysNULnxFwk/XbO4j7OraCTErFTZmwpF/d9mUoQc
p5SCAh/utHr6F5eOltCciReHcPTfvVxdoCw+5TwDbVriVV3BEE5ujcxcQICr5VFmB7fwOOyumXCn
rF0QimNMY8Ki5nd9qgA4uyB11ajIOCORSIxCii0sY3aKqxE5m2UsxQF+yufXyDY3n5vyw3QbPmgH
eMty4GPT4meosQ5vakNOUr7YXTKqRBCEzP6Cc7HT009p6hYHwikyp05WDPvRCNMb7CgFtCvYavEW
M3q7icPesheeJ8w2rnWwAIRraB93bLgwZA0/9wly9etQDeSE+fSDbr8miIVpRbwoTI8z8E9jtzGw
HZrpPjwhtNGMVBUJ4+U0oO8LVSmBKMU9ijI0gWoyG7EdX1O/QrSXLXs1wJ75ASsFeSYqD9d4N1n1
vMKm5c9cWjpT7gs/3dK9FVyKHflzVzSQ4DyLvPxe3SLwq1uwwxTJZE471IxFePLWwWWAS3GI6Fiy
X0B2mcqrRs067l/XdWeGoy4TYXws25XJMYwHJ/1opIvYSQmTlMNobtp/zRHYK00bGOi0xmMpMOa+
DMBxNyByEFsfMyLaH/wZjrPPW0fXAuX9I0PV4tye10IGaOD3QNh3p792+amsUC71gjip2xEAb55U
RjKXXvwTzIFeUTwsjmq+EWVhnx2R95xlivEMg5+3ZxcjZKMj5EyDJA9t33tJ9tROJNd2g6oKH5de
F67P6CL/b6iqaCopFXrZnzhXed7VeszLbnWWSoeKdSwnypZd7yrMiP47L+/d3yaL7ZWfLPNq59Vz
DdOfL9osEQZ03lZXoDaB4vLzGJ/nQgen6XslCM3jk+dxxTT/2H1K5/PiUG+YgfB2p3BhT6E+oyvO
6TvyOlsC4RsAxUb1tym0rhViX/Kjbz+d4rZ+aLCT0Qfl+e0nHv9lsedCq36zdSWMnRrObqF1k94A
oPVOElkZLQENf1XmTd7JQKR/kfGPg4j2vhNPvsnKfxIoA2N9KBXN2MhXWoj/Q3Zt7mQyCV8qq0wg
q1s/K/BVwAshQZws6YegOYXr4AWWesD+yoqx/FDXGUWRCyb77u1fkl+oIWuct15T3ls/25EKD/p2
eUkrGEXzr/di6IBXrIHlhnkXMGOTV1uoFEo6w0C94shIwPgHEM0FKFidJH6uot64mi6f2Z/Z7Ead
fu9COIUVUpzRfyB6eeS67M+46SGqfJhxF0+1Pt0kQSaEpbR9tVn5t5vG3JeWFqG7pT5d5w52ZZ24
vZE0DY5yCKZiYH1qnLTxq8gZQIClui8YShwMnKu3AxCov+9NbxesngpZV9pUqIuItYf+Lyx90cur
ObuGT4dcht6scmRNYzLvHOQ1zLfM/QFyyqrzSGgmmQCtsU5wEEa4hQReMlpQtKq1RKXUlPL09CjT
cHrBcqeYhqCUvVikWsxCKzh9Zjt9XOg6f75IHScp1kjm2+rQY5pipsgRg8KJ6tWoSDk8kHbInCgD
JcC7+eS6MWetZxy2NEP2Za1GwTazOLIRT3exR6KttP+ZMT+H+/VYK0DnXB3Dx3Bsqa/bmaGaviVN
kHx4qKGiGQLskzWbysoWw8q62OItBASweNCn2FnhaYCcKwNFbw4A+ulzJfO3WC4QxmBuDeAtQx99
G1ch7bwa9ZtVHQToOjzHXJvWI3YiDfscByHti0PBWpYjWoQyvNxyf6f0SZYrFfmbxVFM7tYtTliL
uqM0lOVUh9NFvhZgZEZK2X0wKqNhzr6dXSx97dWMZOu9tfQMUoyi5PyyFimd1HaZB8Kb+kLmScYI
v6rqnBPn37uOZeL6F5I5G6Whh8Zn99dA5Aq73Yby1GvhuprGXCkzALB51ntXqPB2YLnWT2FhdE3/
bGz7cmwDEwIbXUTd0dt7EIOCmMu8DJad2zCC776uoSrlkPFBdbbuY3ywJlTcU97i41fgIR0MnK0r
XYvX5yOMGERCtVi3+mWauzHrRwuVlOLunST4x4sHKcz2EB+hQcVkGbp84W4LqkhCXHsLUfvTFFv+
SRZ/JR6eHQAdSo4LmwmdJ/w9oHeaYiCnP4StihW+Bun3JvVmFFSNlrCHl4V1wZVtlHU5Yptn/3uh
CRf0wREI38Cx0ODnQZIfl9keFEYsKWn8s7EpeiNouIBa0KHbkFT+PG3LW/KwOZ+oUIGANMQ7BWep
+nKiS/BLHUaJmKlIvnDwStRNiY87TPckA4C39QnfrRu06b5Z8oT/CyIm7IikG0RPuBcMzC0xAohC
jiCfX3J18v7LBC2eo3O58tTSnb3KK1BJVZNz/3L9y36HsZwTUsDmknuHomCD9YD3DF6yqyDBDwLf
vz8DKScPY0YN8/vTi+OvnYcbwMDWpw135SE+W0D3sNbKIIZFPXiTAZru6OA1lC8ZWzIbF4UbTeY5
ndUU9qc9Cy/zGosOPqiBHVN8tT6VbsIj/znHX32Fcrxmh02F3cx1zwds9eJp6/DCwIlV1O7lLXz6
HSeR0C4ChZXMaLQeCTtXpw/5Czabmra2pTMf5w3hI95sGdsqURXfpkYFrz1lFRnDbPZIM7p9NSdY
Np9FCLhd1tcvwyBY/iv72J7KZCaQPsJsxSKmWQ68Mq30Xt4TTNw7XvoV40jHJijnj7rOBznBX3X2
uinzs9uFEXc3kOJ5P2o/SrZ1jJsEI7rtMYdR1osZycnGCDEkAS8pAqUXbdO7Rywh2mV0wYm8/hNp
yPXh9/sUAg8zrLeYYZWEOLz32gd/I6+O39zi2PUNBdSFJ3Yc9iY/SHDcIJ7IDoIW7sVHVvGt2tFd
tIFxXrMzG1ssJitzWKUzGKC3AGuiNGgDBWr05pBs21uBgQ1J8h4aBxmjuXiZUNmfuaXQ1OfRG/Qx
PXU96EV6cBsn1o0WCKy1686qf0gri/mVKa3/dgPcUJYMwtW4CpApTvBPFGDM4cDY1CCTP/UALqLr
vN3sPfQpj0026HQG1+jfmsCW6p2rsMF/BF6Z5LP+o6ewUJ6XnLxGwpvekczZqm03p0HXcz/4f60m
r1FNYuCwDM+R7T8uIjhnSz1SSqm38KjxiY+QOnI8zw4X2xc2Zked+ISP2G+Qds3giqy4X6xVJfLU
aR/aqm+NX/QmkDiF/lSshcjZ/sJVste8Il7WrVHekIE+4g8OZLq4BPwvaUdF1BLdEuLmPcI0QmEa
Tg3Ns6Yowm7MofNSRJmwgQKVNXRo7o0m0LJHghywj6iTX1cLOMnO7hgwsX/Ii5FtUqME7IMeiOv6
lr9ulIQarbAsc7z1E5HEH31FexSnhi3quq/z76dHKKm+jNez4IFTwo0Bx7OOJefrFT9vsEDJQ61L
ccp7XDhRkOh8VQzEHr6VhFF8Od0egJsCFW7Yu5aGxW4nznnNw2Na6dRyX2L8nKabk9n3hiB/G6ac
XHq3+F3Mpqcri9qmHqBCglqwrQIwOwB8uZ2mueZvrw/q6CnnIDNnVu7ZxiB0v/s+4t83LeXIKf4t
xyTSmQiOrxIzlq2eo7gV1ITQ1K441xZ9+JaAtGL0yWyl5BeKQ/IQWiHEdHmzGE69euRnxtv7TJd6
ws1TI9LGeod6P6hZQovx+the0iuZnISsVFCH/d+kgaDWa8EWKCObZjucLCda6kuGX3Bm0w2zaMHR
e170pAA/p97fWjntKvAzhJD+QYBdyXTd0AYy0l/MyOAtBkW/mJXiN2yAS4dNwoS53jBkGv2JYroX
8OKmTPCoCody1gDf+OpO9Z1izH+eAco2AY+s8O1uPAvFkyAyHFADyZiif02QTyKmSCCXbLV3rfZP
22Aiu3tsZBvT0NtBc1pD1wt9h6rPGAW3w44FWRPhFasYtkdstnXDKCR/zLF6DB/64HTK86o0ZdwK
jnbKy9uRyzTEtPsPA72o3m5s/P98zG7Tu8ALQ2W2NQblQs5/A7FhDmeN92qxIO6+Y8HO48bnN/OL
60LwrzRyyb1JYS87CX7bIB7FBWNnp2/TnXSti5zlzbjySRb0XV6gG64rUbx6YpAWLO+lLY8goVAv
/oqwaA/w37ArUducXVgvew+z3mVhX5Rd0aPU7mkCNFtIz3iJeCneiWgPpuHYFH8nsYlp5Ffj7dD4
XHDpNQMI7DNYyF7Z8Xy+DOL1h6hxXIi2TkCUcN7geOZgwxvgKiUeYu7v8g8HgMIeOxuBdoIFKFjM
7YkmfSBVrTy2Ww9AC4/Dh4GFxxHhCK+CNIs4KjAAaKjWfoE2QtyR0VEIOcc04ryWAlfeFj0DpoSR
APYDE9sJJYsuCLinpJkjeU4p74FKCviwD327vz0X73kBR1pQxKkfOsouqj1FHXyL63TrNInM4wb5
PVUzBwYBXAX9CYFyz9TLrY3vRK/JPnmawGwFsu5kMQDcIsdcAXKVxfN3x9G/Fzlj9BPbOv3fcBha
ON0qIibbJH+qotpL+WRP+tL6d8Pg46SKjC/lfNo54pUpsP6ZTQa7udMByvLEIyIbMGXx1blLmLTd
NQM72J8JDfm5BxrcH56sOJHN7rtzwuWrJFdeiklG2qwmmfbfbX5psBRHELDCoMiwcBUg5lHBzo9F
MOWc0N4+ag6hVYuj8Y7O32pzUZNerxC4p25nuTGH3X3vumYk6zMDOhuj/rq64tA/Kobf6az8zXWU
yktN7fynF/9R1Bl5wgz9Afy6OG5dMgahsfaY0v9wx3kkwFD1aHfRhsaBRY3aYru2J1AO+dLpdiA8
P1HtUz4aKtzqm5/1HmbOb3Xc6bgLAx2BDdjqUhpQfcHqzag7hVmXRTJbp9aI6UDP4YJtwIkDLlny
0Yp1vctMZWk48cH1LeUJr2UMm/FmgNYnf98kjLSjqiAcN/BhgiC47CANcLvKlgctE9Hl+Lai+m5c
i3L4u5+R708lCSebUmjNCaX7vi+LUE6Lodcd7WI6ZUmQl+Qubw3FAwOASyKdz7T8nSJG0OgrVZ6K
YkhNcaGlPggk6b2isgf6Izoyxjs6SM8BpqSNiwXKFx42a0K0CZW2MziW3gP/6/LXw6mSeEilhSSD
eyBedAvef8HDlNRtsMGclJjpAQPcWo6+5nZqQsr/2qS7+Gn5aStL2JoonOstGSK6IFaypiYisolH
wutokjpVHMvKX9J6RQCs72pqQDhyqIjw5oZW0XGduGIiN0LYynbn526+ol00HbRMfTh5Z1XOXwmq
tZKNZpHpTFQQYByOC+i/4prkz4DmyacwiDE4EYH6BUzWG2p4GUJXk1rwIOOG1SEBMlRaD+XeIgH1
OEW4cdzyJJdnHaFevpNbZM/62RHFxyFY+wE6cl5Cpu9BiaILlC3DpsrJpCoXIdjMT3zzcqqLxSE3
liHJt31TYLvOn5K2tuoyScnuJhzGhAWvy5tpCKwrcy2SLvkHJ5c8cM/wpuNo4R6vyun2n7U3Awlh
EIfqKgBe6cPF/JKBPgBTn0xoyyZe1sCQFLvC+weo0GwBG0ba0CgCwHTEsC7H7uREO28Vqr0Ja7CD
zTHQGMMnx5u4xa+Tjrmw8OR71TfXGPD9Cmr5d3y58p/MFtLtrfJ3BUTZL9At0zX5ftNhYHyQse1Q
Ho6E7qmtAE2j3na82rZzD/q8I4k64VCJjDCBu8QI3mY6No2BD48u8ayJZrEU3SOC+ob4/nObhmcR
KttEnNjfnUYVdIIGBxL1Ia9+JEXamdro3oIoG2yfEPoeC82HZkgEMoO6y8BGRGMC3yy5GAb6o603
zp4g0oI3xi2+W4P0+9lH/GyjXdAjoxtXbSIfQlbp4Q2Ur1pkK1v7tEyuXIUmZM3E+sInvlIy/dwK
J/lp80z+EYCkrX/fj8ZDz6/SfHAzefPVQSXq7B1H0s3rirwRyEQSuenQMXadreX79Oo2WlUSynv5
v2mnsTNmBYDjYQ8VWEuBLneWOa5f0EwtinGPmn1WqtBFwaHiZv3oOJilShA3ZY4yzw0XtE6l1q/Q
Hf9/foHOlrCzZ14YHOH00iN9CeNEczAzjqpiEOXRGJL5vyBjf08ShM4Ds4Wen20WCeizlW9kKrM9
WhGAtHO3gc2fN1nhlRJczLtVOFklk5hwY437E/kcISA8cyrThzhD/dJ4wJDAWkMRetzdieSQWBwn
S04aqHc1tRVAGFJiagd2werjYJjbk0KjFyw1nb0O3KQ7ZcOnf1gt0Nz6+byLjMIkVnBGG1sTGH7l
w1OEly1Pjjau7MvvHSW2hvtsaQ4OSaXRbuzf68zcubUu1ozH98ddyhdNXa0CHFDgocD+1Yo9Ia8W
NODoa2fsaZSQoOqd32ZNvx55cKZ8w1lnSR7FldXtfgMrlNJKVTPOMSos466qWUS43Em9B87qPbAr
BeJuT7zj/CQOQNcmY98EqjubzG+xcIURLuGwAgUjk0YSox6+jNUlbR2fc3vYyUwkUyjKKUICbzE5
R6jdd9BOHPHF7ocoACmhY0J6VEq/nAgC0P57OJIbIPQW/2Et+SCa0GP5qf/bvnUPz0/m/Wa/U4ah
qxLI/43540TvwnIUYBmh/D27iNQJDCcTQDQZz15I+yJoFU/YmpPdCE5J9gfHBAd85r/lGvaKcTh4
dsktdXp2G9LULJEXItoa5HSwP6+0HdhXDGm64PNqUbk6SZlauQbHvTXeqD/+pSaMR6eq8IdpIK6p
dOjl4NepOAOg2k0EZJuKhCCJb2kHTHXNTdUB8RQWDAhPadnTKRT4s3t66HVd1XSGAvnN3ZanumyK
4MCagDAEF6fyrTDdK5Tubl66ypFjy9LaCfLlfXwiLJP5JaADvvU4cKDNL0K1/NbJYiPmfBEYQxSC
L9otMJCfgjy54hyn/bxnEqXKSk+mRyPJlN8CSi4JzJVvwsW7OQKfWm1aCjlSNAPYyq0vWi0Jv7Bh
yueTyfirLO2TsYI+4hfOZIKpidxlBa2aXr3BJpFarrNR7lkBE9giAKmr3jnXxxBpzuRf19Jsog7b
Tuv40Y1Lb6kcCumqJTR25+MPoMV8mmHRI3vWE1L5SEwgEG7AhOaZGUGvfZ7NKlYZURaj5R7rw/Zl
Ggl/MLjLcuHX5cNgHtZGOLkzUC9UgcHtuIJFmFCymRD2Iyzgms/yUTraISN9i6eBJe/jhE82Nefx
2Ll5SpYAr2izzA8z1cQkiSMIehI8yYR0JwAn4ZRqeJMI1jNCHx01ALVD21DlCg2spA0tn4lJ7Kla
YRssSJnyUTJkJ0eJ2VpKoNqLnRaHApUPCr1PSC/ApAPCqoTUGVMC6W6QirPo2KZo9kCiE04TuUJS
7puq7jCMGnHn/otjcMc3ebfklIQ1fMLuKw3dXx4BiaMWhzCatbewYsbzciqHJgj5jQjlSt7Wzzvy
X5gBIyZqdcZcR3PwfN1eW5Ms5aPrf9QimenIMT8IWo6531tJ30qnoX8xFCGlIvZ8cJQz/a351Udq
mekJuNkEmY21OYrvDMNYHaLwcgKTS/plwrJwQqJo6wOaAXSCqNawe5gxQsY1kK0lbhXcWp7C65Th
6RSt/JeQWQkcQL0F3frXN10KgQV7rxvd8a8px4vrel2oYTWOssM3A/BAZcIMd5NRqpwok10uM1yK
Yk6Q3pcVKSVQ8E4WMYdQU7p5ipTLjg8KeQwRyUT5dp5p0zt5bFNxgyWxMhgD0YwAjfRAoFvLTCA/
PBB9dHaytNSQw14S3M3KFkgekrULY/RgkKQr3HFoB7DYYecoUhsiJ444rGLn86zbMPQzFnpDEuN8
XqJTWHviQdE3Y1Q0xnvyqx6UeB8KQLVkDeqs/UuXk7k1bSu4Ix/KPJGpGWMRQ1Qis+JsGw9kJbez
gYMlwiiT3N8cCfJzLxKv5ZmzvmK1FhL8PZr4krbK07faQy32e0cx8q9Qa2idj5w9kiyfw+2uni14
BEtVns+OZdJhV7xldCtQ7azBSM/box3BmSJiXikij9xzHmBr1EpvHxgEM02fYmIkWkgr6JlSIxbR
voAyJ/JvIipTxcbLvZf8/m5fvkB+FYISmwfvCT6J82zUJdoH6GWxuJAM+KQRNi20NQ9Ss9MQ33uc
dqNX4LEVHQpKJhcmrsmLkMirrJVV7eY1mRQGr+AsO7xOfHDzCEfmcXJJIRnDm9bIkBjOTLqeuQQV
ueiNi+IUlcaFN06Ef5CQrMm73AEb+6N311PpgJNCZkec0OoXTDEDapGHbeBpCAUcCnsMjYwgdK0/
iAkTsgCv8ziA7aTEbXH8BuCNTXfEMsLTqEdQ38loOGqN7J+qjWStiAyHWVm5MYVXFZ9vzLSGNw7b
95nGRvuQpOEp6TtrnaWtDKjpN8LioIR9ysAC+7XoQQJaGA4eHu5V2TWruIrMsg8oRexIHg6DdaRp
WrZYFTGEdNS4V5axvNFKxMsal+BRjNEsf2R3o0sak4uhcXdSla6CRoCNSAktQYAakFqDUYDKfA9I
ibqDoWNOVX1bxGLCEWl8tXOC+JgiqGd2cQ4Syc7rLzxsykVNTZwa9qyyejSIYNi7HXIdFIHQsXvR
KOsZOZZYa6wqE/EMdj9GM0UmRM1YZMekPG+VDK0QEZSgNCM6twjeLS3imCUM/Gt2jZ+72bStV7fT
yNvIfD9tZzbqVWtOhQG5sQSUp4aO3RBZOiIgtgkKKUhEA7tgYd86nQbFRyYUffXAXs5nmalSFixC
4uCHgIMVjwFm/LMe8WKbG2LAPRKzNJ+zU2mRDKXijErutNhQgG55cg/YyupkmbJ8PsH0JZLMmfWJ
7FPgFNktPaxnE0V4ZVndLhYN11nxBp7iJS2BxlphPdP8MPGaR/W/B9Tjz0M24wSF1IQ3b5ASTNhL
aPRYp3aHb4jjdV6D1NTs3GkuFUxtmFV1tajkx7bvA1KmZ4k6QxDp3GAAd3MduQ1fJuS6T1UBxKy2
YFu6e3EiE1c7J7qAPn0qBDyu0H6goE3E9dlIdIse1P8T0XooSWyJ+WHHkQSrAWdzBsQKFtaV0fM0
AXxhW/xAtnGZI/W5TANeItS6Cc6VVdpWvDZWgjRBVkcfT0tcioz1GnR27CZzJ3OLYkTqfqtQvVlp
XCYMTUXovxpqCzTg51TltrwyCiKZ4VTGeTA1BYogOmoGAe7iYJSnpM+4O/GIOiBGTNK4y3PhLBt3
vx9KztIA/62NZl3Yln9V+yAoMOKvrxoUFxEMT11RbCqUXOhjT7Pcbadxvz7u/rhVr9x/R9ThIq5F
eb7Eu9m8EiWxxHJwUvt4+7pHAEP+lwFSC7ObYWJK/czBi3iezxcBxduO+T6A5ah8YBuajBDDKIOm
u82yGu/IWe6D1/y2n3urduX4XjKd/jaZZiFtRhjBihxWKAgB4LNIUFDjkr0RzJFQjRwjYRnMrF3h
K6l+wMQk4y/m2wQGYyZbbkCL6UGfVm1WjCSIyEB6KtF3E5Pe1idjDyWcVSx8e+v8c6g4+r1BHqFE
9LvQ2rCtxtuOhpm+xARIBsX/zWWmJZ9IjMI07rgxeVTQfpUQGVHBJRV0jh0h8FqrP9qavbhry5XP
5ZXLAg4l/Aev8LVkCAHgVUoJjVSvNTROoo9oBcPRkuxvKzRHZQGBHeet9HSZeM5TKozTznHkzaiW
laOt6lUKhEPg8c52aXbgm92yhb81Iup95VgklzHfoI040owgO6O0ZU+9Vo8gb1PRe9v7yd+pkyZP
Kmwugd85xa2tAAZNVLGyeNuvzDRUwT8NBXNHI68cAvhvpq1HoTVXn85sUnQBXhbSzrB5Uffvn3Fr
fxdVSXvg659FweI1HKCMOvt13SKn8nEghQOlD46LPUnjoOQTtT9Z69Oyo3E1bOrC8nU7RB4S+UK+
ASaQvrCd5xJAbp32lIQqPuWXaKYlz7ntbNTY5ZimFg5JiLrQuXLWLsm1ouPWt2AZa3eChALjPw8h
3CtnbfFhsHOYpaiGUa47Bt8P8SKMEpGJu7Bv3ZiPjF53uwHxcUEL4U3B6tZYcDRLxs8CXZXoY0EE
qtWFZcbPaPj0+xAvqWahe81X0D0qTKvtb14Io8J04cMAsQgofCAwmvrUUH6G5TXl48VMuOUxMEnF
mv0cVPATeYyhrWK7bmUbfr81OHpviXBjju8SlH89kcal8OXIFhwZ9Y91egv/N8g94+IU06qPxYJ9
3M1yqJDt3M36miL9k/BudLUYw9Ya0MJNibCoX69yjx6hlnRASQTYTMqbd8xVMbJMmaXhishS5UW8
G4Sgcj3RKw7IEVBxuCqQxDL9mwopHpCfdtGnnUXfsuBWEozVdgj4DHfL7VEEiZecao30KZZtlyKO
wAMfRuy7HcKr8Ikta3NpaOMT3etfhenWGP5dFUzdss5lJWJnFxE1L2rsC8LK+lNOeYaRmxzUAxjT
PpA6AB0dXZZYeh9ZwE0IimHrY5CgcWeWxuDMs1PMn3lezgITduK15JrjuWcPTiFrGw9LINpAsIhj
rc22MLFFhc1A3+PASrXQiRfjcfQYCFht1owipLWAPKrQfdfsOpVNl8S3Hrl+Vgp0leiCFXsDlaHD
wQ2OjugpgEzHkN/teV7JnRpHXaxaDG+bO0uyzuJmbMBjxVwL3lv+9fyCBK4zZAehDEEeW4o9SDDN
H1rabWip7XnqG4WFRUqOwOPWy7zrrRNuAqfYIHwS5pjpsUovwuTP2QQPZMMDPUpQlPita3o/34LF
Wb+BgPCE4yvum9t9aDgGuVKcYkC6Hzxl2wWSNLcJiyhNfG7/XXzvun2KobsC3ImaLpQU6gf+MNvF
x14tej4ZURf5pe9xlstF9tQgZd6YI8P2fxu7FWnVxkYI+3RahOdVqR+eD/4+lptUnM42NyQlBLlk
mk9v8GL2Cb3ab9mQRxXTGt3DnQIWTyrAbR5CleqQkpK81oiwGdrlBIkYu/dUp4vgcM62Pmd6/GmC
zfgX/5I7IEM2YqStJZLGqa769HLIatIf3grsB1CDSVg/6XIs6QbJ8KVX0c7oMQV3KY/2+PQB/KZU
pJPZRRCJHzYsXvJM3LFqkF3YYugqB8kbnD0Ty6UXLE0u9DZJV9FVZCFdTQn/K+XYbEnJhFichv8N
genCagEXrGdrjANQSrPuZaKQVOgkxEySTvA8Z6tsMQ+wKTV9ED45M8bTLN+APKal42JiU6mGyvBn
4L7/yCwCBINMYr8xZ7lbtmSn0QHGUwn8JLwROjcZVy7HcNZrHI+D/BI7peppEBbWQQxSf7xLFTVx
T5mge2rYsx9KzsKsjOAc2nYaVjjrSYlEirkbIbA339LGGN/nMaGF97kYY5u2offIXlggV54Jzg9M
nf23CH9ixuC0Jdr+dIQomUSOBuLNmWqweDUcnJTxkkYpqDiYJ5QFsHAPokD2h8Ox128+/Xdp5Ns/
q8ZytwZZiK5fHGEMrjQsaff80TzXvS3YM1pgtZ3IPkqkfa2DSl98Lkn55lAatHOzktfQYZYsuaai
ZOJWCshy+iZs5uu0LiZpj4km8zgYQ6bTy6ULm15Ek6JkwXufPGdRZHdzZLoyxxMPDx7pTlc6D3YD
tVbPW0rVKI88WzduopmBWsZrtCHzn+nfoofggG6jX13Nusf86J2srSd34I7+CRt7uxvEWznh9Heb
sSk0dN9pI56Gt+UvsXKgj5em2sATwZjpGTBCBZzdhBllAt4xGDYQd5SKHC9QrJZYMnqiVLIG94ph
IAcscYREzRqEv37em+BHkQyWmp018lk6Ueg0oYTZvlezUZu+PmJLKH2UeroC2BkCgxhmzLqx9Dvp
6kqNZRYjCpI+EH0Mej0LdHaagyA9TMSBwycSuMz7sgI/yn6PMdFS0Fp3TqwPnpNn2hLx7UBOkRKr
J9Yz0XndysOA1+9t/tbNonMGGBXdssgTqw48oHVk3ZDFyY8+R6TOvwaGeQiZWWf6cM4cTO/CN8GV
lg5v5ZMXv0osdhQ51dzONulsth8So/pdSJOsanOG8KoXZ0FIJrZEk3LMkrkuhn5hkM1fsC28XX56
bqUsMzx+0Cmomv9SDynkmMxIo4bZRtZua2kObqcdhmDaKEAr2Z/NUJKZ/kMpsuBucTxktfMJdP07
mFfeCowSf+5c9sd6RwnHvyywLcRCsf5+UrkAwz0/b+1rk7JyLJplw6Thmv3CQkSK62akA9QH/kkq
042HDblJF9YhACMrTxpRuWtcPfkjigMBFvVUDcQjUDlnzTWByKB9eZMOPfjBii2dhZOqnT2ngxN0
aed+V1+kWW4parztV/5hm1njfOWh8Q79w33p3LPV5NGZVzutxYMmQoMiUNk4ilzyO2gaCyWCrlTh
5qo9AGgUAKbTk/cn1VcT0t0rVDGlKflptktj6aMWsZf5D0xFAEmv8XC9rJT1YVoTHb+qiQZcIgpV
2NdEGqEcnrKQGt9PiPZQqKdTtPOUkKqE+JXxtD/tmL2E5Km5H7HLG9o3KmLPry9YHq/sWWQSGeaj
XKfFrUkDc84T6ahPqeYOueREhblOQEgMCAdA9ZmOdgoPwwxxV3sDFwe2sZVR0nTx84rhcb0hPsFk
KEiVgi2ZPH0KG2PLPn+LxnZSBidSlsKFW3PaoFFVv9CeBXwcpR54oEhcMbg6lxhevL3uK9ZqTRsC
HjkFJvD5dHMI9mTlDvx1GmXfWXehi4cCWjs/DhXw53y9gciZYYETZY5Oy/nrCNNFZNGJ+LNbE/+U
8lJIdAFoLOlGVQnWWHioUqOHM1D1YUVKKOzw3wd66d+c1brOB07jdNFaV5Qrki9kY0xb9PKyWXt+
Gt1nPgPb1RfQR+gbqS+0W8DZu9yFHo8vmvLMspmbG4lNhVSmthvuyeyFXfZpqFjK3zqMa3i4zvn1
nDi7iAR2Fe0YGYBzbGs9eLcjb2NcrCRa3Ob7SdhldV5wmcL4TVeVk0t8i3sKQd2X0vmecC7hUM/P
jVfJaXSmRnKxLWtQOe+UH1UL/8BT6xLxey5xzzBsuOeEE0KiRzg6h7/17vc1bm3tXoKjcmFyI82N
w6Bl/G6F2x6MWSLUkAbNj71GCPifRNZfbG3YqAQPxgd3EEYT3EVQ9r0y1vI5Cxgzcax0A4TqUbzq
NNofTDWh/18FrWYj75Tv6W/OtkSWh6x8GZ923w9yy3poYDnvoDUDrzG4s6BwHhPFWeuX/poiGEbw
pGTk6ZuVQL86WrXQ1I4FehjZ5UUiVEfpu9ZzCLq1z4LJ1GqCYwtxl/31tOzT2SOuIFq5BvKcHIfk
RXTAn6MCqkYTlAffT8W6KGj8EjIUbKcOWQunJ0NsmWuHJDhuO4DThrJ2ZxT7hfOEon3KM/EVgMJv
VAxIGO9uSN7/S2/kkD7sL5BCmwxFQV1cZnipc12ltpJ2/IuQLDwkwjFy7nVGEdeKzeKfjyeOWMzp
PKJiAXjr5QrB67KNn8Wxjg0ckWjQ3nUgp95yXiirWncRb+YzSYv7kgUCixFrWEyDA1CQkHqMfX29
Biu3cUwd2OtSyKrKIAl/eOUa/0oOlSe44wSBICdNtW39b1g1/A91I/6rHFiQcx05Zgl16Z0bDqqr
amwuFw/4ra4PRiJZJOFg6zssZDjXdgT9mwY4/XMWcfQgCthPV8pmJWOknQNaPaIQCJ0IuRjhROxS
zgKByFPI2pNvLkdPw505SRQtE9Zxir3k9EV06sNdQkHnvjy2luTvczAs6Y/de8sAeOJncLE2vGio
I6HpVqnKFcaKssleGMMILqXaHdjt1Ya9BLFIV4QVBiRY99iG5gbUWouagxzdMXSvi8lM7sk8DqK1
Lrg4x7inVKk4eBIfwANJdbjsC390QKi3s0Det/RLXiczGDeh8esiEJNr639u2xK+RRg/qEQbceZD
wfIH3WK0M6BXcFfz0npEhtegi6IDFaRqVqrTyh0JwNmjCwl+UHbJgWqMBZwYWXPA0Xz3iIRPO2Th
6aScPVX3F84P95v2/nzisgigHUVqkEr1xMD0gLgoPRjc7CaX/gv2nPJ7j2OBjOO/AfYZM6KULo4k
5enNNT/4TS5XBDC3VZE5+XJmdZMyfcn65zEtpJLrzmVj4pwv2fHgRBazwfHTP5vZsnnbZmurNM94
21lE8nxVUCapnpuwb/t/b4ZifVHNkcJD7zw34w/KHxUGHkgfMHedaxhksjn4BjO5WQPNJA2v72L3
/G4cly1Zb2JhtoQVRQLrACZEsnPSBdpR481rOgkCX1j4eXGVbt9boGGVVq4fh+A7qKtfd2cVy2TG
4oKEKdxM1CkBn89zf6q8teCD67SX7qPjRyggbL9AccAqgsQJKAZEvmPx47EuF7Bv9JtxDTDpyT0F
TO7hr45eAXJtDWTGtKu9pBXO5whv/xOu1ipNaaBgZwuYhoZV3O/0T2rzyFqwvIxM0XLoPj5tTVMW
pHCHPq0sKgnsT9m2XbjCDgvr/3owI2pP5ZmRS8sfLIIztBZ4B0xyt1qOB2WRg0NwnZJ0DBiQngvb
oU60ob+O2tey+NsCuuWfvvfEbktKHJsG9b9okVKhuMxai20p5kUUduVfULTDRtSfOlOs1nAhudST
7f9OtDZtkx6MYeXmVhD1NqeYTR7Tvj7qF9MUg8jSRJqQOeU49YbyHRLt+WM2MYIFTjjmVEW4R+tx
n65gEG2PBYOiA4/7Y3Dp3MocKqGfhmhCnK1If1oK00IZf7RmJwxx94oamlHmDNhxPO2aTz/VKWqK
mrSbrxuhbRHcgTBJXxy1hGOjDOdGSt1E6SzdG4+YtiJqpW/Hd0vTUClyAi1mZ81lvxFADD/8bbiw
G5gWEExfvZRoj4Tubv2/MTEmptxW6rc/I/WAbRsAD2N9vAiMAt5Zzoj2AhqmgLbiT4YJ4sseiLyz
r61WM7kZFeiaX8a2ForCT4B1ZrxiA0GkhFpkYhz1vK+uuRyRACsRxHUdkCDZgVB1X47QKRm6/tX1
xkq/1UZc8kpX5tqoloox29DakXJ0fmN3tm+qwlv/7gm8/PAAYqMaBJQLJZ3Qp2g7PUuPKY3cbJWb
Bhuo5pgrfQqBKW8plytr9TPTPQT2FBipxmW9/+NxSNAgij34G9mtxpLgr27nUhypKg8VmvPsbt2r
c7bpd/RarK9LoPqc0/JwOKjQZsast4JOdBQyXRfdUzntbjRH0aYYHtcyp7bqzZu3fQkrrIzGnw46
c4xHo5xsQ2G/4YFtvbN/MOQoXvlMoQctRVlZrzCSgTJQjPzXD6lLpoT60w0dlBDi4DRJPK0VV3jO
m8PeNlZOUySdIL1HH/F+3SG1GE056aNUM19e6jgEwjHUOEf7Kb3/r9A1ctCgW0XFS8Tvebrt+DnZ
r3YaA5t1EDz2s3ca7CGzCcq7ULfmJdquhdSBFoKFNPsmW3Dyw03+BjJd8TLYvVXiBhGrdlA11LyX
gYySK0yooBxa1M5Wq+xvGZnvp+QuAXwXWzxAMMOlh7D72UmHbNoofCYj6qwoUa1ht1LG147JzNgm
qzHGv2NfR2lsYtLeszWonDrGJU6sUFvOIyHPs9j+b5JTl8LoiMQU9X8ZCSb9u1NN/Qyyu2UUf+iX
BvYt0QzYHKj9Dv/WJbOM3iJPiLOKfMynYnJT6TN+zz2ywTCBir8bdfDAh9KTm2zK5llf8Z4XtsdM
dFf200Ujsu28C9UTAmjNTHyyIibInMJtVxIjoYaZAvwxST8dBOte+ixLSmplE1PvMo+hoPyuTFUG
GzzFwRDiUGAd1ogHX3uMwmQ/TbO5Dgy6V40fxD5dJixgOJNMaLcsTfOcmIIGIDIhPb5xLYtDbieV
IHV9yL4OKhH5ckbO6uUT23lv0yIaB45RjlRhMKrLRx4aFBuN69bN1R0tBpPXIJBTM+LjEUBOD4D0
rDS1XCCYTk/XOL9Tlt83cct96BFaJk34cly5KDdTdprewA9T2bQYtxbYjR94iodNFpAzaynrbCaI
6zUHGHTWJEdc4htSvTEIxnEFRuUrLQJP0gX5VEOU0DjiMcZzYRPz+NsQzRrBkgidFwmikyJ5bJZQ
Vq764hiEopUdGCJcEzwFQyZN/tKOnFkzN4Q5wISeuqqtW9nWSSwEhxccFL8PrI9sWcCvbMA3VJms
E//irXDtR81RXZCKAmXFozs3qDcSWMN7VRsqO1OoenyMGPCFC4c0z6RJFcbCDiCI9C7k5BBV+50O
LK5Gg6oVORlLe9WEqa+OiC5Cd9eW1TPrM7sita1sWais9xaUNsLxYoD9lb5l3QxoQYYFslsKb/Nw
/loCS4l8QvdhQBFJciGheMyhPdsbpNKRtG+lYV8mYiIecsQjGzzXVfTX2lSIcMFUcyO15vNXio6P
1PYNUlVt5ZpsWiegwA+ZYVateI9pJY0vvBi5NZGn0iaexlNfSEmg/K+RMuH4TrjDvTDJpqQ+qesT
AW4eaS52F5w4sK5YApAy7hbZeVUrjNuqvD+pOBUhq8qeMrKaUZ7pXZD0CXZiOdBq5hCviYUMjFj9
pxZAyMR8CoZdCjgrij18/23uCw572qOfNodniVWmEbpW8eiQUgNhct22zhBZswCScosEYu3wCxTt
RjAIGy8Kav8Y9h8IZ5/9WnMF+Srk8+saJF3vUTvXzDRurVEJ/UPzV0F43imx2Y9uCsoIBdmHsPDZ
PpLp7IixGAUIS4unL7jft3+mYpyw4G4ic/XNpi4bFHxnX29DZ7s1Xy+1/+tdimyLqU/eqfGIzl8e
qlcKE3/eEeyq1jGw1fn+rCNIyUmN6SrM2iPfdYspi29C0PAGeqqc7j5cbrxyD2y81jixrScvrkq/
JCqKnaPDPphMadeoCVmlDoCfdTdPjEJJtuZcqrU0Jegp2BJEjTa2GblRrRQsVTHDJhw5oO4Icmn6
lhJ4C0lUkk1KkUfevpf/JNu3ONTaz24LKRP7CpU7Gt7NxsuprTJ7rcAnUJDUnFwgq4jDPy4Nrf0E
1JlPEwxI8oz7CbQlT9OttjIa+NBUfcjD/EpU/FD//ulGx3n6amT1xuR1JwRaaFaSRUPuFD4UJ4fV
OSqlNo2LdpBIZf5hEPJiJJczMHORQfxczB8zY+Bs+MOlzYLli2npshOGCnCicvC5Bq4FcXqm/j1K
4DbBZgnEodBzlT4hEkcgbCcK720/RYhX2e3NwioDMY8fqci5c5zSKmR/ORjHohdTa8QGlEVCezOn
zPe6TraDT0Rt7AX1LLcImjaK74Cosv9Tr5FQx/wYROcvcyNtgGy0lpArMXSDX4CPXxT6P7ZqhWow
uYZruAO/24hoEkj4tbl/BHGVtdXR+FuBEAYCTSrZtOag8rn9C9DL7Vj2bitQRa+4FZ4q6joofaZB
xPjgdqCnhDWSsq5Cu9mzR4ISNt6PvMGVxIAw8h8gJhzu3mIPzJkDlB+g3M0YzREvumUc9wXgqSSS
6TjshDe9J3Mte32T5eTQumlzgitOIXvgJfjpJgpOdJO+ZHUnOknyv+246Q2a/+158Ht4nTbd69+v
jy+nkWC8yHOUQFCiUL/l+y15wJqrbMgLxr98Iwwlc3Fn7EdPpMttkLN4xkTf6B1DbGam/s6k1GVj
JHkoGSOXWx+j2f27Oxg7CMZzu/cPD8vE8JZZ97mmjwvldfbuYONvPMkD6iHCsHd52WDRoT62IGmO
mo29hR+iHgGQ8qTDnd+lCT1mMta3iLop1akjiPvJl8C1SM7c5jEfEGiqbLt8nS5fTfpWby8Cw/cM
VMrJZub8n7HM+C/t7byJrt9oNmJOmNFmaHtbndVgnFfyQuubdvsMhuJs9slhpe1js9EGvsPjo9s/
6Jb4395GV77ywO6D/y6qkt8l5oR/yPcDgZOpQWgP+gxvn4JxDJdbWSgsjdkojyubGJI5oIXPQXCi
nFXsNIS7QKzz0+QTIacLZUbvj7Rbr/5uhsxxFf/mj971wOAifsLNcjO17Rt7PhbtcQnBAdTpyMC4
qA5q20mluVjs2c+iu/mx9NJiufp2blUVKwFM06Q8xSPcUdFiLD4vZzhnX1iQRmiHlSJv7OOJYVNw
NPsFYDLKTclbrEq+G8HzMdWwAk+iW67nEA+HQy6tHfPFbE8IAJ1K/r1/+j/DnMfOE6EDS3MWxPGI
4O/jbNirT+A968AxSzJ9/X7FkB5qKmLlOdkQk8L9mhiNJV1IvT/v9a8znpukXk9hWFXWJL8cPIW1
Tzr6V6y/X8ySlf+hx+4+NP4fvn/zfJ0T2m5FGApD1SnxE/CoEsiWLei1EasXICxoqmAbTljy/oGm
xA/7InbevdIR2dHIjCw5LIYMbV2YBJBGxbsXrgjbop6h3XCWPX6Ai19p9mJcxbV9PZ6A8W10fr2z
I2LHc7T4ACrhS2k1ed8Eclda4royIzsR1sDB+UbCinBGJVRoeL+eyyqIdRDyamPZQ1H7k8wKOSt2
2u+2UJCpawIcXJaqrDmXEu1qTengx9V64i6zCEhBvrmcJl6G1dvz4/1n9V0MIdIu6YO1d3txaEiC
5/M/VdwlaxxnmVjZwkcZ6T+EEUdfmAUVWAl4GbjVR7rqArysS604ORvk6txBRqOSxnQgVnehKBsx
V9yu6QjQ5iyA/olxYWJywQylR88PRBeWlRLzkoupolafyJN4+LmuzZDd0cpdjvlCQCi5q/xqgmO+
a1PH9OrGBg7AS95uxh+hakfAw7ashWOGi50D7qDo0QjjdHvZ/g5w9uBdHSviifsvDXzhXp8Drbvd
bP0pOLexvhbF2OJ9l+iRWPWagP6Y8if2N8a0bUjL2HqiC4rdM57ZMGYchYNpEbvoDUzyLaY2+6sJ
hj/9NGgv0WjqiRbDE0OubG8fwYioMsNcU5Z9VpQV6dW+aGxO3LFM1Ia1Ya/I4qrsNYNjyyJAMemf
OuLjSgZcAQb6k2kxCyQvFcTi4n6O2C+7rO35eYX5jq5h0whHnVK3bpnO65wS5TTTOp5ZT9esXl/g
KFueaDQHafVk1J+rk4mQ2oOmZeNPvA7GJhSUzqSr7BWZzIZG6pMdLTEY5LLDlVAvQ3TnMa2/6Zcq
gkCnSC29oRFztTSHbG6mK22/7XOaix1zaxSM5UOSgLJ4GkPP262HTkd+YBZgBk0hxDbQiQrlAAwJ
/iiu9YmE6JUWHYdIfmZB76nX8zeMOCs2vj5AESGE6LS6pWAfqKPiJIZO6TPdnfJ9tJYuvaX9k71n
Pc9ZqEo/gQisEw2e2VnYLHB+Ib3hZ+SBO10kYj783mR6uLekTwCYZVNrnCGSiYxQilJXEXod2Lk/
nDpgrXr0SLHicfZ6xtVGE1jMKp+MIczvWzXOPdSLt7bG8kW7CZxkj/2xIr2mgGzAVcs6Mpf+kAvg
oumBHcffRTzgxViF64O6z1lW63GeLpecGGrEkzONwWg+62QNThalMlxdutPsTNzqGvSumJppo3Qm
7orig1sAECflHoJJYPi5njse+AEs8y5giMJEy4GVCJXPjbpdhrdir4JUx3VxWHK+UuQOal70MR0Y
/KsqPcoIJ5fg59Ln+ps425PcAKrxoNjVPUGNqGRK0Gr6ENGuttInfRQ9CLWOzcMIbMciHY9ft4KE
wjqmUQeN6o2/LsGMPe4D3QD2hl/yp0iVCrckJ/llxPk20PNp/E0haTKFlf5qrS9PagLYjxULHMbg
LPtg3YW5p4iF0dNxcKIAbFq6GTUeeqO7MjaQ89raEHpT6vKnlfa3Di+AXfyQsNLkEzAm9FhnpoOr
WDX9pST0czFVLGsN0pU2ujY9TILe8wvnlG7L16s4gyrr31MlVyxXddVkZCP83DydpMbmYMryXyr4
6mVW3202t41/k261g7Bi9Nnw7IA4sSkolBMetetk48OjJWEvc+E1xloyl8Ng/OrnSubKYQhSIFtb
MPpZWKDX8/vkGRDA1TWy49iHtUh89WRVe1ofripmWcLTHmy+e6jsyKSi+1dt/3MG5jcs5mrOZIWn
HBvPeedxRw45ZZrhnFdxA8jyupzx7SQaHefFlMjuHIgqLYYA13Zb5nz/XdQXrOPBhKTzkjw08pIT
DzOieIC0Rw0VColmZi65jpyoabitVrcRd2JzN7ybto5ezT5njUoHPh1T7fTkNJ1UwrzAYCUOw1K5
cfJfhfQsbraNAxTnTQT9KPxFNZqiqXcOSQZbiLc6Ub8goG1C8fL56bQAsu5hcopSnjPGZEEjw0Uj
heCr5NCYmLzOr7IagaOv+nNVYY+WFIuinSNNo9Kkjj8LHGK+KrPUWlWrsD2SJXXIR0YpNsZvtFqC
LON0GTKtqRboplOtO/SUFas4nOlPyHWsS8z58ExeauU3w3S1VQCxyGs+LDxi6Pw4JpxkDEVLV8Tj
9klekLBd9qjgnTLYAe2RJSiz2vvni1Pr5Q6SITWLkTH1uPnTeyD9tvkBGwoOD99wmHs8XXRz4Yj5
VrffDJGw8yB7ajfnRA4zqdIiAFPQN5vg04HqkH3ofylUvHY1DeQOcIkNDwwrJHIUXjTsfSqfIIdW
sqjFwLaAGqlLRx9VML90rpKwrjPNVFJxVYUezqY5OA9029/ttlKUIVtX3wXMKaa290lEr7E5hKSS
ysNxkBsUFVKfhZpc+USMsbV5k8GruDXc7+IEKCNyfdLZuUyfd7//ggIKoNRwwTRbsPik9qzZAoFb
eO+t3IokVqkj3hSBc+0+f96TUM2JQRmyfnXRtytE80RxnWu45W0Nby23daj317rjd4iAlLeTSzHr
iraZf76JUT/t0UMZOTLYGKS6krbaqyzM1jrAySylYC6gUKbVt4gOSm9iuw5mZUHlTC6xeht2s1cK
5wJfZ/8dAOrDVyJ52klSiYaPwmsaLDeDsoqyFb0FzTduPCX3sGzyKDOFqLdYS+lkPbShS8XpAr3i
VIGG7xPiIj0JL4hzXHZqW/PlADtrsF9LIXZr1ePkZmkUYT/228hr7GOaGp2cTPS5vhRYJcDhDblw
otjabHg7xMqvX78Ppk0ZJS9+ZxK7v7+w9th/zqkxdb5X/CE9p0BpxvkEQaIDnpAtpCn5ykbGhoij
TXvV719INgRXCJdKO698Pe8nnqGXEf+FC7rA5BT1jjv92eQWQUFGrJITHzbvCVs+MnKSEt1O4z1Y
5vJXDgBb/WFitmGv1yNC1fdMUfFblgXPPU1wqjOhd1XDzt+ogMBUW0q7Un+gXrE/mIFVK+1mZo0R
V3L9P5UchBAzIQ0yPmqaMj9r4mfjWbr5KRlFUXEzbUU8otAJ9zPsO4k0rBIw3M/RNh41M7iqtarD
adc0tdUi3dL2BNMk9AEnx5Wij/quaYlh3YSldp2r3RdWDwuUiEv0tv4VT3cGyqo+aFxET9QnQS5L
p1l84gigWNii3iBFal3QnTmh6YYetARqnGA/taIdUHoQyc/qE20Q4yBcloQ3aLwhLX6msqRuYifU
NbRqhaX7sjpgZzQK0oVZIrkOZd0MDh1g9V6rkyq4m4B0XY38ER15pWnsKV+VpufJEhhE4fVImVC2
BJvivxPIPevsxTAltVt20lS6f+CaFBb8KeIJfn1TSptQSiWdO4sC0B6jQ0FbqpDCzITv0kKwqu5w
6TgjHi4dO32Q/L6GuISsk7R/7DnOcz0Bh/qttcar3nF8640VMzO2UUXflcYNPZXuBzFaH8UzemDs
p5WjIsrxsZScVLeupM3secZD8Ev26UlnOvd/4psDnwU53MYgAHRLYDWw/oMm9aLjQ/EjAOWw40Hl
5kjqDCw82VW4M+NB7/H04db8fNFicmy6+VzgAlA0Kt55GCKzQT9peK9nXAcbpTKKtt72rL84d2tq
30q49l5TPsjKZBETvuT5GovIisnPqFjSwD1jNmJPFVD3NcxQXvz4p3ED/1vL4fEhf63hgDdZ4ro4
2cX7RFykaOcp9/UStzAwtk4RN2/8rLdpx+kK3QXDJvvT5X9lxB1u77NfPXQc0hPBdQlcgEUtyn3i
0hQMtBcQejuPN4DUnaVl0GhvyBa7c+hpkeRa+LS7XbYz4TxvcL9/v7TooVVEnWkE8cCmNHI204DI
9ZMJE2N0oZxjHBhmFQyYM2eAIE9qJTuBaKM8z2/oJSdkPWYoPR+xRQHROS5LCIRAnH1N6m9JH7++
sU/X4apuSm486y0islBpf8OTWWdVesSw6x1egPWTZOutjyQbNBS0UuOrBOZHhhdl/x0O+625io9o
w0J94kXdvp4lodMprf6WGkDlaCE401J2nfHkG5WUBRe3teVVQ0wHqDVn9/gBisDoWdP/j4QeQrx6
DfY+FUBNS+kv8FubVr0lM9nXzYJd4pd+6wFTuQ3apSETyX5hwTDmXUDYKMG0/Dxw6Tf5nJ4HjTHO
dQiZXPPC5a9VNKQFrUdx0VwNozVw1nxDYrml3AFqtGFvEgjMs2Qt4akJZy2Zs3ygx17q2Z6iN3r0
6K92NaK2XAdJ+yqeax6aLBdI96dmTAuqiaoyHor8mp19WcAdA8X/4ui0e/G2D8prD8sK29LW/0UR
n3phrb+A+YcAi/clZdUuKVl2qKpsqibIqIm5Ja8zhFHVC7BK2J6J2TLGSiOnLep/rWd8/vUX6NRU
I2vjem5f8xJWdSUneTIAGDe57wl8MM2zOTXTX8MQ4nsCOpHbMqdRplMBZ5RPKZevtw96AmZk57fK
F6rw+upbSAdo2+entXdpRCfwtpZvLkQJuRtgQIQ3pS3zk9PngBdR52963bpLHi4l7wh5IxOxWseU
1b6jdiLCKLdj78xYw6W+FqRNVKQq6SYvlCHav5DVJ23EHc5yvq9b9CeZjdbOso/1EGHjMuyoRXHV
ffxJGZC6X7qtWmxmhRSLaaQs23Nn7bRtQ5GI9xBtV8CNeSRLlF2U4K7nmAWIK+5au67b2nR/OuYJ
sSGyF4cZIicWoovlmE93C0DhuIewLOTTC6hTHMLmFFS3RBC50qM+9hihNSqf5baHCu4aLdWyHOdF
BSolCecEPXh2ZCnLRZmi9BcC5B9+SKFSwnz9cD+7ajv3X7VdqeCh+J3adMhHFm/XXEWL/7Axnbrx
2AhRbWP5SxKSqU8WvvHCVyicPN8xo0qcp+Cj1QR3IdnKLiPVEHJunBxpOfZ7/EpjlquJUQmu/BjR
iZmJ2cYqjI4OT2bieVZgvL6+xD1AMujyvxdBZArpo+vE58ViH4INyyIvtuDqoNBIkrKS2abduhwn
R8P9gGDiKmVhvFbIxDTT+zt13+9vRX0kpFiBhK53siGeQKvVqp5bk5OECNcCXqvibh3tBX3HL9HW
/xAdT0jhmBPlLAcqM0yAC1S6KN7zMW2GrMj7pRBhRbVoJo30QYqNJn4QUUSn7jm2EiF1UwbJNOpb
UuwkhZAkp+XJ6StJTwLPQ0PXzu0d7yA5cu9ADXP17iUUrytkCC4q4f3CJYrAQDk1uvMUpLAkQVff
x/8v3S78HtqCLCmsFD4deN4BCS1nRVAi8xgIOwIGkq257DSAdN5pRGp3APu4OItR7TeNNTiVRdlS
48+Jjjjxd/WZt+bL3+jk/xWTpxRf1vHXNkNLwcU0U85SPaHbE1cYE7B9CWCa46CLpilLF3WuEDah
QpwNlfkpfn+4LVgkkTxAd5C3CrsWNcAafFrNU++hcj9baLZInVoCQcjSY8Z95T+PeCfYbfL5Brj4
CDnMlt7C1fF4iK+J0pb5C4NgAVYBIJ2NC+udFgwD9Tm1HvUCjBf+30lx3IIWdfNT8bJEb14WjtQf
AoQCUj3AZADmqucQJiQbKc1NYknwcFUFWmJHt25NanToZ6CrbW0yzR+gHou0vWW0OwzdmDpA994k
tJHmReQYnGZhv61J5VcMPgqIJOZEqXcTZz7F2BEyw5Qd7hUDixmYusUd26lONU+BtDJh4YIMYtEp
3pxnSb/qe3tmzoqCNosgXTWfdvMczKUDALNevbnh+4C8TTkyRPuEdJmdonge50Rstp3lTOWfq38e
ShC36KOw8gD2WnPi/SPibxkAalQgOT4RuNLiX01EBPmkDdVbjXtSq9bZ5+4zDsHFacJKQoFq7PUf
JuTdGiEo68hVCz8S+reg0G929r0LIpNpbkL/l4xtd9Rjln7/tBxiHXYef34QcV9I9Pc3jFNCMUdt
HC+73K7+bOBhgkF48bhM2lpA8N9jrEgoQm1Koy9QdPDVVNeB1jRz7N2+B9SsTHdIeX9p3wnaM1hs
fVsoFMiD1iWCdcEWBb2YBhXON12+/FcUjatcMXsHE6Zo93f+3VTggEYShdpTpIaoHtJ+d3CK6YX5
Byiu7xDMizWbVA53hilBv4Ydaw/9togyQ/XDHkV/aanft6+5y1T5NtS0aAyc9bbjboZBOx7u6Hv1
uZyjvkbt16b511Ay+okkAeAzrCWwr2boXlfgzlhlrs4aHnkdm2VLvRr35XVtfdsR+UveI35+G6bM
1nrYr8oCUuKHbyJ0r/RwZfJxI+nra3OkCkTqgiLgftbS8B9XRFIq/OiLhT0GKUmL9988FLiKK2JW
LiEPhDoryfO5sgDfJ+rEG0NiLJrJnl6tz+sDV+siIBu2X/Mow1PkiGMjIhaLkoJW8Cm7dYI3ALX+
WI0IfeSk4unr1IA4E1qIbXwHXJ5eOHJstZR+HdP8B5b/6Jx8dgeCUtXyYmbgHO35ALEwDnHTON1/
cePcbb1lgkgZtRq6calvjVum0M13TlZb9a9vmbHHw9XVkn568iqAsJq85zcvqrp9eWkO/+zlfIoo
GH1Q9EhgiFf0ODaYyUM4yzaWXNwrd9Aom3LzdPgM7pH+QXFGHmw+UISZWdnUNDBbcPafegKMnouw
hcel38+O+xlMcSpfP9Lq+3pxm3AxQ7d3dtX2YdUZ+xkMmCO+LaRJQ7K/VxbVL4Vq1p2rP3sfCw5l
34jtQIFBUJpKjuEJNY9i5REufTQNTHDP2TsG3vKa3QjG7DvZaoB30Y8/OPpNJXh9T19JBDNSMwed
vgllV+abj/V2QeU1qVQHovfhFvS9zGlaq/xfUuq8wfD1G/Cr8JcEw+TLJ2wv2ykcpsw50EmqHaX8
WAbC19zu2CT/dgq0fE7CB7X6lO6okHM9ZM6fFx6yPWjiT4MyLefOrmKTxHaCNN59MyMJww7TrxcW
OCQA07qWWnIyzIwnOCrMq5FVYvLlrQnMXC4wZOjSFM+40afMPVz73ehThmIs6yqaKZdBLhnhrwFp
EppEpdVUZbMgQ3IZkUxo1lZHzbktkL5DP4xWcL1s6+ezEaTpU4UZaYcSBLG53CJiOncRaRqhXDO/
w8yyvoJsNJuRlaAMWsklq3x4Kt66Supi0GIuEcz2p06Syeytt2tXNR1wQTRANYmhzNPnBiJB+7vW
zwGtAE9tHMbl6v8M8fuGqtUMzbWd+v4v9adgPx0utxWoRaVKn4+VDx0x9IzwGBRL0z4YyoJVWE1p
UjHVRvrPrnnqBuIy3bGwHuHPCz3u39d/QOXr3vtDROGo41eevb8MlD5XWN5W/pUg/H0UvXC0Fo9s
d3q8PaDDubyBj2s3OmMG8atLSVkem348ThuhGIISpsJV5gackoTkI6dBz0Kv0MgaMXQ9mZp6fd0e
hrtdCpKkJxZlIYmOdWyYZRf5DrUBPwe9YFvn99t0shIsJWwhUTcdS3AmOqrlG82INgNtVzOCzXQe
oxqlMH5fuQ/n7SJ7SvPA7bp8kUQ9c4QRiDBSigM5Ei4t/7mQHjyVtc0DcsqjKVYy3JYUv4luDdWG
ga0mkmQISiIxT7sZz0EG82aXzT5fHng90Esz51c62lnnkc07szA3TNxK1nYL247rrzCXCMOWk/hN
eicxV6LnD4ZdlvDSgR4zRtrVpWZDok1VQyq7hvBYGau++SW11P/dFz8H4YTEFCTwhuMCCx4OXppH
1HDu2w2L382HrZzoueuY256kPn4axqpNCU3po9JhdgO+DT2rA5ibK5O2tuTq0JlWe1/KbXzP/3YM
ZhKCDlcvjSpKz3mZLFExU6pGUiZWeWv/ZnnW+WEbJ1zlNrctZNUSQz+yyJOcu5SdbNdT6dqFdtr9
lUep8Dn0wlGav7hDSyaf0BIZfYeeklQHFqmXV2DV0ti9QxwHc6SwMZbolGztyyMK239DKjKZajmr
PBFjNY3Fsp4COLxNnECCwfWRw9BDDOUYSfqhYzQJbhw5xo8h5XA8JF2BxYvU/pimByxETNBDdftM
MmnXzY1pHdJWiFTjOEkHmU4SjG4mSoQAd2olot3cWg7jidBH2dRVm64fXDysvE4ydW3gH6Hof/5m
YdofVcAvU8q6gFz0OgY7BAlyoRyFoFwWyl7pxjwcBNPw8+3h3/jEORwzl4A8ET7j6q4A1BVMABH4
6W2xAhKbJlrpFNy7qUWmZrKmpJ9hYhv7rAOjDY7QRShEMqkUA4WHjQkTBLNjqRUtbhgeaOGkjc9A
ED3JQFovZ0qiiVyPKs1Ha0oO/R56ql5D4nTkfoQz7S82wwoeSbuusddpWsjCL53r5RjJYXIOJTwo
Pghe89f1foj/jKgQswcP2xkbQPoU58fgtx8zxoW430k7oEE4UZJhIpuYJDEnweQiyh0uh3ghNZbQ
vKdVqIJCR1BPId8FONH3aLHlxl3g2UM+qQtsoUMX/byQAtlabo4bZ2ekG5YbtXX723oOqxzF/Czd
4KZQu+E5BbDG2gr7KkX9vT7F6FYdiDKh1mN8ztfjtiZcMqnRzdxYPt9smEnW2TySr9kNKHt4dvje
Ztgqssb9eEwxZtjmVrbpH+Cd/GH43EZbF0qIAka2KmnTpm7Y/v11viEBAKyjEZbzCVURnjAiBmGY
NRTUT0m56RAvl+DvZgl8SXW3zSryLI9ytU1pGMqrsxTWDmvIaS7TyGKT+Fqy6dszL0OlGuwIDir7
oAsGZyg+E+YO6hV2UFYBldVDSFhRMnNRiePdfti+A/zmk/7sZ0i9xeRRGfnQk57v9ZJJKzHcEuL1
6jKcVe3wRoqye7h4zMtQBPQPyLUwXVTU9OUhhbnU51x8uXZHXMkpS/uNK2TvGY4NJDt4/7BKv5bY
PdMAwnhwwD1HTJShWiVb7U9bh9iVJUPCH/ZuKZIK2af35HTv1IRAHiNquSdtfchVb+y8a7NV5goM
ftwO3V/TrGPs8lw0ziRafX9W3ZZb97W1GUQx6zSBWOzu4XVePFUftjLhN+wsM0L8yTsFR44prz60
b1rTuZdy4npWCngejCiHo8VOBcxmqIXgljLBoG/6/lpulyEVyK4puzjfxSmrpI2gXbpyVkSd16hS
i8Vo6BcH76mRQgfObFSM1RZBc7JKdqy0y8aRTFQX/L3ywY5DlYq6HVAYjw+X/LxWL0hyxfx9NVuw
0BfV11/elyEaH02w+Rwi8UFxo46zzI8c1DT57Y/H6EInk7T6x7r2snhp0iVwLhG8D08rJv4hidFd
2R+cCwjwVwpvuDhGWSC1YU2KFxI7g1f8luxzUtezRm3Mj5QfzW3gu+EOp3s+LDpjQXtOBAA2I6Bx
6MgKCy7RdL2+m5pOyg6BCd26AUu2dtwhYg85T0Gv0tluYoRDH2wJBfOZja2DC6+CDU0G1BsOpLqO
dZU8UueHeiqxhKNyiV56tb09uTksLw4jb8LIfJ3InLMw/m8P5NVxE484Zdgn0WRfQErYM5JXsZSf
t8Xwg8cR2BxdxV2ETOVO+vZK3i4d4pGIx/54xewXI31f2D/3Bu+ZkKSSfBKOUeUr0eOVTtUQ6RVa
4b+OzqgkUaDStfUGZ/bo60umGh2ag8mj0PZ2HEeEY90Z+6hrOVv0n3ZkucY9gJxg85iACk0ApiBY
w7fVvKpTXvfb5dDgFft+R8IkW2iJ9wOrSndOaBRe+yvNUi3SBTf4ILfo2/pYHuS5RzF9W4Jd1RoL
DaVX7wRll7J1X7KFW580dXAJDu3soOZVp+URt1FAhk2l+ZY/ZQKwCTTZI2niyegCvj9VmcHqRDq1
P/WvKqQ3EvOMoT58Yv42P5RrZzum8T/55hlr5GQ6x8QTj4t5J16vrZCqDroIBOE3PP0Z0CzhPs8+
xLun5SljDWcJwBx5Ctu8MSmx04o2H62Oj55+dA16Dj/xV/+hqV5wBh7bVgoVVXQ9xS8gMWjge5xm
/4DG7qhleygC8JPdOKIjvkYOhvXCwf0dNFGPXzIP2oUSAZMeNGCOnV4kXZOjP7RvUmXByEv2rWiX
i3+N6gyRu4NFodmovrSQn8kZXL6/CPj2BUn99ssysGJSAI8q2nutMAyhF1jO+2Av6oFHRXWc9AdL
OvtkB1zxTCjKivOKyBBe7WFZJ7doPNPHI7pUTLohFNJswxvPLNTm72sPBJpL1PmvlOMU4fm1GmVu
gLMm95uXA/k/rZWyrInF3TcLtPPVdMJFT9PFTdqlfboXGNb1GawsBooqKq/Xi+R/Se6pDohUgoHQ
kj+wTj+N5hs+UAGNkL8rhA230caD1TF2BBnG6LEX1eZixDpum7yOGeVy1sI2UWU/bBKRXE6oTmV5
qugUMhL9Zni5ARO95thdhWTm+Y8sFMRBA1xI8Chtdc2wHtKKG90r2zqpMfWjV4qZCA2j1fBvqrRN
xAPUXQ3u2qSsXQNvcEiQzzoASv8kY0ce7WpWAhJimOIf4XiIBighSzYzMl61sgp+OurluqXnrVYc
2USRvaIAuZe52Da6Micze5wWbcnEsWwqmPUeVvor5MbS+POBymKdJmcceuBQq+Aa3nleqi8yMYj2
19/mqLZrG7Gdj4LnnUiyj2hY6fnyuzBmpmfoqDrfbVYHHpQBsaPmI44XI8uUPkxfsOiry0d5gEl3
siDC4eMAXE+q96HXL7IuyVd5VnTO0DOr9aZ4PdfFxwSnVhOPXTiW8GRAgKjyzAjAqZkQKNMc65gN
X0iwQhGiN6uk25A9lIJBCzsxk47/mz6GxkwhYoWvdN+mcvtH1IQ+9+kwR8ZkhJMBAHT7BT0gxOqG
/9SvGmv7axNkfch40nj6iHtpTQasKUdl7ZE9Cb8xthtnGDHUKjrOWmqDEewGLXNY4eIN3LkyyXPO
SN2x1+nSKKFHMVEjBoZGG1neamHUE7i3AXqmK4caRZvXTixHVSBL/KD5CX4QnjCm5+KNjnKWyCJ8
pvOyu9zzpqSSo8a2X60D6KriRXdhwTWFYRedFxHk/EfA/8sULTudOWBtX5w5EjvXox8LxBmq5hTU
GU9XwueA8tK8r9aVmD89Rfc7W4ePVEidI42S78/PQdDhO4vVsDQR4B8UnMg+408m4bH9nxkbupql
dtoZO9EDAi5qaCMvmIqyqSPeCMTC8J4fqUKdmOxDhdkdNREl+JjgP6Rho8H8BT/8tBiWReZ4cfog
cIzmoor0KW7i/CcO6SjiPn+k3qH6yBYTiQkHpoQPKd6PJPQx6yUyD+QZqwbHkV2hUPu1eH4iZpnH
GwmFKyPSsnmokXlXHsyEmqWum/1m1FAQpr+j9sfdcIHwwDA5PlkvXl6ogXN58pbgqwnXjHAOgzsD
74tB7vERmcOMig92IKIlXo4pk+Ts5Iot+2WJ3yEaLNIGRMMQ3BY5sXP3dDyNuoaW2Hl3JzrBibak
3nehroZBXw8+7QNx5/k0EWQBFv4duq4IOVFFPqV4Fv+hqhVpREPT5hTvUOOUr++/7coyjFpZUmxL
bQ80zrDQllOcQdEL48Dgi8emAeaqUMRSk6DIiKaLuJ0JJOGw5E6Fqw/SSCYAWXr8M/+OwNNhdGg1
VnlxqTscsKhPg64iM1aKD4iea/I0z+n6sKrQKPIYpMgNZdq6bxsqT06LjqrNavhZRKIBpFgngPiu
Vqabj1k+Zu45edCiHpGn0E0+LTyx6z5jD81RkzvwILRGCZk1FS1M1NQ2tzle5E/pqSoO0xC/ncTe
6Lr11TB/EyYLiLHHVUTUve4HuocHCUYvPl9UZeZ4uvuS1CNwMBu9q9hD5dn8bS0EzrQTjSsXQamF
pTSx2T67XwEIM3EmgbDetuBYi2AIQOu7lFPAxDrfuW7tfycEPsTNrWzcnuUDzDLnasrYHVjL8+MX
WHAjhjCFEzoumA/iuV+AzJjYr2cIoN51YW+CGj+V6gmyxFiLh6iuvZqjReCIoizm8h9yQqnQCjJw
lhxhz3e0qmCJI7V8RSPOVAej1NNPb7HDG3wdCPyb70e3KgueZap/uZ5DeuVl33+tVBBcdyL4Ir3Z
GkNicbA7UUk3GCYn2QOU7e4v0nVC4sksZmpIz+xhzltFmFHN/YwI3K05SXf95LRkD3RjXKxyPr6g
uCU1iOxR734jwo7S+ewK16HW/S3Zp4t/Qs8skdrdqMrenAfPOGEMXMRHaJ+Q/heAM97cous6y5eo
1XFwUnG5jQIOjWYGkTxAk4pkTECaaAxbrniMvtRYUEFvdB5PSc2TUItRHBv+sUTXo2Vt7zURY0WT
4f3Hp/pA77YqX3dFR3H8YrNqpl28fA71Hr4BRcBobP8hy6uDdcmf2p9TUBMnnIDIjS4wEEbB8a+E
3I3EcD5qNbLYWwcrdw7vLgBzxA0RzhwSvCy4+/t2/NN8mnf0xBfHUheatcYG1AM0kKAzWu8Psnmk
7undYw2yO7W/t3lbJmuhVBRuWzm90MEj9S34khvC839/8qldJJYt21ccbGPB29MZfG8wut1rLkZo
1T1MOsG+spFq/XPFxwBp19JCuiTmdbcSgqCoKdHP9RVz65hqPKgCU1qu3GCG7KQ1NAXyYHET5Abg
tjvIy1qZFByW6YVueCTJXXd3wjlJPWoIj8AjOjPBPAbMVUCu9J+L3Ul3M+WsDSryN9h+cdKDytHj
st5Y5j/E4vRpKJ01B9uRRyI2yEJD7Ezi/ZB0xfPodBfm75cJjFgu0do2IYOc1RzeLIA20iDd/qXi
Nq2ro65IOK+KZL0xo81VyqVmZSseWTlprd8sxoEKj2mUad8JYMTan5y+9ibEAGQ+LO2/9X+jsNED
D80rbf8m/kCMne6NCIVRh6X3kCARrzL3VeVPxXCOmS8jQmIQwXi3ru2UdtYJHUV1TIbYXsbYf2Kj
im1avW/WzEMrterizDlhgHdReMptaa3qLohjqIFJQKiPBbpm9T+O8lI8WDPwj3G7Qj7v0XHdyjF4
/UDanavVCmZ+VWWW6WjeeUo1+o1A8+3yOsS/Y0amrqpq2G/TnvZxZMXu6SmX3YdcNdjPnOMCTl6q
tyV12CXo133PX/egGzSHQFUSUnU3bWGipqp9gG6W0pSVvku7WHXh3FdCdJyTEp4fx92O80nFMUuy
dOVQjvU1jrj0kYaWi36/I+JM0SiO9P0T0AvHM0W4EM6YLgS86BObhx/XCRImqFfMsOTEJ/Dt56Pn
FHrbkfNOzrs5qCwTn8H+IOk3oPb+n7NK+DD3Ky4fx8XRh1RKoZhIyC9xWD/magGnmgoV+x6uHM19
0aBmZzSXoaQ830msqOOT+gkb3RZv71Zn2kYlJLVwB3ws1/1i3Jr1vQ+lKNgsg5jJTsB27XYOMYRd
jbFgZUYCjLVOy30XnJABzz2raxXb7EeBCQyqpSZHRb/vjAdMD2GedRwQA01Xq7wwaL0T8t8irMIP
Xwp5A9km73VJ/CJTWATFyCLYAw7K50BGIUPvb3mxXix26OOubr3mHIqlOu5R3I7PqWsMvrSkQSV9
v9bkEjVonjGbnXc8zNZtg4R0ixUVwn8V5yqZ43ptlw8cmO52PSFTTK055MUewcZmRfE1EfKVVFw9
pfz2qJQxaWWY3iovDnwXO8lj7/1M8Kb2c3/nMKIeXWbWu54rq82K9i/ckHo9/py8VMwh7fcrSNR1
OYm89ux0Aem5CK6mY/Zi6lE5dgrp+00EPDZdP4NFzA1as17ujqs10NTh2nWjaWeNPb4CA9phpUUk
M14HgF8ivG2grMFCvzjPmeAvro7aA6/vX+oJR8bBEzzL+9J/kKJU3QF36ZK/95KhN9NMh/qcah8U
7JGnwpMnlfvzjpCwWax750FB3msBggMoUj4bVhQwtW2AkeL0eQzyolex2TO04btkXOOrjqvH1Yfi
klgzqCY8EGg2QuYTE2o0q8PATceGRQQ6OqcQDzGMn9rlVEz5sgLcgTSaASzNI44fWPivxAnV5gOM
QcSBDyXy6JHzLrvi3908lw4N2CVFrNDoiQrtriZ2ci3anM3tS8JVvSrWbTSN3JswXIPMo+awk0Uq
09GxXqRpTuka77MF4D7u354NfzM+qLQxSIpgiKezpLpAwqmiPx5Ehg3MQsEEXOVuar4atleNuCvb
0m9ubBTfqF59tppzCFrmEtzEK80YgKrlpxesVRgz3eRF4sYYG4kNjU1J1M2jHMoxIgdAjCOom8pa
wNy58oVeif2bueCkfqlxgD3szXJvQR0aHsBb0ehMdu5oxO/KwfN63VdJcV9Iz79sEqKi7deZx4Od
ZmphEm7AHn+ULBqtYajT+iY1VJcceer+n706o5n7GUB14r1RmRVQrWDWUUORbpNO2wol53640tJZ
BfHz0s6Coa+MJzKrrBw21+xJilqSRmequu+xdImZxg/BqFc9sPnpIW4l9tzC27VIZ1bhOLpD3po7
UOuQuo6dhh4YmrAb9IdXTU7pZ8RgZrCPiq+Oue7gS+yt5c7CAnZ+gXYS3h4jwHHnpyZZeR2MbLBn
VzHrDcuIlVQJRyaRs/UZIAd62v37qMTWOMeTwPV8/74qNwer9A66wfgUCHfPmY6fXIPEpwdliqcl
ikne5f4Xpn+kizndVN3dDyxgQBjQn0ac/A1dj1bc64qVgVoyynBtUrIEjK9qyuTxl3auoNuMaXa0
Psmz5+GtaJFOmmxJyvGy+KPUZqaRPln5NkeZmC04ji9c/mtE+vllnrfnLr1Dt647KPQzQwsKppva
VkIaO4RqqSGYy4cMhVQMluYVRdWm5IGSOdCVs0TOXK4IKR6aU4yj0sW8XSt0tfSIVi80VTYIr4YE
3VylTUKXjRi2H5OXQGS6K47F4vullqK9f3xNFg4I17WtqvM34NvDfX8GDXaqBPGQZI/lVwYjwjBl
fqvoEy5BbaW7izbAZFgT8NeyM7QzXHuseBg4dgHLbRqQZR1rQCty2ose0uulc6pydp0MTu63Ncmi
kKi2LJpfBWkI2MEXZIYaNYg6yYSkWKA2A3Tdpd/aqXrsTjXeMloQFP0HTkMfTRFeR8doDCR0vqE9
zrElS/4S2g7D83pmssJMbdFYOKvxNQgMNrfmLegRrqNxgQ3vg5vjN4eXNvXvyV32hLie8VpeWumF
sP3ZnY6EiipXT3w7IEclrP7er971bbVlcJnoFV317x5MtXU5QNkrzOa6zvsbu4bEfJrLF67CKGu2
PDx/IDNODorUonDmXc5HGdSlAOxShlXBtLIi6F/XyQrrHpDIfucSL7V4iKUv5AHelCTbVl7Ifuls
m1yH+80+sBgaw0EUM1Q71x5bHalkOwDM4WpkJ7erldTehxBd7X65s9e/G8ziefWHdtO2HMjP+Jhu
QAJAcKDA6BVKlidVrdJTFP8MPqPl5ru/yv7qobAU7XAERkvxBx55kBwFZf+TSpBrwH9rJ/AFjg0y
TmYx1JHGsv9PmnDd0uzXPgzbbZO50VBYUWD31YtGggo8mnDo8BoPBReTNWG3IDMpZDWc/Mb9Yg0h
M6ysfaDSLtPd41nzWd0tCsDNxbnqDZ7Qjcrl6nZj/rVK+KxJTHXhmv6fPCh+91KNM8nkdbQh71jE
NpqBI+P+Qh7eoVsu2TtljV0OeG3wAbgk/y3mE4eK0tAs4UgKDXBetsdOsNivTSVGvFz1Hh1VlIxy
uJANJ1cRSH+80vS7gPtF4qCitBvuPJO34Qzrr41qVlajdO95j+OFTAuPcN3IBry68Hhd2SgaPs/q
rXAoBZMpekF9OAz75q/spyh6a/ZJJnlHsw0Zvn510NmETeTRW6Nsh7+yTzHcOSK4n5PSWiDNMB3P
XfuZJwPaU+SivecXBiIsxes1X2WCIenjRNDVRsuorcDteMYj6pvMW1bSVsE49SqkGDMWNkur+mby
z6cKPY6u+pFXyHZm++ph4lLyUoHP0nGYg217Z82eRNpn0zrz9RCXev1WLTSrv6a9Ora4MObpALga
epceeX8G88xZznKT+NukNmZDhfhhNYxQ0Uubc8/ebxtRksI0cPQGD+PDOugh4PkZr6HsWOZIfcxV
FTkBLv4Y3FOik2rHMy6AFG2Jz/g6SzQOVP/dLr9tyW/2z4xeHkxvDI2gXx6UJ+GccUbYtvQHWSDd
g+ZxcKTUQHRT3OPgAaQOcXO8qxfHW8brODCXBJVOL1B63haimEiBXJRwEzoiO3xqT2BwPKdl316X
Hr43YrKa+Go/EfUX1k77Mi40IBwnGXpfeLYWKZMp4Cikc+mx+pf+DAT5ccYCjCCOPVuLbE8D8C96
mgXq4vBSo2KZ5LAyl+a1tgsc6FOeqACeYTWCr+Q1m5hM1/c8dy2cNH9jWSfJn5/19CuquMg1Rp5j
g+UFJNOIO9fZtSxlGGQNXYe1fHgCZSHq4gh9Hp95lej28t2EUDBuOga6Igr/J1+R88zE1F9h7tP5
KCklWXrJJhj74s1ONUWZxECpyAF8MlSgslVaT0otzsSEGDTZ2UePVxWhkweggmygXE1q1uHO6b5M
dKFYpX2Ah71wkXQhKO2nxzLVAcM/4Ij0pdP1cwS5rAjutDhHCpCtqTaotKbZeS1/e1G2/ZsxE0W2
sKIXsaGerxytJnrzaS//qJBSc18hJz6NMBEQuKecMR0c7Dh25x7Xpz5b+hWOk8fsgXX6mi1wtVAJ
PsTqnkyMzpEQ5OpWw5C607ylMjcR1ppbOSIqVUW8cQ0EpY37HXZXPYt/t+jnx9FLQvMeVyDnwLHi
48Ci014c4YkFfuzjCGYue9eIlz0st/qAv9Ka423gtLWoo+bf9PR4n2gheYiOU7bbzhvWQaEM8Wmi
3utZG95n8UYuRFi4pYrvWcWOQWC845TDmr2LZsqrLyhGoQKRoEnAxAoLVYfofV1dr/uUfLOPxgyB
c42+ZMZvnnj6egyK/oJ+besvxgDNE41bn9NL/eT8MVXOh0/yP5NLeLWnC3VgxoMy00hpe9Kdc7x2
JDFslQpIfeYA00Vhr0s/Ky6aL7PlmjTZ1SXCVXHjKC/bLXxrSpTpcYWfUiHAslF/xYXnQb3Bdn1s
IMmCgEcoo795oSDLyH0IX1+NG5IIoiLgMabGGrtPPq6XybbbGiBljsUjj5/T0Ks89cQiTwzs0XLY
EPfjKiG0WRFuKCciXEaQ1ECx9uwOAWkSU+j0etH1xzTL3Jw4qFIM+IV3OrW6PYuNQcihybaAtGvr
3m6GkZMPmvi5VQqYz3V5ZoWnPxsPb7bOWNHsN7kpKsU4FVSRE/bs0unphgF3HjWGlfJlm446xasB
VwrnAUei/6kmjyoTlp6jClStXqjxLhtTNXUXWO21ChD9Du9EaJp4UFg4prEOL/drfnHmcoPSP82I
kLZQzfgqyFA8pbupJS+fbGlbvHs7KITfQUjpBegvfCWRWZPatEPBH2HF7fzZMR/+19QmfS815yqf
qOL2p0s5hwOP7juxQ3faPOJE8fSnfegtxI9TVzFY8ZQFNK3uJCHhNsCk7M9bBLkUtHPGR6mzBkSd
J8J5HLN5odGoQ1D3p72RwKRomnA1EN7kjZsZcl62uKnQ2mwwOOy/MEJP9PbONs5sq+GXVdC6wtlQ
6XV6smp22QO4iKPPfUmpaPjnjsW5EMuGkDrY8lVSDOGhT7Q6dPgHOdurynDAq4Yx2VqH5Gh3RtL6
5VWeqMzeb703I3HvpnzlBKr+/yzv1Ybn1eRypS9iurfFGB+mM5dHMWAnUUZfa3YH4dRDfilQgbkC
0kokbfGuRSWbnk/5e5OuUtyQqN8gXTTCtde952uqu9oaIhtLW75SRe2Md/zq6AwRgTKNOdF+VJPG
KgSv3XVCDmfL/X3FYon/9L+qihZozt/xHDbVIp4hYdXz15QdVOVDJyw8ug+lbwkWuy/GiT+HbXrv
ndI/IexK4RoHEuBhsv2lwZWc+tVPnG4BHmAj8jj6iBvQODD7SwoPQikYN0BTQJMAfWTVg5kJglqu
94EBJpU3dPe3tGJEv9AHSVUg0SAGX/8szjAY0jVkjcgS7ZAsf4V2SaGQs6i6cYELH0g2MQFI6YkA
7HGxKvY6oaGp3Lg0tPcvWFnEZpk/gJq20JetS2pmgcjV92ZkSFX5ZfzSlX0qLDH3INIZOJYCrKCl
LEbddAMXItaHe+Cx+VlwfHJk+DjP6ASgR8210oE+HtXT1lERYULGASSWjlxSnpYrVkrFW1Ji1Gvh
TwTmkdhpmsgNxJT5ElN5Myez7zFZ47eiMKMA+07gwRooNBOtzeHpgb01n7vFZqJttpytuBKYIYUr
9A0X8NohtW94e4Xc87Rdit4Gr2pkPB2iEDGSqQXj/JR5eTN8TWtwlf0JfSVMcF+ltGFj7B5W8dT0
OJPM6TtesxVBmojpMV9Rr0/i7QsmgUQGlyh4PJZE2eGQVn23tsGg8kvJjKoGC4yAPNRn7QNgwMma
MKmi2+3NqLQnPQJSnCPGkLujQZlmWDrghR2faMhVO9egat+zmXSKeI8UGqRaSs9OdtblxEC7G5Cc
nBi5NG3BAmZvvuVDtKacoHJJsiySbsbiqbFrVhz/+JPJZLsmPg+D36K/qxJy+rnHHbssuSfkUSU+
ZkSc9xwnwlcuVdWSFfF8L+Cb/QastoewoQjuldvWW2/5bL4SHhLkCHQcVvOUVRvWgS7N3RjGrNQH
WTLjTdWSpJdkeA0GHSHxl4j5yIHMk5q7QrttMAMtl6qWmR39hJcUFXok/POAn08uUR6FBrXUFq7y
JL4gXdgdhnLUVEjinlZ2PcB1+J6hsZJ4K/3rtsEWuFaez5CrpR+nw+UojZnGs+BZi732zX7OzZXy
4McAqjRgQ/Bjb7u8V7i4+XFP3RWt5fXqupQtezqwnNB8ljQFaqbhCsgWZuTAZ1nV4Hp0cLFhqp0N
oShTQHjC3oqGyTjEzpmoG6xnM0UYsuB0G6JkDdNE48TaqRGipVqM36LSEK4StS7O+mrH1WZJftyB
0VUD2h6qv4QpF1Kza5Ub7fA/8nPIWgzK+D4CW+dYuk4xkbO3xd7mYUjiNYKn/bfrB0RINIgMKlwm
EtYYGBHV4WcOrXaxxIapcx5LjONEu8hf4OPsOB/7qfFfrNl8xR43e3uftJbaNwwv5x6B6f51f88T
4BuBHWY9/sx6tE05XN49Wg8hIdUPCm6K5PMBN+bZxiwvpgURE/RKpoaeg1Ef3cWnlqgJ7LNQ8cEC
G4Tn8olLq/g85awSlUfA7S35RzEwit7Tjq2md4qjZMWkSvRn4tam6F2U7N8jV2hfE9QT7nWJ5ubK
RljCEbtoqedT9VaLuz60siuOhU4ddruCtNiR2EwWQrfCYQ+glkEhbBLqeynhrQI9BGRVtQdHIquc
vGYwjrJUQj1AgudRkLU/8lhlQOiPkFX22m+y1rZjHATNPhFWA/+m2jyh83kSEZm1JJR3Bi8oDYai
pw7qYmtuiH+6kaG6PBtzGxR9w+hZjI61P4kMSAES76n7bGnGI+9fQPHm52WI1EgsmD/pA1pAA0sI
FAQp8lASI9UOmG6G3Ssr14xjpbS0Q0Lok6uHcZs8OxolLjJHowxZ0QG9ZTXiDqdcvAqprAyTgGxm
LlTdlIWd7zQl4Wca6vgUAnX3CNKWvMnRjX8nbxI2X5STxUgrn2RmAgkfHGwBlQtn2N+V/ytPl5mf
frkzsuoYwXwtT2e8Y22GSLNjZERrjK28HYK/l/UmwB/W4eGFTJ0QVQ5DxDDCO+YVyPhcJCQ+IYrk
FSvJu2WPJjM7a+kTf/GzoPgdlRwajgSfNC3U5gEyPrvjhcyH+f5i7F5qQP7hBR7uULr9AGxrSyzH
sfu//fqT+p87QG61qSyaqfm5g9Tl6M0fPtcUHWgzQ8Ueo9JK/vw2DRD5EbYTzcqcXWAD7E/36bjr
aXoN/Pt8MFAcLFfHaZWqfAzSAy3QvVmo+2XL+qKYsl1w6WuRRNXvJwpEoh3Eko/kdpuA2o49e7s1
h5fwPJjqqGHkhvVJ9+HrqFZoJG5D95jIE3NqPgHqyunioJpr0BVlfvZA5Qgirq+thv6w566z58X1
uzvNTBmqyVidmqrBlWgpvTgk/4n3FjmtmJLB8csByWoGlw3CqJlNo5fc3K7AGQMtMJsodG4rAXYg
xYh0FfR6XWf8lbh7rfgDZIXltbFdnseGRNSb8NbQqvos49xMCzOlSmQRreJj/sPSmRy1mA2u4gCS
eE4bBu6nakrPIpM71UEMj31ZMykxqzOKHJ+2FWI3dGEOtFLrEeG37cven5EHvJ8ewWA5AQo2IT+e
s3chYfxpCTkGFlb/6s+5ayPQ6vQgXcqP5E0A99ejMZlOmzk2MHGmJI63mwOEC2VFnQGzA8LqX6qJ
AJ892VhvgFZSh0JXf6Sqz3OOASWvgAivapQYdXilKum4pAEgnONJ0hx1xG2fbnS+z0MZ4Kak+xv7
OjZiLaSuxBkmP6z17WnXNMWIenZtf4BRPVCnJuA/jVzNqTktt+C4DkzVAbGSnx+94gEVAk/pxDe/
FHWnJQgOQOx6QDE2dSj/WfYZuQvXp/fpMuBLixigHnproAGlHZGZxFpUL9jz6mEPAexK7eSseyzC
FiMvr7zdJMmmV6DL0mNzfLJcI0Ggl6rv0txoiHrfC9g1MKRG2f0/UlsQN/rieedCnSn3802y7Bs/
/n3dXcIG83DJalj+V0VaGPYlYrNiNVTAmW4q3vgLkT6lNIeG3MPnyjhsw0eIdgEVeNbQw90aYlI1
odL9DATPyqqoiQQnH0xcME9sCvhUhC4rpbLbDXM3BWVXqZw8hqvO+jRtZbYUEpPQbBfIPExvOdRK
+IJvi50cYLQyvVMR+UHN+aW+bWG5OBL92raRjAcl936Tellq92CVLFFTFq1QDtJCgpGZ/ZDJRFlO
PKTbFq1NDvWfEfy6HSSzhhaTOT9jROvTumm+uEweAM7V4z0RDlXoV2V2QgWA83NBZEHOfmetkFFC
pZV5iFb4RdnWVefJSHyOqyeFuaRk6r0/D6SosxpXv2fM+ul7QA4Hg5c4mS9KiWUnV/Vg9/OCFSUB
9+W3qdjMRKYWGytJ4zErK8ZQSTo7PRGkzhEVnJh6xuP8ceCO7d1AtKwQJGVzur4NTgSiD1DRDozG
sW0qgdZiDX0JMMvoUhvW3tOmmd152wYIwnmt+B50SfXbRYv3xvYFhk4/qwk+AzFQnPC+hajQDx/z
qTo0aFsH1RU5ZureZQVAukzXYVy3NE5I9oayW1nBWEj1Bvb9bdzLlmslABAsF+yr/wpd8EznUh7h
Xk5w2lCGqyCX9tV0YcGJ2P4DbTyCwJzKoVGjvM1mTg0NJ4NmUR/ANuQo+6QoDvwYVJ69xUJa4jah
Y+g/VJ2TnH4fj1mdkUJVJGMlq496NhhMwSrGtRofD6Z1AKAyClxqQtw2MFsPrsRKvx1J7m24PFvg
Wx+HAVQ/Xmmno2X3ygDd/YJz44k+UhOIem1XTpNzTU9GZOvDNaYxU2ILpPxJrV5qXLwaZo3nOqn3
lgKKSLPNq2XF8gkSXBqyYVl+PWLS3YvKp8e2QzuKRXQuchba4Hr8rzquO06xVlcPBjxsgqzCca2f
FapE0surnabaOtCoZCsTFDp+7ZMm4EBA6Tyv5arH+Z1Pc69jKvyRItd89ansoxe2Cgg/iBVcDEEo
Px9OQb+gknY2C6n6wOpBCxR3LGrZgNHzuhOinwRft6fPnee0L2IgrK+iYrVzipm8YHotFrKplSE0
fPdDpDqaWpRLa3PDw9RGvtYSl1mu0v5fhC8pMyk1wN4Jv4WjxQU40f30E9JzCOxGpIhzuO/cu2o7
BkxUOcUeMxx5UelA8lVmj3gXkHEI+p/z4VowHaIpE067YPPYxLD/kr2Svnndp1kht5lU+Z4Rs3Yn
T3cD3tHkf8l3/MNBChR3J1xAKMdVP5v1YLpeqDyNlilUjm0oTiA+PoXeGD+RIcBxD+NqzWqS/Cf5
p+MkHkXdGIHIJ/CaCeDT1Xotd7AC+ztMc6ikVGG5Coe5xn/799uDTKqb7iwpW7Z+bF3nWirqQp9f
UWJNdQOimgIi46M+fj2SFR3y7qtbiziufDto3ZV8EaqdxZ1KR0hO6tmlOHAedDVjMxMjNdFssrrD
3vWZQ4f1/RIoAhze9zBA+hJly+Vv6bxPCdz3R+HNnlM1gH62GfBPMNrXYpkYWfOEIg8ztjIaIPsM
xxc4Pi9yr32p623puLtaG+IXaBy5HPXT1DtRzIOQpxcAF8JgOiYZAJl5jq1B0tXEYgLIXnYfE8I8
CLvXFzXmGNZMBGMwNYdqjmoN4Fqxgp99CjY3hJ8w87W5EJQjwmluhMqynbHq0ElSJRqzt329bEHn
pfcxMv4t0s7kO1QvWcy9S+Ts3O9MLti3oZ/SFMtQvldXNsAmr7dQ498lr7wbvFIY4lb5Lhg/ZZcT
nMZbx8yjzKVMo6YQsMvLfik+khUffVxRjsv8sa8+SbnlQWmmfWTS/y0n5pZ5xgGik8NfzetqqG+E
Mdr/xKxiha5Wm2KVhN9epGJ5lbYF2YYXadSNgSa5D+2P9gePH8UHChE7YKtrBO5X+wyQ4Njzs5uT
J1ISB7bScv70g/EnRwRCQZKzCYgb8EF/Ix9BY6kULZnBZRORoCzdpFwyCCS96ydyUA/uxfBDFSZJ
kjsgEEvmvF3IDvDxlrXvKWUtBBP8spUZhG4OPESYX3qbsh4MjU3DsgVQRGCw36ITq6TLTlWLUbQ/
VP/Hm0GjNn4RadQdwzb7tAe/lH2F1FLnDbCGF86wKWdOuLDDN4VHvKTZmgUpAIRGFRwBCI2hAIq2
rmvNWgY/53iBQJBtMOsyOXnGQj1HDzBC1SIt6a5Hd9AsDXwFzuR3YzfXfla7IQnopMZDPhmrMDBh
ns4623rT533Muq5csM2gvLWZFidUQCYSkBtN+FqSLqxK5M8Wud0SikvbGQNkSoqdujCPucYEOm2n
WeVkSJpjfjWErxn9F/MfMqD6VJuv5dag0mWlIsNIU/7iLEkzoIZ4vx9+wHtaRHEKOC2lhfNBslTk
onRBv9kpCgTRICvLBizYHQ1yRhz8Y5scFP8dV3ZFR0wdJgvOGOqeLXQ2nh493sztaW07wBqHCLrv
A+3GhDJex7uf9yntWpZg8Z0yVoMnHRP9rFC5bGqGjBb2lk4sVZBu2ezRh6zqYrqu4/v/dTEKYmGu
71KKoueIql/59NCdE4h4QU9gBKNilV3bkydImuAlfT0G4RxxRkJwh1YKJS3Lnxt2XtKfdgg2t1c1
taAzUfXcNeLY+JgZwYbqx1ahwrMQwhvTq71+tsCQAKlLH8h0eYdXHWl9oYn2TIcxB8K0r7qWafAc
79vWdp6JjA+HWm6UDrPSM8WnpG15rKmRbCaFNPCNySrJRdjiYX+d7OY78TRIJnq/YmZn+iRxr9M5
KbXGZBM61Yyc5TOUMzsMEoE961p7adk28d0Pednu39PYrJe2UUpnQTVxZgMyTrA7g7airMyp2o8p
xNRnoaebazfoVSb6NJtqDtmEMykrpFg9HxekkYFOeZMi9QG7awQRsvkxV3Etcywhp7PzzKeQyeMW
oiuCfQWan5NA/CRdSVYt8NuyJrpFGytWxihF1BjVKf4slvIVEUTeX+GkV9vWfHf3mprNXNgKNPWN
u+rIvUiSXHXYoUx6b0QkNCJk0vca0fQYHuyOYuNcBsPrQ60m+tAbpN9E2E+RJCfrdM3gTu7gpwi7
9OwBPhTYNQSZV0RN6sPJjUacGUVK3fw/bfDVuzMoDJ8sG44jE03S0f6NQA1sVNRRe/g/vcgTSiXz
XV3KeyLXPTvxV4W4R0ggieREzuG+zrShYTlUpi2yi+8z7tDYqYOCdzws63VfjtZ2Y9ZOmqGCTVnc
4tsGbEmgWjM+03EV8CSBfDDJWlVAIVlMNsoB/GxqDNgsrwA5yNUtbr21uA6R+vAZMZbtsa24J32k
S94Ns2CnXnAy+6Pmg5v0B3T704gdyJTUlQzuQpNyyvIH7p3DsUJBkHVr0CpJ2tX/ox8hNNSJnMmh
vKgnPMvx+PurhDI1Bu1/bWTP9lqDrbBZR/GQy0goMn+kgKerJGh9sW9GJj74/qD+UmoPYrahmCYg
Y/UveKt+EHTT899jgPqI8Ja1RdQC0WRPtlaj1mV6P6beAdAVA6Rt3psd9OCWp+e/hD6PEqy+tA4M
jDwEKZtyVP4RJayEOKAXovsvwrp93Nx2huWl1wD0+I5/Qbfl0xv7bNgoAXQXvy6V04MKpIqEHfgM
Gg5hHFFxj7ggg5/ABWy99diI/rcAXN6O+CJw/f7J1WyMsKk4/ngnJrfL647xFoB2rFoqNmNdIXta
ta87B/hfm/kgD32jlXL5C3u9rFCH6mKSMrGIawGhTi0oF0/4TdFSLLZEFmoTPZDJ+rVVaFCIsJok
2LcYTgE1gwCcvGHspoCvWETtmirk1eCak00QdP/fkHfiR7OFefR9yWnktW+xOM28YwHRG5DnlA1g
ODUHOWuIpjoiZOhaE8aeXFk8XIvkZe4u2T20daIp2nquCktMsvHEWXxOtRVlrhfhRQae6DVw+xXe
LDCJGRr15oiltcwkyq3yQOhmYzShTjPfBJWiSJ2OLQO852Vd4AVOklBMUbqpAuXBql4wTraudxG/
6Woxb6la/BmYLT7HmyZyTiWRCNjFnnQ1ufuBL9VWhQZOLFmgfC2TDMJuW76C4tTWNUJbmqBvWak8
lcQNsWl77PxPxXiFBSpSS7IvVQlKDRq/4epovBwWp7QOw/r806EXJ8rr5jfIF6cy0y6X634hjemb
7gOge59kmuCVXTNFCCefREbA+Mv9gJAZjpTYMz/NFZEMFGxl6wa7atLLf1z0H05OXRfsqybNaTUO
xC2wtLxjkgHvW/CTnNJrJ5mAA4ZElFCftnD502jYDnsoO5bPO03GBr+zyIdYbBd2cVts5+vIZbKS
S5fPg2cKvFoJ6AkfTTTBOC6myZihBokJRAQUcxOTi2WVW9g99o9sOqpeHhVwyLIZjVo0cG0O7LG/
pNELKZsgQvdEfL9oJ3zzPD6boV9dtS0QSSIRhkNVW9L6QagzUtvajoyWzYehNm1F7hbzy/s767Q7
KeXi4cUm7If3POuMNcYrMvsaePZMyLUNId77H4C/rmtvzunQ+CMRz2QFgUBe5XVP1l79B8mQAD0z
pmtGvM5wJaMgI35govAK+N/Tz+CnhizWbBDXEBJuW9wS7kwdT1qVY/bjcsQ51+ZThygJiCSv8rRv
IhLzw94IrZeZbYU1pLR2P09akZwQOoZV2CulJCykVw09VN7CiILF2W0GJ9c+pTRFWWK91AF2K+eb
1Y7F5ODKTTbSjXH4vEyvvzDSOzLPXEn3hNRXoF5DSNJ8lH2VQ5PIcJUWSshs2eTvhp+3w/PmXqBF
u8OogM8ebk4S8pBpmgDlB5/W/QoIV0uy0FcL5DHiJ+nbmwi+PR4QeL74lQVyFf2ExV1PV9d6pgAB
JPtOOh1ITBRhUyGVZY6Af2nViMxnP7XG8k2IwrlPpdexPK0nOVVByGnH9Zla6euQlCwDK3/HTH+k
DdYj/J9riE00YNW2ugJcVUUfK3z8nSLBcYtygCcUqmo12xqKIV8ghmhfBJfbizMjqDw7Ve/JFoJ+
+8dgTQRzl33JU/s1bGDk7qS+BiSNTRPzw8Xi1q2HozT+5w4V/pbzg3XxlVrhNsnIHl8A9sIozEyk
7i/5xS0cnb6b3A6MkzPC7l9Ka+vdA8EtwdNX6k++J3UFrt0UA9XN0z52HwEdPSCkwPcXNcdHyIub
0A+TJ97UZuHkEmpAgoh/yIfedgDn9bSdAV5REVItR46tcuSwEANF8XCzuPWS/GumJwe+MTujAZ0r
Ix9h3LpgDK/abycGTI3eTctEBAT+NQCZRkvWkxZcd0yzeOgnXFP1ljw36y509XZBLFNkJhMo5ypK
wvOgO2x5jCta1b1oK+aa7gHsFipD+r/S8K1WC0EAZSEhT0DT7Tn6cBmQiNDXmgf2VIUXJutj3SK3
kyEtkW1dPT2pgmSwHiCIMNKV4a7LzUssDxD8IZYLOI3biBDB+grn3RBbIIP1p5XRsy833gvQmsKl
PcnG3ZVNbg8l2gxvnIPw9Y5yT2u613X3opicHi/cvGMnsHxs/wK2a7YBbrgpo8lnVWpysNb1PNsL
/tTPWbLIgfJkImL0EdAxpLpPZv7H3Na3ypf0rBuoGMP/TjLrGWsQQHhc5DY6n+PL/C4AkJAdT7UK
lCpmHQ4oiUxu7WsD7nJtsJwVikSpfK0lsU7Zj4CDFojefOISl9euv++DwdJ/INsjO496yaGyt1g+
fbAMJBnZRGjV7tH/22W0ihrHmrlOnUljo/xZ/AFSTV5S0BKX7GwkRCuVaZiO7ecpn3OB0jJHDX5f
1+4HjC6JyHR/I61T2V+pgXnezPyZX/QCZ6HdhFRo/MyyEKtDy/GwiGq9GrNUnWM/UPfcB71uMAXt
NjE+X1P/DSPv6zhjsVhDeGWgA0g4E/aLLL1G/XQk4m1jPY5gNoW5b3XJW0MuTmEgKkU1aLMCDKFZ
pk8z7A4cCrOpUi6gL/n03kwi4pLzUmSaPy016vlPdq/T0CZvXvDEsYgEDGOWWGgjpKj4P4b7RFD6
Dx6XP3k+GlRdcdZeeZIbmlm6cs8RjV//P+Q2EUdwm9bleE87LhbYdaEp3dy1V9pVQSyRG0QxtNQ1
j3t06j2eJ3IxaHJqF4GdvjTb1uilH7LxPUB4r8F3ZuIZDRBp2E4fRLKPM/CY26DxYHKDhKtwHzc9
HPkDR3oHRcPQ93m5a+7rlhMBpMQSF+IOvE5e7Zv2VXcydxqwrFg/Hnm9YvFj3BKVUDDt9UEfUy7D
UB8gnEWJ4V0E15O1wcbfXc2M9GJIJz5zQX2LqxfzTIaN+0Mt4UGGCeHq17WXnHS0eIa7Q9FCgSMh
ckRZ1j3CHbnZhmXxYMyuo+V9z/flz16+Kw+uIqu6BxtN5PGXGzZzN8FaP032U1wRr5Hj8tabCzGx
0ornQ5hnWfIsn665IIcahMTUWSFWiKDthZUmKYeCVSG8CYRVvsSuyk0FD/3ydGAD8SaoapSZdsdt
pc6+DzWxLeQhsoNgYo1wrTqwqTJ/IkHj8DB5QaS/Z/Zx1VxpyaEoBEwkGcj6NzbW8/5ckbv+D7lH
DHR12xCpvtljCi+jzqCJls6XQIgvfriUr3CxRoLyN3+KIhTvVaBw8M+jSZvsSQAu2/DR3XlyUMwo
zKKMDOTeRg2zn2uqRe8/jGOiZ8ekEnPcZYaXkIFq5r438m1g8Au3205Ly8oxV5aMYKLB4kUoCkc+
H5hCEtD3H0pljNPwsSJ1hyxCdtZWXjxnSapvcmKjaQIaZZR8w8KwsCNhQbCkDxIoUhM6554C6f87
rTVqWi/SH0r2W57tO6BWOvsH+QIu1yj8SOt1BeWkfnnjiMx93b3DT4MDmC+XiolZOTonodp7tH1G
8R/SEGPLrsZP/s9SJQp421NSNg/G3vOpvqQ0RnB+OmeiAPjpkDZcWg8/GTrI+wSU+RXqTQdQp0E6
pwfLPGoLpK3aNGQfCx1uscMqExjOwwhgg54SNsu8Y/bRkzSx1v57mp1W52qM3aqLh42ODSPf5xiP
TdGu7eTfvJly27NvcE3ICHlXd+n+N5T1dzDWzFMW+uvM8BYr0eyMCSQ7Wz4hrNU0/3yHoJJZ+TT9
uBXgPrykVzTA2G8zjE0ZFR0Ds9XSK1MvciKA75SLAf+mBemH/ikWka40679oXrWhOAVZytf9wdV9
j7LUg+8TirGQTO/aEHekNEOgENJoFYY/l430QnT7bjyTGSYrMIaAUo9cs1R2CaOp2eVvUSad2vee
VEK+fs4FwMwwh2/GttTFnmpIvwZ5jORRJp/hfoRSJ5Y4DfB7Kecukw4YpsCDT/hSL8xXkVIemnNZ
HH/jyRP7SZV4YaBF+Q1FCkInUR7fuZROCd0Mtc41fKTEWrWO1JhQownUxzEQcldn5AtgRBHhxTmc
jb1+DiRHtRbrdnT12l3UMjTc6K61RnNutHmpIRF/IcJowuMatyVK9n8VEKW0lPcHlCnSN9kV7X6b
gX7IzhM6q8rHG7Nqk8dRAge5sfCsWuO/poQTiI9TAwjnu3lnZmpqouXnr1jIOJ/Qg8I094w4Wl8F
tLnuQB+OrP9zOKSYdj5gUux95hw1AenUTOyQ/4cIrTf49ig/XmXwfvZSjBvg7bpoODUJlz8VhWF7
Oargx0y+oVsBmXIGdJcfsXT8TVXgraNfKbZ+h7kPQL41mC2Hq5P8S1EjKkkkK3ScM8fdEgXoDOzC
j251WnU1PvmDkSEfNCZ15EvfZ5np502b5BUYhAAPRbhxriuGcLPQuzZ2iqwR6r8UOmIBqRPbe7jZ
y2LJ3QLg9aLV+h3konQOI0cm/+aaBzdufyjLZurvibqlbeSDPyVBMWyPATVj4YVIUuBtZzFOelCA
Re9U7Ul8qjxPjM8JbURbGNF6EsfzRvK7XS7+GSKwlffbJE/m9qplHWZF7IF/f4Rv27Ha8l7ymdha
SZ8CZ0c9EMOt2WqHP+2JUnhRYbRmbLR2aDqST89pToaqBNhHAE92JHDwifPWptdeJOGjzjFf2/B2
ICO/qdVGkih5NuTsq+HHGqv7fq8U4U8+kl7f7UwmgdgTaJMeY/zhrzqRChK14Re9ZU9hDZLCFYjL
FS2/1ymKLZZbeSUkqPrXrZMj2VirmY5CFaVYuEPlqfYuO5oW93htLe3SpAYeV4ilC0Dx6g1rfGsK
1D3uf88oVovFL47GR87tz1VGH7SGBVYk1X808w1gmQYMpZ5VkHTfr8Qs92x2QrZHfFzqJy6ogqOH
hhNqS1EJS83z4lb1QIvLDqYIePAjBkiJ9WhPU9ZPZmzyO34pnL8lHfVoXkuuHVgjzCoYMNVFVwJl
Lb8BkvykA3Bc4xy/i2qRKqoZRotMAYWgl7uWDP9vNbpwJAcBD2efNp3FXUTUAc0ZSz4BP678osnd
FhEnDuLp5BMZiwwzKR177oA6FgSN0K7PFXPwAytKmYjdJ8GLsErD2K+Xiv0kYhnn1MfRIQMpsl4a
DJsV0ucG5mu7OvtN7gi3AIuOLjWiOqU5yX4k/WWS3E51jSpNDuoKozv1KlDjMmZcMZvUEtLxAK52
NXvOKVWHe5XyurOvPrDQpQWFJn1Nh7OSGjHbXK7egud6+EMllMovuQz7JdKhAhM6ryBRSHvBvVWO
+h3EHbGGblymiZMOlRatdjaYLi2+Mf7OeNvYpaLPY3korDvRqHSeMWgWBQoQiFDWQ2vWt05hAKGR
X0OrmQtgreOeDFPXRdzPalVfZbiJ2m/OUb0GaFYUgkpk2gwQh9EQjd3A93C4YR3iOl/Ttv1jfNhG
ON04WK/r8bSHOip1r5JCjIZ+y0Yb00Sm0+K65Je3TbHOqTwInX2XG+1M5UlPHmWNQ3Miy2JQ4D3Y
KDvlE7b0vbIGQX5S4fRX9XtT0l7vXHLaxVFCqTZpr5mMFFyaiQaw1DtiJCvEVQdF2x21tZiUbSRX
CgYMZrJ5nvDub67PGGtwQA/MtQ+F1IyngfElhdgfLEkk0NBm7uDz1zkix5Kajjyc83puYp6d7cuD
Iwn+n3ShOiy7XZX2gqAMPJMjIq9SZz7kTwWw0SMaF037L5nl2yVkHRLvN/UY/GCtMq5B/jqg1Zs6
DRMCmcXNit0tg1pikD7BPyE5ieaaTUNU5aB1FAtNlYFZLqqeb22YqgKppy9FXhHO9MsDFaql5oIO
qTN/yL3olF6ODnMDAaxujHifNqxiAd57KSyCAm3avjPkHmkRuUY1G3IGOLz4WnGf8ihWepuvU5SD
NlUx6pnpIoNv/JiS80b4s1f9hBJXG7eJtYgQFcNnKdkjcnBDhIM6Y7g4wonUkQiVD9GnCu+ZcMut
4kh1E1Bckk2OcEcKSXHW8gEfbuKDf+6fEvDV2vygEYfl4EfuEP9IUmb3I9cnrTKe8K0HbzsHVPAG
uDcBvPdUvKvR+i/W/RfN1HWfhRWerUKOWRiuU3pbYgaDCUXn5wBRTmFJ43BtI9tT3EHKVkKjEk7D
rFZRb3SlPtrwOVUFcECLGi7lCH26jpGYrFjvWzByCNLj700sl3Kwxwq7xOL/LPjIPhAeHvoR5/Hh
0+HTe7dW1TYKC9KZd3FHrHHp+mEUuGcFaUETEh/KwWLP5SrPpS0KoGQOjMi5xZUSd1XO4YdRuot0
mSscwNwu6imtleqVXZmtZuimI3q+IX/jg1kmqqeeCSnkvGVjXZGRWjZ741lYbIFU2w6gN+h6LU0K
E6pt7JPvtqJtpt1pTUVT5yCBOrZY92feYtkHUSkjYM0lRNWFgvhlIfM7waAgCYQX0ZOE6fLHKDIb
PJ2HwGW9GE641HOXbG7+vpE59L6ENprctjuEvhLd4TojXjdDpzdr+Ho3SQOFFoF7gUt67AaILZHi
g2j3TlkAqnDvfUwZVHgABHPpGZEjPlqqfJ06XeqOQBLQmfQEJ53iWINNi9xQ9JRTe1HftJpQ4dov
PbFKsIzFDBg48PIXdOEzkL7P3uZLnCpk9x4Z/BKa8bcOaBjkO4nUDKzmnESBwaZaxHJ7nal2+K1h
+EmHahH16GR1uibVtc6YdrONq4PwA4wd9SA2cUkRcAy6ixZ1p+68fSnjAFjFWpD7zl08uE4Ya5Rp
aBpgwxEKY4LZK5t0EIIJUUawS5rE/mRy9IyhSRfYyIHSAMLN8r/SJzrYrdo5HQHj5Tlx6u+tVUaj
QS2QO9xwAr/IEjZoVFpqbtLFXxsChU7ty1zWuNGBGRoIu2hJcJ/xBoenBA7xlaXPxfo4BBbYLK+o
VZYM1bZDEicuLazDndEw/eWBLtjPKEJl+H4SN30PJIZFVnf+HnvZMhWMgPu6LkiidkdfnMmHNW3R
mJl7dg+iRl3WnRs2OAVw7dL6DE75qWbmnrGmFyXr0OffLZQ9BC+ae/k3Bpiy3ejIvvbZYvv/xDYG
+p6VWXgyW+j4Qd8PGNosITN6JGjDLoE8H6fXEM0iO/3KL9wxny6Co8K14/ZZqyIZcHEwQA80k/WC
/G+R8ODOxu3Vg/ZKUuBq0gKbvLGatSBpyN6wwrR8ZRcNyOJRv4W0tog4MpGHg5g5GkWP2yfjubHx
nRXixxLNzcaar+W3VVXSYzTZb1SyvLp4zEx3oJ+4qX3NRxniZWlMidTkyJ1u+/Jl02e0KQ/94HM5
0fbX/BR3tS2a0oMDhOAHE23jHrrfo3yqRA92TRngk3PS+wA2BejAJrkyf9Gifzik+OA7g6tebul7
JJakbkDK85KpqYrpQ7MMdT+v4sV8lhsiQRKjBYIOfrf+0JZq8q2xlVR+nRGGvG1spLaH1s2D2yve
ds3+a+B+2ZtAR+Ibrb615MWOL9P5PuCZwWSI45ECKOGuW/xCnWpbHVK0lWWv2MvAXD6Z4bLgN+Hs
nU/jvW7vJMgaqh/DS0nfcOr32wa2+TPvnY6KsDyHTYuXL+DudE7+BqMJxpLSJeo2nATg7cDrzvqn
xPssf9/HFAfofK8KDdhoSS3xGoDZlK812syiE/GPWHp2/F1TByq1LvTZ9lRSc7HDL3Xvb417caOq
+Jfd4fKmD+zmaDFVPdKkSBuFiDrr3ZHZPmPPbIKJfE9gyo/gthnMNrzRR8F2xfxbZ76gFh3+L+KG
G4sSA+RsOUs7qfEPFcwU6XLNtCMrB5pzmpBxrYFaj4oDyIyKBeVaoV7O5+aXoWUYLZtZkcGRy2QD
WKDsIu4HB74nhAM5+hnSy7C6A8a7FNmlcQ9brHAQwc4RBX/4UeDBJT8eNRHTQ+BaM2qixFNennr7
MXpgPry16mKSfybT5lKCV7oTbzXoU1aQ5c6S/uDI8jla40itmPv4mH+oJiZucoMMpmXqSRTI1Rtv
zg6sMhpdf00Frl+qANhr5YcMIWGQ4RRCMwJR6l9ikH4jlRMEUmxMdp85GGPXh5L0ZQf/7NxqEG7h
rWTcL/M8plrFZCTAVPRDq8yd6wEvmqusv0OjehOHcx9XBYZWGiOLivDeTCyMJUQ/VLHXWoyx/kf7
tuW6Vq9N+s3QTeA9qOrIFyeLs9bOmQYk073W3bjY7z2i5MHmZ57XwBWCGH8RnLWIFzYRM1nb6YPl
X7SJotOtT+4RKYl0u0CSWIIaCvVWlw/jAIZz4ezY3HD4zj2CLAGtcduMeAK/ldCK8IpmcwcxWAZE
5xXGH4lGngwzkb3AilFj37qEDzuPAOTHJGo0OkykeXThdnvAj3pHkSOzNQuQXV7i2AR9Ypkzy0RZ
v4H9wD/saSZjYeuug95iz1e8hMs+OHIPzKRz7D8D4JQ30ypGIioIF76O4tBtGUFlg8/TwqGBd3FP
n3gbfJc5NK3p++33qFL2INAOeSCSJbdkZ2u99l+9E5SZzY+Y0eXr6ZTz3fxRl5Rw4+f3Brvxvnbd
QDgJY8Eo8Dw85HUOt6h7XabySqYnP0wH8KbBM6thFgJ57U34GOEqKXKYkfMpIIcm16o/nEVBXm0a
S+yQZvAzZrP59TIFKY6Sszyr/3+kMfRh/WJz2VU5wUbbsbu/2WYUYT9MehvUmuzu6dNDDkkemOfI
i4XYNoGBd52ofrUDRiJyCYycEtYnSVcYSB5DjzGFp26rf2sK5ZDv1SnrXPIR1YdXQSvIila7A3/H
d2DhjBWA95AefCyRs9l5XKvgbORq9TwKsx5CQMKXgieY+aaetCXBo+UzUcXsiav331JFFQUVdLbL
MG8KX4c6AcIFwl02oj2/JOqoBYMhbHBL8Nm3cLSYbjXu88ZsJfNFND5QTveSaDbl0lrIprk/Ufee
PUb2z90vpfZsuFUEHPYM8gtkFoTCdEDNRF28HkIAzAZmDsWLVusvk1x0vAiInRwQQfW/9Wl/CN96
yI41clj4wO3EC4Q5HEyRAA+I1doviQGeXvNnU+r19NFfO+yJbnJBvqbQufp8UB3OBSDNNgfFJr5V
/nkyPVVgSAHpL8Ykn8ZDqA1KEIcIp8vCArGflAg9FQIgqo7+eY/3GXfx4jgS/KpZJo9a/DIy8yc4
x925NopK9SLKoThYb9aYMEOAotdv+yEStPscZKnh3/dF63hbsHEiZUhb9nz3Vb4B5ldvtsD8pHKn
1hUXm2RO2yElmLtrD1a9+vPYEDRK/70TA1dKY9ejSUk3UZ+kO1fiWadU6tYkwLOz/YjMJ6pHOVlp
9X9I+MDDX6DaL+7dPwTcrP2kmJ412mS3ci5EYQRks4dXPMzQ7hWRQ4oTMu/8KseE2A5SwiwLesUA
tJg2LXtXL8Y9LoKLYFbOGAeSugz2Fpjlf012NVQ1XPr7dbEHPFQA8cbvvXMpdaWFkf4445+XOg8f
c8MlvILxaAadvDDNm0YNSd3sPL+I37bYb42LZgDzbTCv8ZyVM1bhjd908wHprrnp6iAZH10alWTd
ew0McjrdlM2BKGhgnlS2fT6G5qLFKPFb7A/AAyiq+jfJY7BRLqELlG7cKU8DN0bVbLqFvSXqGlr+
Jq/lCQbIsvWDFb+/GD3u1tTkmGTJ/Jg7jqZFQnul6lqSZNB8ALYwrNJLjtWbSP/RTj+CaNuQTHjM
2MHUUoNTQKuBcARlrGAV1xBCZ2RXe5W95ofDiBNjXSf7uabYhsF1EiDRLTuU635EwY9EtkjkPdR/
SVBfrXUs90fx2WH/4cTMuGgn/PjWWwxBSABybBV/athn/oW4ddzDIXl5fAUFVK4DpzEvILPtCTQJ
a4V5KWCCZinIm2vFwaKpb8BHR9hYyoilEumK2BCFf3ARiNjFew4eryXmslvQprWZlxYhwqYx/FdC
zQX0BtjceWaJeo9AfoZy6FjpnvOfBVm7D8Jze3t/Rw+EWfAC8EfEUDUtkmqJIkU1DI6jioMvEkgj
dmEJ0CosQNxWvh2qvS6+lPf6moXn+n4EF/RDaMhnZyU2VHNczYZH1uMbdadM6+6lRrd9TM165Jws
8Q1zInzss1fj7zpWHhzEwSRGJDw+IuAfdSli6NZSLBVcI0NhiifW9k4y92xz9Z9PYwh8eDY3A2XN
UZRjtinGrkPGMLq4PklvcaJP20qahGE/U5USEn8AM+q09iUCTwOMCMAaaRHGiR8tWNPXL0jz3BQe
pv3cyBKaJu1C0vPnUkwVHpF2E95ravDJ8zwUF26JWCLm0tqlN3beKujm3EGsMvfyvuw2pI74St2R
UY0+oVOX+Fgi4pHWRwERYwDeUtVSyKGvU5VYP+NiHqhUYsEAcc1SEB+3B4tzM1svfH4GI3feCV7f
mT1S+bN23owWlb0SSAMb+KPMI6Mwa1g0WzHZokLGzQYn7DUaW6SuIcVJMgkUAtiUBp7hrY2INcXh
it/RkyFdjSDLwQRvtqtxdXlFqfxq4fbJzdg2XK+bogsH5FNpeFbTzwDykHG8OoFnvNB8SbvteV1y
+TtOdFvGVw/45sKBLGuTF2zcao/icYqiY36X2ixqq7f55fkJOe0+GMoxERnQX/vLQgPnHw4gCOSh
FYdWIr1dzhBkZSoEf3eQKRiRHsJnjZo6tnh0+QqJ4SdyUNK3WrFf5pSGFP6Vagv4aKO3BD3ntTXI
fwK4pBq2a7NEYWzz+ZSkDS3LGXXviC6B6DbhVOpmvlGfN3zc9NzcibCeJ42NePswpRfccwDG86jb
Zo75ecZluDkO5r6Ht2r0luOQPt0V4XJBMS3B/UEyozc5jAzHYSdc+SaxjSIbkLkZiubRHn95I+Mh
xGGxHFssPa3oDVuKFIX53cgKZO8aFpnUBbZ09ER1zSE5Oz9nKI+icg7roFpcehRq6wI9ecR7t78F
KOsYlHbQC6m5T4RdjccitbDyJO1jEpT2zE2yODWbhLVZJSK76VJlhgWVGYzjL9TKxfP2s+xmvSG8
Qo99GK7JbEbciSf6yTR8wzpd7i4MCnbkW1TiAqTlNiK34mfZKsQIeOGu0SUnqV0v4XS/8gyweTVZ
V46nzIQYHIK1C8+iHYTvTxQh7ULubuHeDIam8s2S/uZ/CUgk8RJ5QyYcWQ8fhMGMiohKwi0kNuj/
t63P0WczrubPFNxmrAu/iJf0R93dnwfjxnvln6dEyWTplfFP84Eg5MHMbnZ5pNfYTBAPyJgRVpt9
LtsR0vgaHQ6zYyFyffatCYguNfd+oiqBY+5J2ifXm1tPh77xgFmZzrowXJIwgUdyGgGuaYgsoPb3
W5EbL0zXSXV/D6jGoVvlsj+2nwSvO0hNsf98g3gD1PNpek4Tagj6jNYM9ptRb/6Nnyb1j4ntz4ZB
6XNkgyLOyMYzcmC/ZIm2VZuog8A4sifj+bNQs8z7Ye3d3wgpw99lONVXlM6ICfXwS3zZj9ph2/02
dQcEB3wWs+uXdxyfuGu9rG8UP6HUu13r25qe3uhlVVk3r73CYPt4X5Uzs+9HIn+7pWNeq+BszdVO
STmYQ9c1gKd3ZcZe7v+wjcs5CC4BAUgOjojLPBqe8W4nS8lumt8LpZYmG8guiZ3csw5uivXyLM5i
bGRzafmY0fUuwYpe2Oy9oVuWcrzrBS6G8p7OK+GoRzjC/mQWfrWS+tZzebyl1JJWJZopXdwDoMR1
gzulLq2lf0fWq+j5P8neEOr1BOR5oTqwB8hzuHkraH/ZRsU4G6x82v/5C3himigDM2f8zZUdBTTf
Y0gSHN4dFrHOzhFoj5HlmWxfGA++FuNw79Iv7Gjp6oq/jCby4253Idsk1jsQvclHsNNbjV/oumME
p6jZuWy3sevAu4+eEZfOZGmaeQUqVm26hDokCKmgjj2teT88vJ4OnodBtU4axiNKsaY5z64gUrjJ
a+s/MbSdbyY2WQHx+3iSQIuAJEs+2QNI091JomtN8DmR6eT+0TGvSWor+B/00TNV7Ku8EgmVNBrl
uPQJ825JxWpWpGtbJjOvdtNwbYgkD/vDH3DTyWcIYvCLmJRodpT79+5Jwp3bS08EqrVgt4wM+l9e
AxaScdjnEWqjrxd2Go6UDgZTVRWE2nJNFKojDsqID7SyurrbvnpcmpwyswQcV8V0RxCcg/mePQfT
LFc5TnClGT4lsUZJS7sz/S7RP0qdUyixCRZay7R0Vz0v8yw94RA5Xy2z09koUeCY+z6tijFKJcWr
ev5urAWfAMRDbDTtfNxlB0MaEMbXQeM1nm7x1wGEmSVnGkWfXFAXVCd1rYhVjq8OFfE4GqtYYVMT
A+pI9iIWYdo9It5zrJRpyl+DZtwI5z9gOsXp69hzx1mXuRTkh/wumPcyOIOpUQ5V19qe1GwRgxmv
yqLLB/tged3SNxpSTexBY/HCHDRMd8176kdl3RrbQb6MYbqwEnVZ9t9xi3wxBTOAu3oGIe0CVUNO
h9qS/UNnE92VqocSn8g4FqHzaSKlM+DrhJ3eUVs0QFqNDNBpFBUMVBvExuTyMO7QOJmfmhlMnp9g
0QiPU6wBSKqH9mHTRFpR48b6GS959Jw8zmr/RD4iqRo9fMAQN7c1iSpYkzv7aJA2+yMJYTX9rdV7
TXIJbXUALvC6U4WcZjB+CbjzBxR1zwEBOnkK2d3SPfedfCQzqzdiiTY4l5tcK8AYSV7vACv8B1dn
DpgcAvjmrwHCNU4PsDFzrTk91ZGStU4qT4C4bMWajcZYqQJALD936B+RhyDZ77+ezrqUYFinALJr
AnH92O0VD4e4RV+ieBePaErsPErV8lxv8EptwVUjgdpwjtnv0Leed0rSi90299/54s63lDG9F0h+
ilKtDMBZY1nxJbxx550hd/+s02Bm3Iq1Bu443ZfUhYJngXyzDxx57sye9au1SCS2giTyZujkdL/9
6pXt2diZDWDvyMHMUj79y4DUZMAq9kl/gLC1sWDX/qt3V5QlS8HCRzP6YWZZxs6ySAPX8duNw+by
hgRmZIaSn1NdwXDj9SXJczgAz0ik/VW8elEWhZstBKGge0MlPMHwHTboxCfqyVf6Kz1s1LzFVFAW
W5WE2vkIx1NnhxTsoFAsd4R0+Hn6DvN9uSECCR8VsjB0JIGF/rd7n4aEOi6elnM4nsj0jg+75OKL
dw3Jfc9KSFCVMEwefRFkRQr5VWRl0JOKI4FeuC4PQUiVDpLEx/ZP2YjUKotreFU2ifKYVobU+vXl
VxfRlpe8o0nHVXDz4fFuu0ms2pyn51E3mP+0v/qYa/7E9KeE7SUo8o8KTBtyEbOtVdwxzLMKSkcF
oe3m7OhiNNBKsRGiihYu5kgA1VoCfrk8mYIS0RKom+KQDDiFyNsuTbfkGj280exLVOxKvQqG7i1z
cMTgmiPoKnyNC9fiLXg3zNeyLF+LXmqris2Lz8FMI0k29xSo9JpC69DMxKy6mO6BugLmY4yN53AU
+n543jsu7oi1zwx3rXAKrJSY/RZ1NW/TVCs43NrmFzkFjckGD3T209uXUu95/AeTMhrF0aUqX8MZ
n6oQ7M5ALFJfcuUC9Be/5lNxfK1t0wHaPuRUVELWcIRq7sdACs4mcQ+j9HtXx97oaiF8t9SkUV0H
b/eBQ51KnX55SN7g+9k7VbELT0747rrRVxG59cwAIiXDCCaHnywjYJQPGfiCGeRfOd4EheBGtSTo
8Z5dfEnooCByOo4fJmeOkWSyZlUYr9g1dnf5Yq1D4+cfgbu39CDTo3zRxG2yZ9bsiinZukuL30cg
hiGaTfFV31OOUvtvEisdol6+AdppUH1NlVYy4QWohIyoFtpiZwOLHJxerAi97GuOnUVmF/1NkyS9
QF6AXA1iiktQ8x5JBd05fPuZdVt9Q+wF2I5VlfkLSx6SFGzTGPIkAZMDrEb+Pb/0xGNSL3Db/2PK
FXQXJgclmnqANYLdhSZGAmtWLECCjHzhzjVyNrpndlWLvbpK85v3GnlhU0+/gbvk1FXa9EC+Sfxp
iYc5A436yWQSitatBpABYtoCS+Y0UWBVSjWPZbKCkheAWekDixoellgo7hXLFmHKuUFUyi7WMQP9
pi6ywvCrXaAGV+/2OoWoyr837Vkdxv9hX9lH81W6QUU7XNzHxd1G2Crm/G93h/YWZ6Psko3duLs/
9eCt6s2//+rWyI0D4ZbuoSCH+VwbJFp3YeQNrzcrSqrOpjJ1flIZi1Mvox39ZEJtP2VteFCtxtLf
psdgIUfw9XtFW4y1s02UlGKD3Rv/XvHxl8svnT2e/29ZBghEzw4b+34z7SGqlrV9o5J3FnBmmxck
oOVqdqDJlJPS4cBuvU0aJSrjTuVQLJuDyPYkBsvGF6GEJB2eHvIWt//nY9iCYADWplc8Ygmw7sOe
4HqjHQ90CU7T8ZGgSRc0/48lOx30R/vjWtOrTSL+43LoxrOO0ftViyRR9rMJPefAr2gdUMK+zdDB
PS4OkGm/E42COWzu+U0Ku7TiVoIVazhl7XU/3gcYTXPDTXcCwFXSFoR9xE6+7W9cQRyYjPdeM9sV
kr2Oks9KToWvJFRzY+9LzQkA9yBrjBOVz+y2dMb6NpUIPorHQA2j4H7hDk7t0Clx+BO/EOET0QXZ
5SUdKeOtKS1eXFsiQAC8TzZJZgJK4POuMu+P/GvJUo1uiMWgy/fkPceXBGyzNA+yRmGGJ74fF+dT
xGnTI3qvOHb6gG058Xjh6g327w+V4lZpSFlERDBTC0x0AzCfNt7WJ753orWtBl9JRZN344hGj0qV
p2Q9RyRLIa2lVktYSws2RTg4u/SZklQYmxnB4hj8WTDeY8hKpt83t+RH3uS3EuaxiNoQTXVPXxNv
uGgz3XupCGO+EU79rHmHnV6sugGhWKIIc9vApm0WepKRQymK2xvNPUYPklN/xQwKnHfc3mAEwvH8
tPPtF763FOoo639kqffKlDV+RSbAkoPpLPR0f+CCamArj2m13Nc0rWQDqMfTFzQNCxtAMeMR92kg
13v4ghDydw2KL6ZcstkYB4DP2ZMv/HNQw/hSfkLKeC0nJvG8X0ygszZ08joxEMXoh7SoTr7R/9NK
86hrl4XdMITEL5+FvyL5SnBoF98HKIMRwcZqXJvq5LYHP6X3NCfNwOAn3hwyC3ipuanop/wbcmDW
bQdWcLjgTTp/AoUuVfZeIk4AGt2e4MPFVgEVK484L9Merl9vGhVbaIVy0KjRygWqPjUeCwGBVz6d
N+Bmv4Dq1e5S0vBdzRV/PDwk6vSaisfVfiAnjJ9r/i+xHKDkjEvPa4ofl2ehfq+RGhMb62S3CZ+Y
Cs99XmwQHtmFqqK2E6xyLj6rdPRpnkyUGbIcXWwIZGyvd/yxXcHQEXwllwUhPxra0GED7214VnZL
1BbXHDIylt6OvJnlDK/4TV+Iue7rmJ1SkSgq+H8pm7dqBbX3f2TGbxOulyrSzMoYpADKf0XjlRyx
NRTatE+aVBnU6qlIWkpZSU/uQ9DYYxb514e/CaOa4cCdQzcU+zOebni04d5maEY35oY0hRjKFxr9
6Grlw/zdEuEjli9WKDR9/pKTzf7zUXXMaxzbBgzQSVu1Bqxo05NARi+WEaGP+S1NUOvpiP4f/dJR
jQkFjoRO/m0FWoUD9AulTLX2D4Kq1/V8nrY38ZdMzR5uGGmKqNiaTzssFakp5NQXH9pEuheRD1NY
8iXTcao3kKNxEPtyuVt2hWKShxWqjy7NNjk0g1iH70xbc2TJTWzAwiPK1RmUsdIQTZdS2Sm5cXqh
/VX5VeBwUgB+9S3xD8I9Uj32kA6e/7E6e/gCHL7FiPEYUQB6DXJmNDuJRPv8LUMETTj4re8BC8np
rNEWQL//as2/k1RXM9WxJvG0+wNsiiiHFdkI1jFZDuIBBBKoxuU1akFIm+lIehxcwXb16molEith
E5rV/iayvgk1Xcl9CvVnh+VlXWSTdNMoZCRTofFi2VNfTmmY5L1MQcnpsDrW8+O2JPZbMEjqwHkW
ldnT0OQ+UdkAvoSps/Hb1tsnTXFE662eJG8xPJm2+UBHzGDrSxUC9r0YlgFw5eJa7wX11i/GLpv3
CCnowkN4TPvC/6AjkfxxWNvQs1aLHYBFPLGDzx5DFSGBRjpcuwOq9gJxdb+qwTJoTKlP/+3pF/yv
T7OEV8rKCw6l/W8MKkGPYIhIL0/gOOzLhFQy7c/1gVu0k7eviLVvRLWEa/VUH0Q4PjAPr143M3eZ
COw/E0IUa1m8PNTRvjk1scMJzVACy2L3P+YBNOAndll/ghu02g4Sore0XYkqexuEnazBcj1CanVJ
0Qt4u2zAswyesMqyasjv3xkTjK1yyx/YBB0M+YpDsfZNbcWxBS4ZJ7r8OJ4fynBuW29bkGR6cfk0
D9T+6icX9OVNr1ybiZfSFRalM3TXy7EP6yfXGDhNMEts54R17ea1NyfbhRVLijBAj0j+Cl2T3rK5
A1MVRgOmUkQl+1pfaPfAnddRq4BbDTwr26GUFeQlAZe9sgKLVVxwoIt3qjRdmg1zQYnK6ObVLKp4
HrziycLBVidLlqRqjnaxo+C8qb32/5RKEDv7cZgbF6yp3J0odcNwWDLCk6wgGsCF/yycKAyh89uf
yUm9nyIcmUwhAQKw+cNDcuAIOJnJfEQVYeZ767Zx5lrmz1QrL2fe0t8nvrgsyiPpsGrAKaHvCzBq
jufJAQHgAgpms6uti5ELSxEUj4X3UesegNvpvBuGFMxZ7r6RYVyHcvBz3XZEAtRMNR9hRPlzSwJF
9oHWTaPar1p3WO44yKn/mCDcKLHbdWCS5KYIybh9YSm/JfOV2f+id4Tg8oJsQxCmMCRqOAFrvkLO
tHTTpkdiDvTq9U+yPl19hYZSynCLYp5VjNmpqCJXLZfAZbPSVJTGFQNnYBZHl13CpooFBXioQIMa
KAIMYMjG9IRWjOOUGs4i6oxUR8C6jlx9JjYnQOAKroRwHSh3Ci7ZenyrY+lMkgNQCrmXg41+QZj2
SfdQ6bNGoofQb5pZFY6PcWK2fV4AP89CvPawkBVwc7DUL4EFvEutCe/mmcizj88Ts2IyyitncUzG
5jDFWk+BzIiIrhv6pTlxwhN9Jaz4fji1JO+zG0id8hTS8IIguH6F04V2kn3LMP90lTctpjVouVU2
YduPFtlu4L08+g2quPWshFgt+IamgSwL8qTrEqaESTDie25DPCTSVwTMLW2kYdXNcWuvQ5vPlfV1
yn0G/c3oppFquqwtTW+AoLB4pNWhafrDcmmaA8ywK4N5lUZNR+OcuuQNYLjcrFJPcsNy8/lvwhhV
skdhXUgWKP0o6Eo2T3zT51ThOnYlz/qh42FJ7jCV4RdfaPIaK2ZCL65d3F4uYvVHEVwqhDX1ChMV
xFV25laHxG3IQixC5+PFLI8SSyuBwqD9XK1pN8b6P9//kZ2oBbLVO1tLKQua0tLOIRltseLENh8U
NUcyLSdCZU0Ylk5fMj5FFhjV9hchHl9+X00WWLwXfhNZE1i9C2xMaNXK3uYSap7C9G4FPS/oiVXO
AJhn9LJBWujKWDIaz9bVZOMSzx7Ol01T95YJmoKl4ZpKPOt7l+3TOI0KDaIPnbx2YFYMk3bujVat
lPsAxpwPfQJxD6BVL6tNoeGxClU2zHPwWnbJ4SqpLqcDlU7wNjg9KwIOA5iKrLYo+kqgDVONv4yp
3HwIKQjCPJ+YjONUotR0g4+8n73jQMiCN979HcLNfvshuW/qdWxFLn3YJSjavhEX6rz861TxcXD7
4GsIax7Z9qggCWisTPb5lHQP0O7M5opm0fhY/Cm9SV1vxn48S1MD7YBsMZbUXB/7Vu3Z/2UfG5sK
APLekCtaT9XLY7L3Mi6ieniQdB3Tz9w4YX7P2e3Ifya9vm2NALGIwTJIX+JV2/+Ik2bi+x1HjnCF
j9MhFdecg9MBgVEgQjNX3dA0cuADjku3f9ehB8JBrPiElTLyTeSm1+jwWWYNdNe0y6DO2hxHEA+C
R2oDB3Pz0VPSaHgQoNEnKyFCtVZME5o31sd8alMm7jnRzGAOi/7wcUkNQPO5p6z24h2UIlOvioYx
TNWL4EhmyWLAwV/FE5o5jqoMmm3hDB+xSXRDDxb62hE9hSKTTddmv+nddwtMC6nq1KeDE6zn/IhC
aEjVIo4bq3Y2+BPIPVfdoT2Io7EH8TUuad5ta29jC8K/Khcc1bSNSfQfhFYLYHw5UpCT/TT+3luF
75RUxb99r7HG0E3kqHRJZX9a4V30HLWvtT3DpIT3W/9WOFt/I7c/6zKPTl/SCflI5VLTJMpj1aMf
xgtxMDlmDExB6DkAgIr9adKj9HTF8JuYXLiPKOzQq1G8z2Xwh2zGV9nyWrBeHSMHV/ID/7M+3IzA
IZyHXKRWsZm3eOf94K6ElCVIrobuChUVrcmep6nB+t4A1RTAHpvyVgmBycNmDeWLvd7U37yXNQ0D
6wEsbv1hJAAVeXGAtOKM2HWgEp9QoF6MOlR23mi/xbk80gx0GnCa+4wIgSLNYQNl8+ir3dR70H7w
aye35j/xUPPGII/XaEN2oYcyNwmfv+SOdeKTq6NKjB27IUi232O3wD9Sl+WHE1VtPP6qEz31etwg
l16z7jRbnaAL3MyourkSUcMXSEs9t1l4py64koLSpTE0jrmgvD1fieamyhW2HNR2AwbHO0FMEnlh
7jF5eftb3Joq2y3BIosrRE+UzZWORajn+FJ509X1NvTFFKsSgUvG/xfu7mavTvTQQvs6Q+jTeRir
ZrLXFsBLYEhS0GYKhw9G6WIW0kySCVDHLHWDB2sBIuPh3li61c+hYR6ttsvZaQJH1Q75ZZhyyDsT
fKxcL/T+l4neB9ZBsHbrtuezzlg7fa+iFYYgJdJ3f6BfcGDC4o2Wro+fCu7a4/OHew1ivSTrEpGt
atMLgrVgORCHMa+pl4Ij0pBJWZGHnsKSMFo0yZJyPIv2mD82/N8AezMxUTSlfcFC9yZAQLT61n/4
/EM5/f1V0HgQQR5phi/YwlO+u6ArEMYGClKC4t2djuQwMc+qk6jfvwyzcJoW6a9BaS8S6j6tiEUR
HaSzE9gzAAl0yFnY+fF9YhzV+WsN+YTwlKbEJ+va7s0FMY380C8gk9mQ/T8ZwYxqOrlTyUo/YcV2
Si+TrJ/YubEtMHbcpDHg3OBh9i6WzVu42jT4ASPC3NHi+QVl0rVH6bXOdGdhZ9nMaS8eGCdiHF5/
MTEzOcFzB1reHh1lAJZGbfq5MBbT7tGeC4J4eFc5wEtTdLY2eN6gp3oiOXoJ0s7TCerytrYM051N
SQfl8uCWSolkLuUqxbY8bJ5yGS5FYremjNsyb7ZakXuVknS5sv/jMHwj98s55Nb6SQ3dzBp1ByUE
dtLlrpDgc95kNDI9jY1RrVOazUHGe+OzzWYFYmjCrNgX3nXmOb1Nob+eTcB8nUwQwb2dhsgw3E9Y
wnX0XCH9Pfn0N9rXluOJLyzwiKzQ2EdhZgOZ8fj1hEJ0+bNzAxfW8ag8DJaxeGXJbY2GyUBJMy4o
BDaKoYAce8gy01zoepGR2fWrW1KBkx4PAyx6LYCBBP8PPH/kQRVCJuYEd7P/QmGekcwdV4m3AKRA
AwnlneREtJYZch+MMGk8ZVGfOVOKdh3Ts9h7x81Qj+SIghyZ592Jeq2o6tdt29k100+XaMrsK7/R
m5WGIrnvG9NRXT7BunL4sfjfIukXqnpYMtskhPIh5zJvCkMDzvUMOBYs4sy5AuQ3ekBYF6RtjXwc
8RfS1zKgRMX1qSlXA1Jv3r5ztEfO+pCxCeBXZi5qXuhHia8R3A94BMrOrvL2IoIqSiJzjKloNijD
aQv1wBNaBZVZNTkdub2/JixDvsDsQkkIZnQ/BrnkswRpVKF/wdWhXNI8S+IWvqCxQ+7A+uR0K47t
YnvKD1KPI36Zv9pc5U+J0DPPLl4eVC3OmUKApcF2LZvcKbsXt+veQtf99AnM7zx1ywoZL4PXYnWe
0Jls2xZy+QRXLRjL6MYZ8WE7cTkAK+qIITXmH3GpuqefPwGi9kX7mZulil8AS6nNObRF22Agu66t
pRmYmFVrK+G8jTv1XSjEB3QJ5wXte96laC4y/7HtKiMWY80MwMebIkYDdN3cmxhoAowjupgN+/dr
DJ0uQQpXqFqNvg9WLM5LXHxYzYn0U3XotkSAiSDsWTrlAp+f09AchpE1nawXRfDUstG5Zs5WvVGa
NdFhKl8BsTtfQ7lVT9Gjd4i+IjTC5VjQ4yzJmTuu/C9oFrMb4AkRRfhzucg45yyuN5Bm4Irn+AEW
ESbZnV7V1aJaB5z2r1+aLl2PjP7wzEmZJ2Kpehoys3FnfmgIYh2VViLeCpvBrsQEp/D6yPOg1upn
jhZFHBn/F2XTAFkNskr1Sk+7s5xkU+cOzm+dS4oiuVVR9MtbSSwMpjaGHSbmIv5hwkcZ9Lz9ukle
CswY9Xfo7b7GS311t8Io4XLMxOP5cAf1x0XXp82biYxwCe1Gl7DFmbq0K2408JQh9M0MLfSTwbCz
SJfaN+sMe50F+Lf2PMNJyh993q3kFtGay/YT33LUqsiVCaJr6ekOkjgwyQ9XqwJh7seUlhCtb5vn
8wmRwoLhBvcYE8+0Ttl6cLkEOLkhf5LgN9L7YzBQ7lS0c6JNG36cFjSNqQnHxXj0hI6AtCs5wxj3
E1GygPnW/W1CvDP/Own6kt7dzmymepCfpNi44lVT4BYp2uiQDiGydwzByvaR1YeDbJ26N0mQVDug
6lqH30UFtSJV/1auvHYgk4WNEHUQ0kbSk0/7lEZt/CIBUHJFcuxPVah8z0MaMY6JU9lMb7PHDH6L
pkIpx6ciJ/Uoi34drlo93fwvOncWhccNiSfEMW/+NnA3AnCUwMhFomtqM0zEYcuWfohkgTBuTuXH
g9YwAmOPxl5veBeKTKSC7aQ+CLq9QXBRDy9segZcArCx74Nae9lUHqGfKlxIN74+BzqI4cQPHkmD
7qRNFDd9Y7OO4Fb+TSaKQXBs+4m9tvYBydesRIuOg/3AelahdXb6keICo5jUxOHpDEc1Dorqrh1a
UDm2abR1bKgqLTa7rtF4jfKr/oKEj3iDN382bH3j/znyu60+YLm2Rohc2yIDBzpZtFU/L/3QOSaS
14uL6lEYtI3wLWjlbSCyu/zs8aHv+lmJOdGL/kz9JBef+zCU0OBco5i/QmSbz9UXTBaooPNzIhmc
cTeZlJkN2nLiVZMH4daE5XiGX6/4gSpLVQItKLQO9L3PxL1+Oz6tAULQ73Ysk/ymt9qCxXpSj8BU
HQgIVRT/jqs/m1E81QNWB2xNM9m6lw64FAosSgtfs9+OXDua5IaLxTYfZRJhP3DyyAvEgoBjBtf1
/VTVCTXRllCHs0E2BSjkTAjj08Jr6HmBKRl8UdQQh6r58W/fQHZhc8oyCW4TGqHq65m+WLkMRkIb
XqayH83M4g38BDNdP0HzxKfzqIkZ9OOS9iuMXxxNAUHZwVhxyc1c9nPcL985fJJ2zhCNOkrmGOlV
tLg9XGzzQcxtmbBPOEP5N8diqwJL9uHvQ3537z2djR1AbM/45fXq0LWYUEonVo8t3LFtYGhyPgZa
50NmROznxFJ/D2dl7QCvX1yayNSsHE9Jx3dHmVOzWL0jYvx1jqEsFoozCdDbkwGiWUi1ydRGY/oE
xJEZd5Kzv46ql9AJ3aIBmrloVHHlwRNy4SKaLGhB19Kr+EWopG71Nm6q36BpZcFLYhjhBfeC65Co
yu/6lsX49RjcBtcuyUOWxwp+zVWLjCHkdlAcIMyDdRAVAHUqmVlxs46c+3Ze5RUcVCzrDpmyoePR
J8k4OpM9PlhGbT21u+H0f6no89rqc1sb9TbMh2GG2HmAXoilELGqdsfIAhZRDdZ2F7GkiAGmsNvp
srQbKCwsDGeIDo7FJh5G8+QnMmg/zOUi75+q8VRhYipQjpCyqdHQA0dviXh6rckZnXKFEqc3rvup
jIqRCaZUR4MykJ7cAFU9aiplmaTj+9N0XyBfvU8QW7UtWrr3t6J9iVfuEgAJUKJWqrNLORtnrtR1
DNQve1fxxh2E7pMCtv/bGTuvH2N4185Uw9EBfPuPuUT1zB6Xo0khisUO7BpBmYZDosWVoWXjfpTt
VJedh8dXkOj6TEU2wQj6SM43kHlkIyMF2ZYE5wIKjGpVsXNv94ewmSx9RQx3Vum/vsrNKmmSwr3A
527HwThe0wIIyofQ1mu39HVN95IMdjBGctVd6konHIZ9UYhduq1jcz4UzNKKpWOSEQo2qGEAIlXt
zO6joGQs5td9+uH18IMehqjxJj4ge1XZIC7ej2gCuqFkRDGDUSqMqJyksEdWexQwf0XSOWc59CT/
pWeJ5TRZfvf7EJdooCj66liSbFIi2jSuJePw1LJ8RYykVEMnY1fHc8UyI1os2252IJKkFMZigVf2
NL7UrAr2u6z/jSTk77yK901Dl+CjNY0X3eEvHpvcOIWMuc9dKurkZfXUpGasTgOeae5w2KsZF7+A
VZwRWZndlJeo/0HkBpq4bMLw5Z4rPR1fofytZ8T7ZFAIr2Cgvsk+JugOIJCxfC9YkjXjg/6cgzr9
PuAnGxWpKJtseQNCCvSgl9PiaVuyReAvXGBToU9LUwS3SoOnuPDrfQUbgI8FdgTXaMw3eTknBIeX
IvU4OVyBaExRdVkMy36oX8ScrJVDNOdJrRFfYTJ2GXQ2LEFCBjFh1Wkdow6VWsRMsMoHQgvDC0qs
+tg2N0mRXW4oWp+R65tgObbBmEl/RoAK20UgDfVD0O4JHeV950EEQXOyh4M9qKktBxZqqNgfr9w1
gdQ6Xe3Zg4u5iHQzlxJAntTZqn3udn9aUc9t77moDt2H7sEtZgyEvpCbGN5dVhoBjk1OAnIC3HdV
CuHVLufjlJVEuzgQBQ0yja8PgMQcrbj6PmN0njRJlLLlbB2XRvzfwvF2CGgdDuUG4qmBQJ5rqBVx
XVj/VGSgQ/znnYOgW1Lly9C+8ahgBjWmXe2VcD5ScMGmB8ZwaOAfjnPb5+/4/TszjbuzS76gptdd
wmRm2LodvfYzCFzvFBeUhz5d7nzPjXZhudF0GuS2MqY4HXMSCYJSpfr4JSDHehGor4kaN7WlJLGM
83qX4tn5nwRDdfzwRgFFBzgLZziT0LIA5/p0bm3kdVwCJ4e6gVrNOzo2h5cYsQrNNGx1Nin6tgPo
90ToW5VQZElzisbzfLGtDBJLQG+axlmE39YOo1CwKCl7KGGV1nO1CTQd2o5WkDDsQZAi6w9JLnjA
FuAZPftch1b5MqZellHhol5lUPToPdK/9MZLlOscAy5BGvJzs9G+SYumzc9w3YhOaGSGrRut0Lu/
1/XZAkBPguXsEg/ccY8rq4aCHN+AXpXRM1UTJ4PBYZODVNMD8IIOdrlDyG3Mf7Z+fQMtBfXa80qs
+5cS5N5YEj5BkU/lqNCOoQrK2+P6QjQBIFZ4gCMokRGI45hBPtxfwrmSKjS9hfiRv7V8TiJLfcJ2
6YTyUl/TD7XrI666oq8TLAFKv6oOZlFQCo8dpBq9YEZRrE5XmhjAm5N/gFZ1YDO3TE0Z9cozXo78
p2J5kaUADUpuTFY3GiqrVpxA3R7exFCqQiOfB8aFOVlM9WNwnki0YF9LJ1TRlP4HMZYECyJlsQY4
Oagv3OQ6EPMlmXO/rPQbR8TTyQQkT92cqX25xJ4QkNwyRYfG43wB2petybXDa5XyOHLVCEilyHmo
Xrbf8FzZduZNktnUHea1M+xjrfyIxts09fboQXpwYr7T6EMS0ZdZnPHr+8YOzZmBdUhXBvGX26mX
182UOmvgWbRteHLZAuRUK3+RhF0/crYJn0ICfpxKUrxo/In6Q8WDextK78w6ESQsO0PjbT17AC2u
uPKsL25hJYYsQ1QkPCV9sRq7HVjRmeP+t/XynEE8EPXkeiobiIp/y/5L5c4XE5vAkfqTBXkMWeLn
rMn712G/rCOoG7Oxx/rG7XzgCIcC91HHF/YLLpT3Cdy+8dokVpE/CU5mba1jeMVKrv634E5CQX02
TZT5j9tWzoo8dkdWHN3ZSK9pvXKWkfFGEaYpiP2rLQOxDWZxBKUqJyZ+Ei6JaNOsVG/vR269R1N9
NH09qt3reMlBCkx0ktSVOzePoq7w+uw1LEc43A5t6ijX+b1RjoyvyLCqShx0e7tq4PPXhnvbUAFN
0xZO85sM1c8vSseM0WEf1p3gGUlpMIUeZxoB88q3jV4/rCapHj2lygw/o461ou3FZC5RPB15Tpnt
LyaJPckiNg2AmacOy3CKBfAUQIcte4NQzInFw1GAar4ERbLUkNvf75Y6qPTunySRyeDu3OpcIczT
rscabm+I6W0pPT6jNTLE1E9co5CCHMVF79uE0jCmg82Tf3sr5QbvqzOtiQjplhNdvcQXjJtPHRTN
c5X9lBT6RDeClBLtS7X+x6epDsqzKt3y44BFt4ctS5Oww6B2cU0AtL9qf3evoh9166Nn+AoqVY24
QzlWyv3Wf0hOlvDKzNiu93ISJKsttVtbKn9RDSY41JerumIhXZE+cy7rr/rVajuxprUi4ZMrWHFN
4zoCI4WfktYHxdRV4uwrPAda/3t+lUHNdRwxWewJVuhEY5o/+iLN4ccWwETQVx0GdXU9GWcBIlZV
K5ho1Pr5dS2vz/pq1l52lb1b7WrCWnrHIT7cNdPdomLtv7tlNbUkZ2mMotMp/bQhEHaPW0Y2MRN/
Ov14cG0poxaTdS6uv2Fl1tpKoDhTn8LveQc8s+Fd0cAC58cBb+7m2X+QUUekIKf0YbaG9sPIEF+t
hHD42Ci/NYTFgz/6d196qTsoGGjrxBsucDj6J3l10lWqE3QwM+IhcBnlEIGMynMi6amYGSiLhzZK
GEmywCr/9o+spoOn2LMwPyTys2RfH+Bur4sfx2Abc+N4N7EumUABox8+URXyOtdk48kLu92N4Ed6
X5VR5I/KxOd/MnGD8Mb4yp8ECPGVivKu9MgdaCTkrt3qskUk+PYvPNE/TaY0C+Lm8X1m8Z0OAGY4
QWvJF0Q/oHuTNOn/pI9d9xfOy0XafGHvrKS2Z3O6PdbxIGmQYf1jRaSUlYhhDrSOxpw7NtFmVT2o
n/kctY200eSqBAkKpvxN5w4vK77f60sGNzWMjHQ/j9tA/ppRsHKwsTU2soMzv0JwQdNOGPsd//ge
skBBkXa7kI9FSMsc2HTId+yeN4g0qiLRLOUezpXnlL0hYBXobZ38NBYrtyAYnbiZo4YDz3dIteoK
s9qMHidWvBZKVzmH+EGgge1HNgAf9Zfum37vBzcVBsKzbp47jS8Ld/wxuiCbsCzngu8H7kQBaONC
Teb86iGIDuE6y+zzSKYt0fC7IEBuiwedJHvJZoqUCcxLPRYNLggdG/3XEXwBoIc6AgXa/WYd1Fcz
YfuEirGojBWEOldZRhF2lV4Mt4IneECAVSLAzfeGaKrWuE1AmfOB6iYhrlU96rTVJdlFFPvWL4Bx
yNwI7bsC5LA1wvWJmNmP2O/O4amhPxYg+GTtBhkdmX2m5q9MIetVX+1W8bJoIMIBv4dv5b8C5U0q
a0UEJ34bYdPjx2a2iynlirk5HiU/u69L1FiMyVua+1wn/u3ctdA2AsqdsvDfcRlW0/JHkXi4AmLG
2yJMudDYAO/H8/VQluQGrthCUTNHIjDYqGdURNo4k5iVUWuV8GS1oQIKrr7mD1/N/7bEOPLst3NC
3dqb+wK4n3FZRUheoo0Vj1fDshP2JVMAtTb0djidDwokgLVh/ziTN+0BjGzybZS0kLARnIeAkrk0
BtfNn41KcsqnKbK91k6k0LXrwYSF/WFJyOaNMMqn507hLoJSjpuh6z69pyaXi3EV2xgUK4lOum7s
zOEV8RiX+V84bT+adn7KkYMoZj152p0pUO1Oy1J94pN/jnCd7hY3u6WCy4JaC3SN+AbjBkyuLSTu
QXV6XgyiYDAb0yMkJN+P5mXPsl71Qmpvx46YmimAofhO4FN/0VG6CuAxv49v4fSL2iN5al7V2e/l
AhFLxtLuFlyTD4m94WX2V9jhmqLuccCXLSjPu94FPxb8SqHE6leVT8CP9ORSFxn6WVPgTzlee/Iv
FgfjdB20HhzjPn1hOblZofRWInmpozFhEKv7wFEys2oRjVe14x0GKJNrEnsZuYygqmIvOhfoQjyz
TRcdAd/V85pD1+mjRe/hUIz1275rLd32+Sc0zfxy/4BdUmB4SZchvNOoFOywm1MZGD0Qj4PDTGU1
Fs716uF4zjICrTwXb+ntZsKTlXsJ0x97uYiQvNdesZzBjJ3evA7wV+9jliXm5+sN01/+22xMKcnQ
K1dhbT941dyxXZwpoVKl/E7XB+td9Lz4y6g/7mNtYaQVINNYCili8Ck27t9hyfLQl/jMiHuip0JG
4IssQhn6xlCy2fk2h8d8pcT5wMYqUKsy/QRY9EtoVDrLiDncof+QJ6MSX4kKYdUSmy3Khxo0LOvd
w+9bMR7/cqXFpLedjVbJfIR1epjw1NUGOkiMJZzIY92lTnaVuVVbNCaSItoRg+08CGsY9bvQ8mv6
YAkq1qrTSl6hxeBiPRptbVLrohkA91aS3GqChjJYnzkBf9+1p6ZFGMVZow9NsPfkM4kstAcsStxE
q1npO6XqBuexKbxs7btTYxLJRaQIyOQfn1+lAe6nw7pWta9Fz/CNn9OvQ/Dwc9IcLvSL7kk/2szw
pkgSoV4ZLn8tzkA1yvd28s/Iq8TM0q0UXMnQSwx9v+iPOWtSIs2cWJqPQa25tD+M80qLEcZiD4YZ
FFLz5AE6/VsC7WmNfuJQbUKBcQuym9NaUFHD+1R9bK2fJqagCCxdpblo0+9fQF1bvZdJdb7fkX3d
JP74JI9qhDoJIkKkuZ0UWbZe0Onl4QbO448UbhVaW9mLcm7vmLGJq8OTPsmtUMPSDRGML9528+ys
XeS1BJF2CfHijNnwfR1W8xEAqqiKOKcABjgb4/ZqVrTPSIhGM/3R3oEzWU9oZXkBUOpYS42fO9KQ
fRwK4EeZsjNHK2UsugdirmjdVFqBE3I3x2jmpgEIAODSZgx7kxJwmocuKcy6kWGX2QWCPsKFTevC
yItLSGvpXpCyTBv8O4SQ9cC9yHijKyNhnPMvvxZr8aY4+7/znZ2PDZHUPBgDtjoQkXwGLnxQV3Cu
KDfhCp7qvWLbEb2FydS31cKF8a8JWWHTHr1PdIO6JFbIlejLxo6n6aHhQNxfH8saF+zMnAr5Z5Gv
ELWMQ99WmrDcR6Wt5AJDFYV+aqmBvh3WqDBfiG6+fRsM+QKOfCmmE6mtOR1CV6negTzttPzFALlz
rKCthNXHOFlq5Cc19jdzUSzNE85Rr7Ev4PEqSTOTf31LSa7YP0EloSWGSmllYcTnxgGbSDm7PWoC
lb4BHsU45b4W5paDYSWZymm+pWiJJubjI1xWSprd8k8J8wjnMn4MVGYXalfjVR0xHNsHX5gSON/z
RVCpQRY1zXYnch/7pwEgXG6lrB9oLuZjh9EarOfqEHOL8n2kTJn6ypJIBpLg4a9xtNY1CJTLu5uj
JN1azGyOBxjIjNMefSIRWAA33gFMZEnay+KDD++VgZSsSGqyh1Cuvo9bKSwV4PaYWH8Hfk1rTCRL
91KrBJH2wIJwGEHgFhJx5ygCBkpciazhhZZz9iQV+FsTK0QSvovXK98CDH/6EzvpPE4wUKG6qFzS
miGhUXOu2rQDpGwkUsv0mRAcdvsFuqKjNJhiUuq7SSIGh+vHvFC/xF2uXlQWQBW05bUHrvvxJktY
pwO1afuu+JXxTcgKE6zrRLFKOGdtq45XDzUCMAemo571D8hx2H/rR0EqGedFLPikSggDy3jvfZsn
8Tk4J4BA7g5J5xmlwsZpbVffeJYZnw4G/UVG0XWIiq3W3mQeqU4YwgKEzoBhkeLcr8HaGedODeh7
A/7fnJDPxq/p0tBwhVMBA+U1Nfnb3f/Tr7g5gbdccsp2wgrsZOT+ITaF8ZOlAPXTAt8cJFG3OS/d
Fd1cikRJ8o9M+W8jgLsgUbZWS6u4vNSUAZSYwEx3NH9r6XqVHI3Lr2ooyDphTBEO0hA2ZOU0kfCY
7ErWlN3XxjbICEdRg3traBjI1mwMJpBcB/EN7Y5bDODudcj8/6Rya8glKKmOkgPthcCaGwJpkZ59
ABClkI7jEam5uUtCIC6vuvFvOjAtzDmeEadXOHDzzsCO3stKRJ1/SPdxeD4JHU1uqCoSWeOOFgmf
HBhlAdez2z4vf9xUUzCwl+OvCXw/B4SbbTo7Ib4qwx0Ckxr5wbf4bUqkqr5devYyoZYhXm93vZlU
NnfSGLksPLpsqzebeORdq0SAww7D+00pMtempgZPuD8RF+ysriToK9C6tdY6BTafZTgx5VA/X4xH
823n5eR4ydTrIwoSQLInFlVv4Zkxzz/wD5aM3MLJg5pcbE3Nho3XRV0Jz4/6DDZ/JcW9TQWEYSk5
SxoGeDszf1Ekj+lQpM0E5TkNDPi5smsyxI0fGNOpeqQQl9NiWoJojgn53tQoojq+X22RcoeZOaIi
a9kmQxeBzwnqlFk+zyxMwnuH3MePYSt5NKf9WLltR3+Rw+qu3eN8vWLBurvc2w7mQEAmtf70bj4d
rstkRwUSL+a5sdNEGwiVCfxo5zKgfCdlLGSdqUcDYDELCUewxKFNwywLiCDOxObAwDQOXUmodXhE
/amJl2esBz3uX0fSk9i9J4VlZ6ugy0vH9e4CxbRiVaea4T2r29aqLFvGEfHv1sALcouvvDHbm1Sl
vB8BDXAJO2co7klcS4ASvu9sU/uvNiWyTimVhyEu9Jb8QNquftOB2TJohpsCHko3NbfNXoGbPFSs
K3zO3wNmxKDOh/CE25WrmMsqE/BHOCKr63Php0QyVurSYHcjs/HWOgocdA9YYUZ/EiMy0wN+36C+
w759wH/BpLRnUD8XEMmcA8bNHa2hahzGQkW5WQunmdAnQOCpytMXLhbA9VAK8WUVx39B5ytg2fmW
MR67UyHwUhy8K3N+js1gCN9uke/QACMBOwyV43lX9OiA+Dw8EKwwRZMAszysziKbD5RXfjQQaKaa
00+C5Q4I9pBZcqV4exwurZHxhYanENE4LKMJPx6ZHlBp5Csxmef4MID+GmSNR0fL5gxJ/Wkx+Q6N
ZMP1cuPYIXRcHa39rmW78RccMANaaZqE4cBPoXoS6xWmeahmNIdf7lcqnM37Y9UNdvmcEiDlEcg3
rjCzlQQ1Cm0U+Jn6CQ1T6o9FoCTZF7YMcYnpxcGhCpRP/UjkGK7pXGYliOCNiW7CqC+PGvdEzGaE
MRsdCLPADDlOTC28sJhx4P9YUXKkZcyFdY7d+pKT1rgQ0L6J60/+cGyFoFkdYMkQ8WzR1wlRiNx4
n4jlFCAdxD9wVlXxAoGjSgBb3Iqas4EyOBV2GUMAdPgu1BwAiAL2cDUQnc44a92gI6OnJbtgcw6b
SlLix9hD6vAzJyitYjvjCnIm9Sc7I4wky3M+w2YRqjpYmaEJQvRMRwQTAkfUz9strYSGgVHH8UON
qAGbcWyvSzqXSDEwbtBImMLmcpZ/NjgOubVSmNg1HcIuF4zINeawgKseD61insGBwVJRoikhcTL9
BcM0BoeA8382g25J7/uQRjqFLlDpljJL068wscplvNyxfN5qh1jwdrRclDLPiFWJ1pgYocZpyHNp
I9mFOEJCY1khcMawV/mz6Myht1UTt01vvmbges3nVmtbmO3VlrO1Jb+GeoEQRjBOVg+O4syfIsms
MxsTOk5wuWSNHAjM4K645SVECFZn+GNcGvIoIx9NzZGHpG6qWz/l5jEdmLJqUunkDDmPLzPdM6aZ
BnRQE6U7gov8K8LpHxzVKmFga+Q0SCmhai8nurXH7umkrGI53VMfEzqobjuQrDYfcooNJLGnDnOd
j3PFRQmWNMHDPCpR+ZWeKx+ND/E+3uOAveHz4Wg6SCe8h1lppQIW87CEzmeN2mn3/lrqGCGh+XXQ
djlgjAnd1zcexDPfy5mJwmKmDw8WDP3a5Azyzd73C/zYML+KhnYJr7cy6/dqCp09ExngUzgr/3Ih
GCn6qm5GQwcyEZHP+Y4qI4vomsPKVSF50Zp5ltaItJ8+1bp/Xn/WjlISEC2aEVVtlTPdQc9EfGkd
bIKQSc5XieVYNtYcYL61YvREE7wmc8zoLXzWJjyrm4YoakT8uhJ653SiULraH73qnxFQ4MTlhcc7
Gx5eZIdjVVYyUiiZQzYwGDiBHR7B8Yz22meVczO47RaUQrb4WW2Ger17qnwrfKmiuAaBPn9lRRNC
x43Y/y3CC/d4aG2QKwBIcc8JmX8wOvRN1+Net2VrPElOcrIjKllnR1qDtFNQMQ3NQaCkS6QNEgJj
wdnFZqFvd3rrL8rlz5pXcKGyl26+nK7jfAtX6x678itizPN/4eoQixXvwDRr9od78oJmOP/NIC9u
/ZYNiu1j0PWS3cbcz7dw7/cDgXncVppAv3DKxbkeqKpsEnaB9sZgI+Z0g8GtxuJ+E1lLljN/f4zt
m/fdI93zrMmEzU6wQK0Wf8e3sgNyNCcjL681AppxveVlzbuPKBsZINsUZqE7E/iGtLB3EeWg2UUw
dOL0UFXOwBI2JEvndmmF3luV03qAZemxNMunkNqFn1Gzum2w6kGa3/FlJwi4FxeEhlpeJVsiTR3j
bWWmeRny34GLFZZPzi2W2u1NDq5hWouEjU5W+LhBYvuJBEbRxRg3ClvmO7b+S1K2plfTMmSof6T9
sH1WTST/zePlbJmebIbZ2CLiZt9vubN3u42thguQvfoKR5aLTn02+nAJfAeoExA/9z/kIyM5Rzpt
euXLwh7zMBvZgiZnI8yHGnknXb6lZik1A1hD7lZzcOchaD8nFExGoSu0F8k1HBi+DmdmOKnn2OGW
qxARY26aEIe6GChbitLynduVEI7wS5qwv5zQVmDftm8eyrM1tg4ebvzPyBQO+k8cqZ+bo3npt00g
hEUZNvq6cAg65yOoD9Z1QfiXFFqnpKkDeatCVZS/VLUOMYvMLXqi6nf2HWvBlK+t2MmacrekY71v
kFBiJwsX1NIHO7Ba2/v3sIavuRIFG63Xn9eUhPqWAIrGRV8lxulx6vFweYX6IBZPzyILuO0JfuMv
05e2ZF6Er4Mq08p//8WrweXmCIgEYv0C6hHtGfdv46g9ruSFAx/zBeGbs03252AG00n6LP4jFNkv
TvD0vTAUE6LD/s5BJYvhfjuQqiF5WjlF8LTOuw58YXELutTxVgXtOvOPuKEyBmyI3W+emkaolAlC
1Uuseg2SuqiBa+WF5P7dhb3A3wNt88GcUNVOuxPC7qic0aY3VZqHKmfMae75y4CPiAw2CZP/oAM+
MtVYkoRdx5Ti8rEB9IHaRHJ0n3SQV3vZS+NzBnROem6UAkB8vhYKTOHOxcWkFrD6ryjeoQsR7KwL
Dif4gJNLMK2JeUrHUYKYNBh8E71IK31qJCMLX55NIAvzgFRTJ2zyDNxBy5lCaT+rLmEtWBdRktmQ
1qsHrpLe7k4wKtIVt/SB/Wxr6Fyn0EVXBd5Ssu3Gp0qBc8wewqHB3SjNXIhOpZAflNEp/fVK0r6f
RsQ+Pa9DGARUwRZemdCqcR3fmj2NeAo/90LktYa73i0WvB4AQt1I4Hx0sk+6XqkhKtTxzF49YNqh
XWrdL2jDI1GzymLMBBdNPGwVc47SJKfL1k6nFKVXefoCRztOtdIQ8WNK4dQS85IgEqIhAC8Lwapx
vUyd9skLU4fFXRRAIDpKgZUdB7WNlcY5QOc/z/pbyWoWJng6WlmhAs8Q0lWvbHiFdq6im3J6zaqB
oO0aQdyv2henGg/mDEOYk2YvvmTb66klY7EPbAo/4OELjGczDM4YCS3ivPUnHLmjfVqk4wn+a8Xx
uFEbOwNREvDqhgFaJGNyhxNs6WODacegHymYK4T6qG0MQTSF7dAMQ6mD2M49rSFXieeIBW7UlAh2
UCgLO17E++whF3OWyCIIUAXpNpBekiJ7Pw46XHjSZZfOqNptdoFgo1jV7PQpnY5GY7BihoVLmq86
OUzhHFyJ6SwY/CSLfa2T2hFSmx/hJ2fgD0srOckPXO3DcSHj+AcAfMmNQjB5XyFgMn2C8FdvT/y0
hn5S77yKA5gHbk1249rZoqEEpedcatZ2BaT90Re6T1w/WJo3Oepc47HeW2zKCfEE4KLpjDN4rkTE
QkbbpP5duhChxUmH+hcX7wLapDgq2K71HCM0xcaRKa6FLRgi95bKwmaeJbUwAF/ggRyYhJezoODu
8Db7oBTvHD7jM22CJ3GyrH+ZMIwdDvuY41eQKn0QwiiqWI0isaFtYwaAt9nzBNlRsamXUVMY05Dg
BvFXrDUg+62prnw1VItcxhWqhG3kUMLEi0xygaqFmyxljlyp4x0CWIpmvjWyDW3x3gAthqJeOtMn
aOZnv4/8VO9uT/LpwveYCmGqUHVxQhcK6cp7Th0T6/lXSQyfk/bzN+aIoZGrim7SaG6wo3TCIqEK
qSvXHEbRPhTgndwrNda8zJ4Z0u5h0kbDOJ10tihQumPuIJzRwNu/iYz7peS3Wd0Ixq3XjZ7JLh4d
zYdj6MrByKz54Ox+UMWAA4Y95+ytYwa0kMjmzEvHZoRnUjl2f33QqASzP4DSSdrcmWPS9INxIxQW
rmmHHEezmLbbaHjW5wi3DDTIZLOdMfVjIkh1PZ3QE+QQ7CHE0D3+ESlEgIkmRJNhSD8gKgDcOHZZ
/bq8YuFPFWzhohTjbZnMhTs/4vz5LB6n1odoK+n3DzMPHEcYNbH/acB0JMKDK1EDF2hsEX5ZUmnD
RMAb24tVZx41rmrgQCJUyKFLNrUi10n2ZrKV9kZofxO1fZiVgHvU/VJZuEV9golNzvKI2wqVWmXa
CUGS87v7iamIy9HmKP7FxP84Zhtc5BU2sCjXmkbJkZgecf/LCZW6OFhm5BYyULdjJ9k1PagQz5Uh
FNFjHQOql7D1/k+ihrWnLiMdx9RklSmg/RHzijjpin3tH4NnJEmkgVkgfBEjpXoTGCB4LC/IZzqq
1uQ8DaWFBgV/HMxFRnWLcTh1zySKHMaKWK3wkmVIe8UAi7CAbGB8hIM3ZDQhSATD9q0aXMvmcFLe
ox34JdtAM57YEeuvUIzGwDjELs4NG0tA6eY+Jy3k8/49PUc8fK6d7MHlRZSmPvrRdEounCanp+Uy
J44fXxhXq9yPqaI2eYLpxGTiwyNXkbpQDMERbAJbpCtI4XDTw6b08RFPbMsTAt2zoo7WbRr82igO
FyyOXNhi//Kh6IilaHE3vrtdAxzL/PaPL9hauQQnhBRRsOInWMbiwLm++9siYvWtb5IMGAt/Wv+3
stZgXvAx3GFMA6rN/VYAr6y2aRZEedUKkaAUEoV8VqHIdPsDCttRuiYJVYyaRR1W06gO3cZseNE5
zoOS9W8XV5BRPRnpo2+leTcKKktV7JOtibZSY36yIGf4uNXy3Vixoh3j2nWzx7tDeL2H0pV80Ton
styf1DtFYD+Qq7eyd5EfZP+GlAcOMPseYIuwzkPc9ajOlquMSn7gRHfxOz7gaDUO5+6S2NAPhUgm
IJYeob6tojC0Cgqrqc7W2jHmICiY4ZRuB4+up2sqQT/mo52/rXLjsjE3sQEDJjokz3MlkJ9GXys7
QGl+cYpfSNkFLGP0u3lcLAcZfvEY9RMIIc3puQBgUZlS7+/F5zIvuQVnpGqCTfpGBdFBcI2ZlMqD
R62OQE4XPIRCYKnJeTzXDo2Jn0w/nbUKNcTHZBoHmJcmNczTC1X1XJmHwJX/SasS6u0dbHkOJX7F
N1vAykmnKzkRJQPmNz3YxZQH3n2OSUYo+LH+PqS1fWWFGQ2cPgcpJribHvCLCIpN+T5wp0B/CE/f
6k8OrmL2OIoEYjj9QpOTcPtFehdSZvjg/JKh789IzMQBQtesVN3dVl2Q2QdvsZV37dXscTVU8UmQ
HmhbOKfB2OOVc6ObfHxDDx6ZyeXL2BEpl9WaCkk6EQ83nFXYVSptxkJjK2SeTX6/e21WFSHiSL11
gKXpwc/2tWwXtMrz04DDMHyA41OSHmi7Hopjy2NbPUdsnOW1PUzg6mDq+l6fgTEaKydl9A60dG0N
B1hoX5ebyQvjDgkbXuiN3f5n4iMTTiFqXDh3IAjRGPaOoqnwOV079RkG3QihnK5qbgqEXKHmJVMV
MrSOS2eGbMkBz5VyZKRuVAS8bPi4RsIf0rcXV0bh3CqoLM7tczg7ZiZtzL4YAj+pOtTfTbImGTWE
jABp46aEfFsQF8f5X9Xc9P2AtDHve/TcXHs0tm3HjezC9IH/ALA9JdplZ2Cjpa1SpFQFZBrgl7De
JadDezRP8HrGl8ZcyPITktvcN+0+o6170/awaC6pCja48hN7SKSJe0fKdWQKYcbONq4Xo7BiYEmm
HSMjDTW/QpLITsF2cCueT+bEhbH7QOrj4VTPaSRvMKG6HkXIdklaXVWv7k08z8iFD4quZY7iTxVp
9gGEfHZtdO0q2ymYolTJvL3SOF46omnug7Pl+NaaJU/5gEsT+Sm3QJThewdPOZ8rLHy+VA85xjfb
KWlpGUndCZUvm7ovYaCCwkfkGW6ZeGoMCugIKzdXw1G7nAOA3uP9yZ0ix6+gytadGNdrhCspYtcX
0HYjYFzJbdXiPqy35GF9/ig4g/wJfzBPSXTYNCUg7GqIQoW38hq6jVErCuEvEQOFOfaS3pMEdLSR
jmK4GcuRk/0C7lMr/RwHWy+Xs7dX6Bjj3i+bHx4Rpq40D1GXjDWUHSaWoAuXPpJNPPuRlGWGKwzS
nfkX74OIxJv/39jcjjoxVTvpG+Tpk9MJcWaYBhVAe13uOZnIRBdO0JPjAhQNX4uXGUYn+RYZI31Z
HetFVbWRyhjJ20sN/TybEXJRYRXEuAdOtm8dkoltvhJQ2nJVMsca5XXVdNhGr/NOeOblpkRaMpPS
53B28m+0eJcyQ7FZRv4Mv387CYs7lIHxIiagS6V2JzKziESPXo7fWJLV5cVw9cbjZko2eGkJYFd7
Qyt1utD12d37hBc9IIVX4JeYki/7AYRm71I/Uy2P4A4vq6jglYak1SfCKQAoayJ4/BGJzWd9GXSp
YWJON0OU61rgrtBFGs5OnXeBBRQNZQNnvTqIjyKY0QovqNdIMvnJ5+KJhmpy6+bxTGzrR/VTffUk
7JlhX0l6Pdrrt9BYImLbGjdjeaqF/D7rPt4TuZiVzb+9xzy0JIBNvw5SF/HoIRNsJAIQbvboKV9w
D6C3hjf1siiJwIpjiJL+Fc1uT/NAWIq0b64xir/+qTRF/PtVLw7yls2tF3+m6lt47wWHrCAq97JG
iJawRxr0vza0sG1hQ1x1lPMhtkI6OxkGRmOQVGfTH5/w3CfFodoLyexk3+G1QkC+fpLf2o7n0uyY
8MxPSF2peeE7zq9/1FQlqcc5E34GIDQ3g5tuWXI+yr1POjVnAs9Bomn9Ndkx4FHoWVbEgPb40yt1
zlQCDYEISqmWCYyxOXO1tAX7C//wU+wJLlTTqYurvvIS4d5n4UBnLtIEpq4MUAeuaIT3PBPuGHJo
upPKmAD3Hs22kE7asJ4M4Jx5Sny+z9/coTi8+IfYG30qNnanf5mBSS9bLs3dXSBpah8fgDNMunga
F7qyfj5TKXjbLt+ji/AH6RcxUVWuxhdEUqob3/MwzZyjdagYetIWcX0NFM/JekbRhqfUhjx5uTRC
KYR6I26pj0Dm5UdcfvNH5xqkbWUyiHcTChZJuN2aetSlWp4hlcFPHVctUtlign5ONhdm9nf14+J8
7BxNBv0YEJjGUowIyNAotZ7HQ21S4ZgHW2fYyaaJFsxhmK3eLkvOZk7/DO4rtIOK7ZB246ylMd2A
KtAdNd7au8hKkxJzllDfL/w3GwSUKhSV4oypw+Klx9aVgnkOl0yjCkoZiL1w4FDj3L1w/AnonVE3
SN30cZ4VPjdBWYc4Egy3LqHjAWBR6zVa+GSDLg9U0w0W+mGak3x3pa9D+tvvPKPNmThtIP2u6CbV
SAjYaF19+c0Xq1AljgYyy8hR2bLosKEj5xbEtahhP0pCpEJN8h8emDI5JrJtbFJPJdAh7l9rFP2C
ETggTWvUPP2V0fNBiIGyM2oqJL6N+amQfoiDXvrgWr5JIHwLWxweXi98zARjx7sJbji6x9yWWVvs
Ohx9HJjxKq/vm+WmbrrMzgVEikWZY0rKeC/zSyS5JtWRg2qT1gjQaSBiF6ejXBz6SUQZgiHzySIL
W5bALC0K4Ah4JVEl8dvmWZW03EbTiaCpfCeG+KezNUCLgVMMAb6+GvuJrloD7nIKaZccY6t6FkoK
3T7kKD5VU2qjdKvuj4tQT5cKDim+lcEDa3C9GUUXUprqnbNL295BE0HaxT3krvGg3babqQEUP0wb
PbPWQP2OcydHxbsguOlCfA5FRXP5R+lQz+bNsBKwUQDIImWDhx8OEYYBaHkTtoDPMTD9I2MRbyUQ
X8AgH3FTCSoZq/FAW11ocZLbCwF/q+wHfS5xYsOP1Yk5CNMR++mgPIcx1Kedscmxm0ZU7Yt+ABoc
N1zjNBfeCvqVcJngYW38cCkLt25XxzV15mux1+9S3YqaYZdfEe5WjY7Mob1FSQO6+2CC2zec/RGY
yVaipCS8fXVGid+S5yM9Ar1YiflEOlDZnBWWHS0A+iDZVKoBed/4HDdLkCRWa8c01Krbdx+fHx20
6HsLOJknkUrLDGAW4qfCLm3hPFV9N4qyRoRm2cLHjrKuBpYVKuAgxjmIXBkoGIJlQrVKLdRqr1eY
r2KhD9VHnk7YC9hW0xVghF0Nbam9Z/Vuv4HUNCdpBFhZQviFJB+AjE+NLVPWKgDe8ovT+prVeMtc
rBtReW7ScXLrYaLLd/M53DGf8+rfisg9C4x4O1LFiMxbIcWTOYv+iju6Hb4dPMZUrECPVtES5Y+U
BAVln6UQhZtM8IW/x7rTp4D8hDGZjLO2juot3U9Ui716480PcHBAEDWIss4b+GoNaIujoFkgrfCj
06PHFstY4344+NUBT0GZTE8U+RkKioPyfoXE8PP2QQYLZ2ZTSnD17qExFgzehBbmknjsGsEDoIos
TkirNVYlHfyaUSivDKors+USNV7HdIlVM/dnZ9UHieOsoJ1rFxUiiVpJ2WE4BMPnSeg1RBQzUl7i
h/mOkQ7J6GZMeZKb/L9+/B5ek4eqjzLyO08fKr5Ka1w/KCpuko8NjRwfOdyA/qUfbrZTKKJcK5zt
odV4xHAdlqPrmJriGVvGE6ciEamChXB8pSzRjMeNTJsb1G2FLrkR8SYkzZ2PDOfOCRqhiJa3XhFI
UnIhtL2hfrdB3yndGmiN/zTej/fEbK3MgolbvQ6I/qFe6bi5qG5seKg8HnJpujc1tq7bRwSsPGz6
CgAWg8Onw/cHTocHihm+ju0WnjRzFDAHVtKb8O3T+xdIbOwIPoUjSZvA4S03hF2VmNgpMPgZrvJP
J4momGtrgShNpzZWuhwlzYGU1AvlvQvV+n0G6shPO04xmM3SDUaAwVxgKHp/fi9T1P0mO0H/y8cm
LlUhB+7xy7bwUYOH34Mt1+EZLy4QWB6u3IGkiQr8pnGOBSag7yx65fYnpIE8sildf+J9PBDNOQXS
kVUTvQhthM2UuJkB+ePDqiRK+gnvifal8NWmDMosodxgkU7QWYN2xC+GkYqD7ozBeye4x2A2kYbd
DMQCUMiCKCjj625Tdg0uDuIsNYVGwcdig+En3RmZYlRi8wSkAsYcv10AZlFWR9JHdhMtZ8PzW6Ll
eEcvU+iUIpZZsAhI9vPX4kKx9s0N84FKyCZTX+refWCPKV6gHT0697Gs63ZifoREmNAz0lk8Bep/
3XolssJd4grP4Oy4KkBPb2DAr+bk102R0w25HqWIcHhpLlE2KMjRdhFW5VDOW6PRQ/qtp9GAonNI
NbLG9Cgn/62dnwUcYNrVFIFVsADV2QNmhVMj7UvHqRJOotFQuhwAQz4uMBBzmLMJGuEzIUe5pF/9
5NdRGSmEE1CYOvXDGZNh8kcdTvN2PHHI2r0m8eABcYqQO5KSf+0X1mgLP2AXi6EMi2h/bSK7LAmo
lQQK4pvKs1L+YVP4TkzP22Jgll71YxNzE8nfcU3pipVBR8ioITJaKW4xRngq5iIdDZ4mBjmNh63I
S2Zlik2/PTmrltDtm2JIBhp7ovH+B5vD0hNUo+/yNwMEfTSnff6eSk6gszoY2JmhkFOSw4q1/qfK
DOSEXUZgN5fyjxPyDtKsbE/dFLAPDrpk8M/s6tH/ewdQ/ppIujXROTOCmtvyM2wDuRpSmEVqtEkj
uSozi3kBwl7FEZ2GOV9CBJ9JH5nA8/85HQI2/AcEvIArahi/SJk/FasHcRxYlbTkKo4bf9Ga4lxa
azzxTlV5E903k+owE4PoSRNw/VTOVy4lO77F70fPCQSFAE8s8smalk/9mBANtzXfC2Ea5/ESP+Ng
hbYiAxGWmO6fVov1ZY5vfePXvDidD3rrX6GMvpKro80fTDiBfZP/UXSXT7LWrTI8BwTib1hHxg/K
euXb81usTxtJFC5Tt7PP8oJdxE82pkZ1Pab4JIoQ+VbGDmKaZv0MpJULCvsGeuEVf8k7cVVFfqJS
89adCdhmOEU1pX/aQxUdcM3OqutQnITm3/AGnCGYG+29r090cb42hH7imqXXYhsTpiADFO30Cd84
2RsxniNoMjtg2dTCQ/KfAFhQLZYszL8AYvgAPTqAgK1BnCA8Ogu066WZ1gjzaEJaa12Tnbzq9bAG
VOwXLmNJUza/7hOFNHnkF3qS0NRqno7knPz+1o2GHL7zt3jw4jpGIsh2xTM+iTv5FhbayCzJNTvJ
ZR1YLSiKVS9ZFDkuEcjEi9rppYXquYMk7OX/IOYkN3+X1XNEI5Xra30wrTRwLbYuI4uhN7fkZj/a
gKFdoartPt3+72bUh3qngS/cCSwHZ50dSw+wyZRuFAK2PRNxGMte+zv54/E/e/p2PIHDP6amYuL6
rwFVgB98CXBX+9sc9af7RMk79QLgEW3PsxBDkqpNAcALpY01WKFA7tVyZDH0b2Lzjdwl0pDncciu
PvkR8QyE02Mfud3Poq+LRsm7eJ1tpsH4xLFx1u01m0EKq1cii/SFUwyMrCOTse9fWbfgReR+rZkl
TcCFTid47MpBp+wGdfb1xcM9COMrgtGFvBCPD8HNnmFWZ9Y7S9soIVr4AYt/O+/I3fVAWEQkaVzZ
DShcHP2TFzjS1hnsSg4WzdQHJqiL09TGhd8VkJp7TqkmbRBrLTNXdPA9eq53Pp/gwNVITcJEGY2N
AeqjadPDA2fZyTx9dZsLqfxgQChcFnxOBedrEgDt3ptXM6fy4mA1fjP0Dj3+v7ncafl7xId8QJgs
ooE3VDaHLRmeIOEWB+YQCABhgMkjKWtK77s+P1So+s9yckbW2xfZ6q1CktPjKlaBK5oPuw3uS5Ga
YfmpA2UvmdatYDGHo+KdQWDYI06ua2U/nsUXIDzQfl1khMf+Vi2HP4lpp7I+7KgutZ2hoJ6XCYCr
EvCNLRchY00l2Of+vDbl3v/+dAc/gVpupUmb6FIrG7HbZcCDoNYxkJydoHqg2sgdialXU97vOD6r
SMd3zZ3b5niaKDcKABRqqDSdFWUrVyKjekFIsgxYqmhSvehUFiBHYcnoadBi3NdL1o44noGjx/t0
6jxH2zQI/po3LAQTZuDtTFnfXEBa6OvrP3IM+1ka4rQSj3IrBIAmrcI2vfBIGks+CruAKJuIOq+u
xAzOY99tJ751zA3phsiyJVzZpiHGvVl7eUg9Dee/FwzNQCf0/Q2hboiuoQDRpPTj5JhrBC++miKg
XorP8MW5OwjDw7HEcOi/W2vK73NE0EYRQK2/pLiNt6dHd+avByVgk77Mh0QEwq0jarga9A8q21wS
SHww//AKGmprrA3uP6mbFTtnNU50y9a3TCsbdTD3WvOJapinI9uXdxou6VWQG6EDP/01lVMBbFsg
glvfJZbVd5cckLWZNGFkrrzsugDUQUSjfoWq1xR8qKoDiQGndfmqMok7/+/qgIVsmxN7p9MIqHEI
MUYAHstCDLdvWIfojd309/3mFveSri9JfdtFfPWnnwXWeQ56ZS8Bgwn6asNR5CyxV8ON7WbIVcGj
wgzUP9fF1Zq4HqfEZ5fWxdChMqBrImcg6J/uK1/Q7CUEKKqUdSlIDSVYLCs/kxjrMQVJWf0yKiKB
mAk18CByO2fXH9U0Ixxx9JuYt4xhldNFXLQnLSExaDXhrREYPbgeP9KlSNMlI8KGpLSvFCzH1Rft
q16X2WlohTekf2lvk9JxJnGHKCBODcFvmBaFyxnpqKMVLpX5la5RlNhUl6zuV0kxRjioesLAD/ac
9owHlLrFgF9Kys7a/87kLuY4md0uvZj2TjANFbRpo9XLB2Kp8oNy4R/FNFTJ8XwnOvWNGWpdZfkn
7Bu+S5wiGLAJ1cMa9tsAySg2Dpv6IAY8PVKkK31/mIny3p51B1mNAIyxiSOYIVCpwX4Z9/fmbaFt
5LhDYzgtQAEANqvZkz6t3vRQZ5yB4nupBOV37Dm89te3nZt8iJ4ZiP5/ey/UQHCecdXHPXjbGPwt
7O3wfzT6HXLuUx/zKxt5txT0jJZDGiTXHjF+X55UMlEHUODs6y5FPov3Xz/r/GBteSdR055C+lb/
WGNVg4sqI5H9uoRXaYELuiNPHh/z3gdnQlGlkHo7oKTVA6v7Ogq/bxflf464sMZ2LSJc2tEfqh3P
nLTkOYiHS2m/xsvCKiepkfVOlxxpbDs0F+m+JVmFLDMvI12/sh2yoeTu79DGYWngSCsMZ4Gb80T8
RL1+6cLAsczwAd+AYIgnUCLdlgH9pbjPMC7W56s1LZ2+IBp/GWc59WVC4YU53tejjM/NRDPkVnru
ehnlBr4FngVCN2+TDkPOHzQ/pzW9LMHPEgZypbRnnmuZtHmtvTOR30bYPshM6bry8riULf9ti7wT
aDkpOl7V5Vfu6/P9/432wZmkOrSu0xRCsAVC68RAGWLRj4jk/FTsyEFkaDWf3+RNHDghQs+mM2Dp
fW+C4jKHJNYECyzkVpvmRJPieoIZnQw8D+zcEI2QwUJGgzs3OQHOsjAZcUypC/rvkvby+gl43QpM
cs/oG3qLtwtRIv2S6bdhERmb9pagnReKbvafEaYFsZ7OHJKLoZz/27qbvmNDT1Lh6UvI3HiahYf8
AYhAqvFWx8GO6G9sVJ+XZtjU66w1mfm3dVYfsx5QfQeH3m8FduLsFticVO/yQvWSDiMNx71xL5ai
ADGk96yt22R1D7Yk9NBUiuJrD414fMP+fOgJ0BvrcHihFKiCGjlwJaTxrFLtmI+70AnIhzfFQLGd
cZRSEpMlQGor/BRs55yBiXY+yez6cUcLubPeE1Z6FeuPAa1zHQ7U4UbwzEx3ggZFOG/+LVqLjPv8
Six3daXpeyTQyUxHFncHHCMvUCAWwu+CW3X5Qz8SYo+lAgi7etYA1O74DA7LsTWCqkDIE+4Isv0Q
yZqwUoIaKmoRYnPSqdC3Nyzn8Wcxi9G9gF1MnzpThwod0qykqR4MW9TvhcAsamkCwf7I+EapkYdQ
ho8Xde5dTa9FUex/wrerfYVOdjC8GcDlk0/zRclY5F4Ht0xbXCjbWxgmNAXH8wu/+BbvuSWeA6gI
NchRGor67vYKjixONtTtsxvQ3lNIw3HalMmGZHVzOWr5gCiuwybz3YnierhMS+73otHeNHlhvtPB
0W3jv6KHRKE2XSu8Mr7j9NkBXZ5sSoMugvzE7nqEE+Ui4kBqVQH1wVbnidAqLdCy/+sbbgZmGemH
VvyuZenHWSGToXhuuDwtwmUgIQsPdXhQ78mZeI06+biIfYArmFfQs8KKpc9JTxrs8mvGIUwKURXP
AcAWmcy5NyHM3BiJVdhcmca1jteBtyA5GzL2OZAmCAq4xbJg9kQmAEvXTLemuJesNE+LAA/ak/fM
PAfVvg9K1zzK6qZTjTFs3HFsJi/FwiUkan2e/pErLuEq7utYjVDDd4FOTaEg4FLFCdfYQupvBrQR
UOI6NDoyZDakeULSrGj2R/RgLgvS5mmSRhaJOVWxIrTxR7ynSPiM/GSVn3bNaEkU943eDcIndZ+T
YwD4o3eNrnA9ZthLtJUJMvtg9+NiIMnRSrH0zdbi3xLUCgX4DRh7zyFa9IKcADW1PrJbBwNhppbL
MGWsRNTYSpYrcU4oZJPllc/++K+cTLsEnfp2407+gk80WG8BSM8WyIT5R7v8RslkglJu2CLmcIyk
cgScjo2/f4kwApuY/oK/Ns1Dir6Fc6M3mKGQcYbeLRFdx0D0xQU1v+L+t25TkgOS0318qKRcxVlq
WfU3f6llwdXjy7vkUBLJZmQ26tbDoGvKq0Afu6sUGaK9nez3ze0lL7BO0dmGr+nWQxHFmYisQJgz
5JcmVLZlYMxdeQV+4yFrl6bx5V8RbRrRqnGjseuB0sRetqoxCIO6xapAT5FmINQ7h9WobkKPDv2b
WbSbwRIxoNw/+q8+AUvw3gSZMZuZl8nLj1aIIOjwOYYAAiECPQ+ot8PY5CMyDL7HWz5hVaCIa5eg
tEP9lmeeUsJJzQFfxVAwxs85+BDE/UEyzJe4Qm5GpKs450hZp0clr+K1CnTNzp0GEAjLSM0USmhf
0rontLfoXMRkjJK59ecFlPiiRQl9gPAGwNvn+lIkvJsX664O0P4lgL+I5zHIouJKcgMB8kRY6oaA
p0Uwl2WaKLEVaXsetkX0p3BHpDxZhD/GTcHrdSJek8d23gIUcfiU7+PZeRYiH3HM994CSVO4+Omq
2HIVyJRuvDDjw3qR4ElmgpImrrGpteUf8ZoY3Y7tcUSxwHtBllwESk2FDOb9Ufn6ay7488m+eHYQ
P1mqJrbT1C0ttLW6WcBL9VY9mmpNMYcSVdI/2PataHN9vsPEcdVx2IQnxRu956Wx1tO3N1dZ+2ZQ
hKjiYlVwD+xN22AAO0iQZjumZ8hFrEky09/FjoMB3DuJMU6DeB1OPw3EScLY99Fo3uOm3+GX8dhq
4YOvU5u2T2URiKKaILvH+EdXZF/dTUibAon9s849xBlQv7BGqHyFYK+h6KsaqlN+XzDWpNg3HcnB
r/dAr6NfMU2Ji2huCfwcMovd7AKYpC9OWe4sGDIeOr+w5e/MnfbcfnU/mLWcnZE6vFuJah38WUgP
a9M0oin+If1KE++Q+tIzzRhSWKreVrvVCja1dhY/TecTUwUEyY+aitn3sjFJNy2THD57F4NXZNRh
6YBwQlqONuLwz7inyw4fA2uRRwwLwuHjBoRorkNp30ihRfISOU0r/AeTvw1dRL42aqPBqt9VETbl
t9CbbN/GkIq+BLsot9PSBfaBYhILYXuACDDULB0Ahuna4RY2oyHF09CGqxitUnWbCS0iuVgmA1FG
MDgI+oDiDUYofY4Fif4PjZKa49hPzIrBy+Egp3CP2oa4sf/DWDv64Yt/bjE+j/SY2cq7ilecEJLS
H3f1SIX4MBG+4tHshbU4hwUH/LMYahPSHaEetEct+m0iDZn1JfQ+WlOh8+OUTqIHxDHysvbKy/+j
R+IZfcY1Bw0YgdY1wtmzmjuDRuXkDfqws6U7gQEdm4Msfh11s86B+UoA1FJN/gzt8l3M+gxNy1+e
c66MDsJ/aOFnymbKcRe1Fu1L9N4P9VWbWkkA20fujWPTpcpjjttB9vNyspFWwKV3s6jven1TpFQ1
eHDsX8BmCJWAzXTY5OZNLsP5lDBo+/lh9nePf5AIXIZY/QCs3X5jBlz7JPPr1gH498rspc007poD
FeNdgp1lkBNx6XWPpVZQGwBzbbpMwdgzux6cBl59yAz2qasRYY3ggxTcEfxTJWGc59Jbz24MTpX7
frlwLgTiPXM/5JJ1o0yxmMcTvqCf0irr0IK2dFefNHFwTWSrG1WHZUOHXMe2MfDBXcht6uRTUuHM
fiqMTr3VqyohBI2sXPU5SFHhd/BwALAM2/jfyI7MwqxVwffCB0TzwhtAEsWv3+2hV8xqQwJolLcd
apwfQau+09eiyCSHp1KLkGg8yHstJZwIXmeEFvjf1Th35uONvFxMfUHKKlg39P+BioAinyjblZPA
CaWzT7yzBoK+YqxiAfqHQcLGKGlgnFK4a4doc12t/TbSXfD4hQa5ZiSSVLbhiR/Sur6aY01PpOs3
vxN7+p9TBVZf+AiYIfK9vVNToNCMv43txyCjzxNSxs9QdYe55yGtaY/cdb8TY6klvJH5xuDSfjOd
gprWLq5Gn3xWX/htGXgmF6ATCm6z5kr3kUmcPpEDC6bWLLEuS8y216p6n/pgk1u+Ze6RRx0=
`protect end_protected
