`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ht9xCRtn+QHdfbx7otbuN18Dtjv6vWbRn1vSmQAMFh5nfOFjLk8JrB6tW/Te4iZMoH0QBIOsD4qd
VBlklaC5JQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DIENKgN0Sqku++0Jjt0w6pmu/lI/r/xapEqkEQ05H6objvgXO+HoQDEpXemxbpIkn9tipXHbW/2b
nqKap3pvqXw760s1kzUACv8cEpeF9GFynZl0+nf+O1PzrC1dX9k+lvEWM7bJU3tCsjAdyuDN7Px1
Vd5kuWEHUxIxPzc9T8Y=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RJWxbT5JmFnrkgFRdvO+wJOOsGYZrznBB+KiCdIHt/XRTIgPx5Gn8gaR925APTU1SIU3SaqcKkzX
Q07x0e2HOXH8jdIHRDOhtDpFA9LhAzv7sMN3HdVeiYFb5mo8bmLYrKlePGeqrUA4cbZ0r1457iuc
ATI9klBjxXQRtDZYfSY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ldyF01LE/dj5Jj07Vw4Hy9JYkwmo2irSintksruyhUK41mutswkJzJjZOqBiAfemn0+ew+YfMcGd
W++e9MrctBPTtIe3LMfanugRUtZJiy9GwDAbvG5cifGJyMqWWALBeh7Iy2HjqWF4XlJElJ9BWW45
3+hPTc2PSV/cENrjv279Qq1ejpPZfq7CoxnXvd6xEk8330aNfw8dPDFODUhUqvTZHUXLugmSta0r
3pf7G0oBNjDptwGroGMxZ/5IWlDf+ihmafUemDJomBFkAOjtTci7fpC+fklmXmHRBWAk9GhQo5No
EISiLWrvTnK8k8ZYb2YfkGBDvo8oSqDFMPnyLw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ldUyeKjaMPlr62HbfKoDQIKLUpbX25SkbceYdSWHmbC+qQJt1ljuvyKPiEHsxKKysLUi4OfNHtMV
8rxGjZcC7RzUKwjXn0UjzN37XT1v1De/OQhZIcbSsM+9ubVN7NwzAsE/5/eiaw/acSpoVu1UG1WU
KE4sHOGF54YAjS3VUkGMARy8Fh7Nh3qXihX7NIGG2X75pFcSfrJ68epQ9vPtYGEsVr/SqB9kGZOv
EcDbIi4vpTx1tVtoLzteohznpwOPsuZlUGvbLht/xjSDnkPtDaTc0NWa4U3LPL9DC4CCr+zHQ6mY
S3LtTSz7mc1CgyXWkAgMjEEbhd4kB3u7RwYxfQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SDeiPdGRq847qkRmJKcp4ibRGBmK94d3MB6PDja3zsw/hA6deMGLanb1I5uycH11VwUwJRX+N95+
+AQ3aRsXBtIeiXNw7XBowtBivuaUQoEqJSINWsBBcY9mP599PNHZ4x5ENCmHjHIut4PVSOnb6+eY
h2EtyYD5weeMw+gLr0sgeDvaAJS8n8B2nhOqC3jkS3xUAB/3FSxZ8FCKFBxJb703zCnIyuKgvcw0
l3W/PFtmNBNKDHmVqij4F5WLXqYr9yHJniMMKotgaedhDnSgFmMBv4opZ9GGEdPUiD3VSlEksruF
UI3Fsh4GZ4XVSIfh+c81XElXEgYHtoQeo+8TFg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57632)
`protect data_block
THo5OTsLGi9818EuldVrSLsTdNcYFEcDzA4WhLKj4+LjMOrkeJES/Ucl1/7RCGcN9bap0fT/19Gs
tandkGiX/LkHBIoyNuy1PKai+qUegUfVMP0NJlykGVveBHoLhpVH8unZoHPmdvkbI/i800x4uMWC
uh+qJijMt/uimBwuQtB3fA4bN9QijPyALXcb4xQaHKRjnWB3vEEFlN4nSyek97RQrm+dYs/KZSEM
Ph1FxxMHzl7b+9I2Z8Ha7ky9H+7UHb7ReHH7uJ55NRVjdqUIfT+vM7n8C6GntyZbU0B8DA377lqo
6XFmbTjilavRnVADWioUp3AgkJw3y1fmXQeBihEpwhbuh+uJspZvcW05McjysDemTEEnNcIikHid
jIuov6BaTlFvexbwQ4WwOsOSexxSH+suDdXEMChtnwGlLxnte2kkZjmZNbLZXF7sJIQN4jPt2UO3
onWwoNTfGID+0xau3slvtRDsk0Jz2bUI8nIhdN/xIK1Zyy28QvPaYkXPv8q2yLTcRCeXVVJ5o2dw
5K36MbGMXeQCfH2rMrVoP7jXQf12Z1aG8rzWVh56WR9vetJ+zjpc//w8ZEIJBsJhoQCFKey++eUU
y6nx8zI1Stj0uZq8tiq7GF8FrC5Va5eDd2yHd1tjuO6LENNcQTJI0NMSihcKuofazwoTEcZkpY4r
Hu5aZH9329USS7q2FBK+zF65Pg22Nt4cMqOwOXIgbTpEzqONlTbWtvOsyqbdH+luqLioBHTFMewt
oY/37UpKQ74PakIz4bbcC13vBr73CuWkatKqlpHF+Tb5cYj8dRiLr4l/nM7CL7GMoKtzDx4tGUso
+/owKAodYZ0UPP6S+VG5R/qrJpPzRW3Q3fjvejbs/4vCMGEFRE6B/flilk0KHS3Zf2w4aLLDjjUV
B/tJVVDPCo4anupRNkCgmlp70R3PHzLcBygUTPKJqejGklIQqG4xTn7Yd/fMzbb5NpotpfSb/QcE
pMIdxgiWj45leIjM+1jHD6TIpNFX3GmRHwDsBzW5eeSITydjOjJX8la1y8B14ppEWsoIdic9soBU
RBbvCtm5QfHV/LI9NB5YlLfPAQAsBpJPI5jLab10TXCJvF1C5ku74RT+NIOsd0e8aN5sDaxgrenO
bH0/u2Yy0/PLHtxQU6AQP52M4oNJIB8z7F/OvQ3bi4uKogH5/BOpmJghfXGUuctpfY3OnVhL+Yyk
29F340MK3z2xirbU8Nmln+lOfDT2SlS9YtEgV1EI3jhXbO4+NiPtp8bp6Ly4QnjE0xBR8kg4So3H
lQFeShD9f0JSvslwG6PshNGpyRmLu7qrJBI4daA1DZkNFNwy8Ymu4IAgsmZl9PU3m2NcaxidZQBh
J8XV7ZVifOhSg36rGjHAR2fFAY9P1BPG4Sn/ecKHmydggxg3bNeQQQ39vodoeAJwITmWq/j01zpz
rW+V+fBkRqHwSbURdqAtfC4e4buhlqzHK4YNZyXSMfZO3KUoUAHvkoRjiT7f15Csj5PAeVNOdSz+
eI+MKjuNpqderXLBJPBrszD+zTxkXh9foY6tQBOIiLK1VdleJRbc4TNp20/tq1t+bqDtoy+H17Lf
xTHtI+EqglNbXgWZRpEBeI86TyptwIaK7E8T8Z+VoKKHidYGFwGOVrQCu9jrfLdMQXkqDAkCn+GH
hcnH++GE/+Dz/iR1tbWIFq0C7OxCLrLCDpO72+2uiOvKU50KwxSj+Zxu+4bwEpLMxPORKmNK47Er
1De7XMVeXv5K0gYb0bOxF1LZ1dBxbnhpfXkdYd1NJSywT3r14SzUg8QU/NBhx5sulSE3bGOMnQvT
DfEhq1P+6+cOMgxD42AmLSEBrs3LUBirTGfmLqk1xxwrjimUAUU2uDCT/V31FBTUsSRsgh3PYHQ7
EzEvjPN7vD1tEhMvORKCf5s++g6D6UWp3dE14rb72LhVf9hUCBNbOXNEAtAw0mFEfpl2YQQVuE8M
m1ZC24B7WSjrD8JqlsiezSf82JXQPuY39Irqd+eOyuR3k2glRb4hJgBW7/R0r2MIpWVfnW+ayoTF
e8E5Q54o3md252vEd0zkmCjEjXZcj7bMNAJPNiYFYZ2pTs/CVf1mdIMIgvelds/WChkSILDFc/sq
mBrYagCStj3iWfhyM4sMghKrKDPGEiB6gXNGz/QR7Nhda7MFOk+G5VU0mu1zGqtmSvvZUgqocrIG
ck4c+bQeW/6I+TK+nuAWKLvgsNalMNZvIp5LM/SyM12A3XyuHhAyt9Ags37TFASIgqZDNpbDuxy9
jJ/S5OBZE+poltesckkc+YUIcbABS63D9BuEZOwGtoukpqlxiL2IGw38fuYefi2Cn6B+njLYz8zC
V2aGPRzRiX1ngMpFLGX0eDMgM9XSMx4OVibVkwVFuEwtf9qE0K9crCnonmuE/dWxF6mAMEnkYDfb
y9ANqKyv/sa9F1P2hH/1EoGGegYP6wsIelb53kt82SC0ZcNa06KjVT27ZMz/bPIPtOvPYhtY4a1W
o5khAuVM/KfCwm4ftlGHDTneIa17L9K6OWNgaBEyPRzo7s7gvbAnWAAsvgQEzqcP50c+YiBwEiZh
CI97UnGb6PkHh94esF5wGtFfxduNOJdjvvGwWmkL9p4isBRev2oWBy/qAhPCzCGmexx3NPd6isrB
mu9RD0+R7v5H9VWui0LFZU8nWPe2VDUzyxuegFEYTkc/GTFYE/7KuqLlmQGUhiUh3aOOE8ohyi+r
o+r1Q6KZJENV1K0F9rqsD0j76NDYWACQkxoBWQK1QdzCfofp+/0TQQ4Wh8DeYvRfzI+GQdjRlwCq
Gz8gEFIfGckcsYzTvV91ldfJYIkSmOHteZZuxYYUJhBEt4lr7alBc6/XtrjxPF5O8cbKZ4mFxQie
jU4Q6+CfsPEEODj3Y75ZGw8xSBtF9uAgb6tUfWIzw2MjWUdS/0W6Xu3mhkP0TYr16rbZlRkg3vS5
5oEu4PmjMJrwcCFFpc3+jZUo08kJ+sieQhJclREPfgb6Pgt2OYldXaziqNyPau8FPI7I2taWSF6L
YD4nemx/yINEvU9FMf3oZ7XANNdC+2JvZs1wGUbA0D2bLY3/5oBqguiwY1HX+Tw1qrIyLAHoSPJX
epl8JmgS1dkEMWjN/9bVk95aIJTdaFTdQQcwN0YasC69J1pk8gMCL2b2ygGbG1t0pwqF5ttgfwZq
/fLwoPCxIgT53ZsXYYq+V39u2em+xHeJvG2qhacDcQaNIlgHSax37dXUixNennxULZ0VdDz6cSL2
HABY2+ZK9ACxavwUb4NBgLNwvjK51nppuzBhcnfy/hB1IpFKAAhizOw4JZGtbMuHeKfOtmB0D0tJ
P5UW4UZrvbRnstMSqaoyja4QvEmauH+QsfZvlHuoia14vfQbRynVHMxQDyXZgMNSWefpvKX1hdB/
AC6Oki0lD3YpzhpLCm+6DnwjLXAzYNDgBBtKZmEJjqKTtj2uJUYRkaOnaENo7GHdBTD2jIy4VBTz
1trFlWsGqevuZmOCErClGxvgWGwojrr4NmMzx6BEeXnKZJmOoygCLqV6EMjqO5MgMD39TfkOhWS0
9OiMGfHGdBmg7aoID9EO1vkVk966IOJVriULPOMs7nAoN1gMeIXqPGJKR0uhJ36jPi+SkdIL45Wi
dqlKdLZXmK5ttppWUjOJfLjRrxSGIeRtwopQvROXXOMRsaoCysOcaW7wo8pxKMiA4zU3sepnVkIy
F3DnPsU7yqwTXPuasHSk77t/s+y1zIJscmQHJaF1Xj8aimQYB1PxfnHieyNYgsVXUQSiDH2qNm8s
HsQMaaCl17GxBTqzcoxcTiPyP3RPwYe6krm58a/aaZxJxQR00wRni9nI0bFR4h8WINDOclAo9WPJ
Ke0HX5yBwqG2UXnbXWRmF2eXdl7npUBZAFrENbVie96uTlUm5tCBK18QhSYaw201An8CSg/uJd4J
sZzR92tm0OyXeWxyOhrb7lx5O7EYAMAbYua+mchN51f6HEQQaso0U2VQv50Y+lAonOo27yHl2f4B
XD6ca1p2dOhiSuaYyMn8WY2dz87fPG52+52w+1jbIUFrY8kEyBL0EgviTgiGUFjP5eBaWkdaOXLy
RYH/HG/fGuuGHWCqi8R7AIj4SSoWI6OEp67divL3n0dmWIGfCebc6oHCvtDg0EQCF0DGhu4SY5fK
I4vqAjSoPRiFCcbJWSAtpqMj/k2XpGxc69V1eOe1airNWzQb7XmJKarmkGLX3q67N5rdw5EKFgpO
vd2ZQjlUl6CAn9Z3fPjC1UZDpPbJBUz1l34JK+T3A5wa9OHJqNczgHUfzZaidB0Gx4zsHgPqDC/e
WBBYvHTdTqXNIvfbaOuGhZpVLNUTwoSt/iq3F6wGSGCpC8krfUGYXePM9kUb3AWvn1ldlIvf2q9e
ZcQgE5SE7JRRggube31bGC3+tMW5p1x5KpmJwCKUldcH4cs8YxxqyfdutDOiu1ixBPihGa10G1Dc
CIoOaFkc8oo6iXbrGGudF5z2/y2iqVRed1ibH68M/53qYEN3WvtX7+5A+DaPsjSDgQFDnla/z6Cm
xYD7R1U20mWs7fgl9NHjALHe2gFsed2jJO0yl3z39YG92awFogelwRPCKrePhX3YKm63OddWtG3Z
ToqhZrJQElbQWmJscBgMoMozevuVZ0hiNIDpjVXso7hvicyBXIlqK+pZKHJw9bM+XEOJx8kUtG4/
RayyThkgPYUOY3PPXc356dalklXGuoiH40jxkcuPDlSkSPJQqdhfQbvFLlswfXGq2FaSltqhE/wY
xkVNU3YJCVjPNn6hnWquqbjVy0qtE6XbeGGjPiq41oq6Aip8CUw3HzShEmtvpp7wPT+M2l6eu5Tg
jmdtrZ7gVgJWJMXDYzZdqxsg54LTXCUT2GPziowgpsTg7wFdiX2Dz3EHYfAvp4HkhjgmPz1BzRY+
PU8qol7q/+vLVZh0e6pWwIzjgHBY3KXWC7MWWS50gUB9CkC1VXSP6zSlSvPE7tR4oD71SG6Oib/o
FYjcktoLdwoI/iBWfkPfOMBHGJ0aaJRUZZZUIKTUGsFa65ftaejisjfjxlssX4OTTmQG9Sb9yY/2
GY6nC3d/E58DPjYL5imAuPKs4QYSLmtKN4c2CFMaJQ4VleozJdguVlbu0w/uEqouqPFUgSnv26dm
l4floRUiEyM8qjswUe0uTJ/loMQx9OG8N/rQbXUBuMbGxPhPN90PYI2npqGvnwvNk6B3NnvXbYYV
Irau5UpQxO8pc0JMH1W5p4NVvJuJ/8WmAs/1V29GB8vNs5pGvtkDGpEdvg4CmVVI/BeUBk075iok
kd1XXIJRNa/PF9BqrW6NOUvPJZ9pbob8SQJXfSRUjbjeCyAxe16CBhRjbQ5drweFqXJWRibBT9pj
SzgyITIYCOGmldTKig4Miews+Qh/B1b8c7K3rvp6BdKaTP4xkXQ1MkITNaNHNqct7gXwC/t4jL5c
/a2DJ5OCdt5l/NUPoZr8HmqxqN5+uy+weWer+yuPV9xmwJwC6Z4+pfCV9unvmt8dYoGqMI+4aMB8
HRlBxpm7egCAwIrkGqKL0TntexZ7L1QVvy0C5VMyPvEERpkL9bhQrl9oD4nu5LdTrpkX3ZbqBbb+
2bfrWPRZXp/jlRUwjeSPEnPHF3ct70rxDYgpuYHJ1lTVVzTonkVZ/mHL0YMNJxj4c9aB3hrFbXK1
7orEcBjSCW2PJtHhcdADNfC79PDLSAKQkg3fa7DaFyArbEFbGq/pn+aYBgr5asvrtKPiktcsdAzV
aCkETdnvAJQ1+486LLzknX1Q4luNuCCMmZLdd+GzRJ7IalzD6+j8jcyj3eTEY6nC9qgAC/e6QE5i
3Vga5lkocuLeurHjCMpDMTYh8X1J+0kSccO7kaWZTggjbdfzssU04lp4jREpoEgvUpu8mU6MwIVi
iR2OSDctqOEjwNMzpWimU67SeLs41We0QOpYMg4h63oJL+CBPc32Rsh9f9C20faA23SMznCVLvfZ
Ze3ouH5YYMBeLzw68jHAeEVDn3TLZXxU1qUBWzJf1KI0txYXTFrbhS1hzOKKsEcXvk1ox/mp3/MS
sDfK6wkunkB4cHAvlJP4jHvusVXHmFNp585BMI6NXSCA1X8/weeBsdxebSMom41aXmEe+DUpOSBf
pPSnIUwBpER4ZD5MRcxQaZ5DexktTrdwHTv4CRaQfspLTyxysUvAGyVUTNU4REzteh5OmvtCXE2o
NBrOeZZb4vuDyisghaCqwY8ltVy3emUnYAGhjW3zH1zk5lYBESMbOx14u6VZJDWbv1Q87Bl9apFK
4l5oTP8xR64IikL1IkAwoSxe4z27ada0AF3cMNBQUvKC2Icztn8a+N1XXV4VmLRl+ZldW/DQQR7y
uUeXiPpH4Gi/ZZBHNXoUvyxaA1rBbhvfuxWO+ct9P2OkX3pJ2lXqrPbmL7OeO6D81gSGRoQo2mmQ
xZznGde/n3axsFCQJbLz3mQz4uSCaOMQcDXemivTfoURVobWtude6N6KBGf+Aq98v1rRYdn/BDGO
z5eREFgTEsL8eY6JFFq1+gMyiyUcgPoOqdOfNBUkb54JpIVJYD+y+YRU+ZzPAPhyJ8PAnMlOkw27
cZae3sbFOecSGUq9tBwh71ypZvUkj5slD3JHxvoS6gPHInVoOV+6tGi05HAlosXYG33czPaAJ92m
xvmxt9pfoQK20carlyLHCfvLP3451YNQ0TCjT9HcXqdo1XMS052jIqKs+3AQTp2yXXXK5kRTVERm
iQ3yjK3FSkYVr+D/rYuWsiGh1U5ZajhpcGiZlufYIfyDFty7KnCdZRDGe1GilsB0XWCBDDjXE/Ku
5K2bGT/O9lF/+N3wRFUGI37RRXwcroGkHTMDaDEc3KM56/00suhtJ6p/Jb9D53WHrBvAeyYOB4S4
q8OXRcyLwEXFN99njJX9rAo4tun+vCU8aUVx6l877NKG/QtZXtWzJwBgaC+d/hf110QvNTX1vMNd
QkJQqNwhfNvzErP3bJFwxwPWQmUYw+w6/x8z+VHMQ1zKnk4TNGI0c0suxgafcK/YWTo9czc4SAez
Oifd7SxYV9vIK0/S5NPriP0Zf2o4cy4y64BYe8kvqCraY6WcVODl+IDCw8hHNburKcUDu9VeJ8Zg
g2yi/CFOVResdVf5c4fmdEVHt1eimYpMLUWKWoJAcfdq8GDklz02TUeeDCuTTBabk51/b6ZKJih9
+MMRD6S2kibn+JCJZvLn3k9yVvTB0MHhG8kTfqFhbL7hgm6Zsqe6dqC3ds5WvtgZQnBXVA7XONvp
7QeszE3c61sqxvt9WhMv6b38WgduYshLLL8Lw47RAB8tGHChBaYgYuc9ohMR5rswXYkgOiY/f63v
A6UtzvNiPI72EfVTvqGDPGET/64zVAV7c+GZK/xspkDel2Q1tQPW2XgyYK5i2etJYyNaJsayYweO
tqXr5k6WewAtb+uX7l8KIL/xJPSWad1WTx0qNYPJfSGfQjd39zYQYv+t9zyDFPvMO5l/7IjCfxsP
6YKgGP9RjjOupwwyuMdP+A4pubp8v5zjLN6sKfh1bXL6J5rggLZmkIylQ5swqx3DO2vHsl0Bk0xG
WHXhZuhO8ktFO8UfH2qTsplR85ueO5D6r0BS4EEfTA50NqiAA518gKDWnkp3kMMDQk9Zw9jasMFn
3JSJL5LERynvPryLmh0goSyh0QeJ6N87DzQoU/UHGadIjdUtmIt1tzLZn7IzpN685dRa1cDlu+TG
pOsiQwI1gqZ8GopWfJyHp3HhvNBTkvpUrro1iiW4y6ZfB7R3Cy6S2Ekq8+/kER+7ikbVo5f5lOEi
wt4uLD/ANqGNrkjgwgBRWojWzVswhFO2nf7CFkcKETkTh+GHmXhJ59j3XvZhgYBeNaA7SBJhU1m+
eNUyleA9WuYwpPjAN9VYw5PRS7fGpgGK0mkCEx4eaAgC3LezsqohIIhbKkGCxYUNyOpSOr6F6MNO
Dtlmkei1VpJ8Pre4FX6SaoEBlETUe3NdfEaBL0SgYT1y8o2MnVi1otTVPlQGecbbPVHxJpth0qDw
jpsUOUq17v3m8+dmksAGndLWoxzmCgVLMeyiH/BQEHk84T07rawR0YgPqXGEi3ENlv823qD1pa8E
PscJYKsVSSO+KGvo4i8YU61ha17+v1liwi7pG25hrPgViwFJLAoYq6Af54Jw1cWnUvbRZ5sh9PSr
nOd0wmQoDn4OLChSXySnayLLzosJ+Hfd0pQlNdu8WsK7tkvRN4GDy2MJz8wWf5+hV4QjzRGhnDm0
kUC6xNQPSaQ6Y1/TCpGc7dsa38k3m8T7HzlQ4Dm0+2XVrYvNxtts0ONSWpZqY1PI9RJb96aP/+L0
cXdxh4Yj8Zd+Qm3YVtDRhTn74D2V8EiTAxkX0EM70hnF2k5M4rJBW0VRePJzIscW1KlR0cT4FAKm
vnxTrS+HheDRoEO7xlhhYTEAuF+uIsp+nD9r9JUUyDIIiBWvXxWuoXesoC3hjae5gXzCko3mUdZX
36FZH8Kkhajb29Hj9o/fFEtiyIg7H4bfO4SPPB+mQlztAtA3VqZd//14mAqUnsFnwQfDlRSdXZAV
fQr8OUXzYPPuB20YTRwoHDR4eRZJbi1pHlRxkSVPMHrshHtPlC9OcXvonJpvxPSLctftRAw4xZlm
Dk/lSxhGv8OEo5W77sw0I8VJmNEgsQ2di2saIQ//wzcmzuNmH3G54xAi8bvmXqycgyAm2Ho6bqBQ
BlXqziaYLRVR59MG2jnP1DYHvE3qsAHR+WdhLkQdqFCTFa3CTlmTQmeEZ9CXQBojyM+jrG0jhPVn
yO0j7TvepKutBo3gHiYMidM2skB1BzdKoD4ou2IlvzFmS4SecX7Hcl/G8tYryGYQkKWDRZoqCzeL
RRWaivBLmIwQ086tuhj0jjx0LTRYrzJMePSUQFV6emq3ePffuizO9Rz9Oa3qLsbJUe7ep1CXgw6i
J61PwE3vb0N1WJFz48RNznWOT7TtHU8nbReYcATNCgZQU6SzyG9hlWXWc3YZJR5k4dsLWXnnDo3J
0p1t/eJ94ZsnmPthnP4ggfsm58qpCTK5LgvIHSf4ROOZSWzHsi9UV40EudXVZt/PSsMs0qCMEGUy
HuHXgHNH6Q4HXjK4ARbxESNAGmTTzppb0vG6VehsSoyKhw3m1EhQbgKEeXPoWu4jq1MY8qG1cLgx
dUbZA95heLOu43T2f08JgfJ7yUiCPJpEK1o70sqkRWUXzQC2tAmbNcIs+y7AvtyVkk38i9gOgOXa
Y3jnh3HFF+/L6VXY1xoW0PifdqLiRe3vAoMP5J/IOterDsMfG4Gt2GwMdxICYh2XCRMd70RQuGYM
hfiffKGYtdK8j3WOvwp06d+dnioaOXLVXfn+ZEATfJ7yKGKXZdTIYGe4Cx6TBW0zZV1itTqYicRA
I81Q3bCIJ9gu1lCNFeQORs43/8s0U0S+onNaZGKG6nfJ99fNeZocHIFCQ1pIA3H3RIYXkUf1f/D7
5J7qmq6XeUj4qF8KKaUVGji8RxeU4YDqeO0EJ53jxy7G5ayCV8xcAU6zya452/vfG5DXfM01ss+f
Q5eJEI/j1Su3TGq07p9GvVzpWtRjviwbA0GVR6ZgpNkouILp6tT1y5JxihEyBqC8WiqAra6WH2LK
iDcBSBQGkbymmvSq+uHLQPPjOlI0VlZWCpwoG45qwHsmIGJMN12PGOjZrJPOydSwMIuQUo2RyA4e
M3auk2+CmSs08NvLKtIyZQZnY0cEv9dDk98GUw6BEHpUHhm3mYbnKLF2p4Rhycn8B4AaX4HZ47Hz
niDlEamjgUwdIEEF7skG62sAH7phfbmkb7WbVyp3QR0NTsFdlLZF1V5Y40slCP26paN256RnIzN6
uDmGBBEsLvvKuagkg8t8iPLHBScBjL6m8eLuTHD/il2FhQfhRZo8wKzcFyRgVxAv/PSda1fvmtfw
agGmmUNfpiXNuvUtSE7ay7HUZiFSKmKrn4DNUQbiH1lpZp7JfhuB/vASKT7qZu/wn+xf2mUqdaN/
Gvvgj4h4TdvzDAXdvPnVmfUIZYg2JFHrmr8G2Iv9I7RPcgtaD4a8TdmgUmOMuj9Mt3mM1zjJZimv
wlM0+xGrdnEoXL0vE111/HY5V3eRiSQLtrGUzfVxf0xHRo8og1RFHH1RXadqYegoPnCFNln0jV9d
/QDziT02tIOY6mRVOx+i3bCNWr84oKd+B9kK6lkdCiE26yumTTSg26glOVGW3+hrbySoEZi7ggY5
xFzQnKR5UxDOR7zldgPdHqmdsOKlcTOppdh21aosFHD3dGYER6bmSeYY+u+kGbnHPiakolTXQP/+
aKlBOMxyM5hlQJS2wEc5lXGvINFa/pquC75LzIqifRDFC6V1IJqPuKrb7iaGhp/uSCpdbwUl/XbH
FpyNcsqmvfwlj9c8dJWsZPH95fwoa3CCMNO+vcjdjgrWm8DaPYfHRGZ9JCdMVr46urChZkutXJC4
3yszUFlmyBxj+G2IOT3MsmAJvADtfJMo8nBFBaebhOeP6iWa6Uxlr6DEYh3B5BTu6IhCWXHCR2BE
DDs7Rno1k9JytqdN/4fulPsyGYSjicFZFbty6v2JXJXgdn3o+1oIFIGeSR2sw4/9GCJCNJ7hrlsx
mW8+12sWR57WVsiXWHJ8qByk3kjn+6SV3lrIe9GzvwteLjK02L2trNRtO9k2336XtsJ7KzigLyzz
rmUsQUEELZT9ZsAXX1+z4KUmpZxqPmEarEi0Jt+bNatWelWqLY1v+gu7BBl7Ny7PM1UK/sxrn1dO
DRLZ+o+AFJfutgl2U+6AWGc3F89mGQdEST5F4zMgG+YwcO251OOCphvCT0FFvDKKbVDYUQDYa433
jkBUQdwMavlTl8q1Ys8F+E+ixVs3wxQ7/TzX9mP/JhjxvzUj9p5EdKjJAuyQ/TR4SmtkKGGYP18k
upnEhVUC9FKK/3ZCD+YLyt7h13GTaheWj0dxqgBusCbEEs/LRvL/4NXR0edPA6+K+bME6Sa43uLh
66WbfBRir1H280rpKRIxHSmF7WC1wbXqxzlaXpsLgs1vvbwk4dQYTBcxI2RQrOiyUO1cYr8EReSf
u5iY6ark4y1Tr7Zohd2nukitDWGT4hIS6EdIzVLNZXcWQTaiEthqxcWcM8tc3xW+52v88qB2hNSq
iPeAdmkgASYcC6klktTUwt39iE2jNAYBCX+mwY8ZmoO3sChUZ2ipmM1WJWfBJfRqjo1LTlblxBdR
AjmkuHhSqkRkTehRMMO8r3cm7MLwgyTlZILtq0g4DYZz1ZhMHeWrb5Ly4xVo+swwY28sMM0KHyK5
INhVv5FtEwrxi0ArHlY6Z4wabnyw2a4SgZAM/dX/xBcQx8ducAUROpy0nSJnvHzguYdy02o5c++w
EWEMIgQ17xKCRqzmM8Em1i5fTZytCMlvY3Gq7p/2ANIjE1tGe9PCUhAt45V2a9nx7xSxtwK7bUB2
mfTRU3jUeaz7sR+pfUTbz93XGDh/NLyFj7VTV9I6tDUyabHGUkZvmjyLWq280haHxzJP6d+4jx2u
32kxWlhBGZ7nWRy6zgEp8xIO/u9wDw1FWYNGz8m9Z4aWNFNcfN4p1Efkpj1Dr8ihvFbQKpJxuwPQ
MycF24PP1pcaxQLqm6tL4F8yHf6GYUKV1VqmMaLsg2wHmiwOAjhpXRWCN9edT0FbnBKYJCkyx/NX
WnojQxdyQVoGXOts8x0U9CjBnzXOE6PD5a3fktmCjZJvd4P+AEOp3jovkYu8sVtd/noKNZaGlbpL
wtAATH4rmMV+M9LpnoaZE0kyfwMD+lbALCC9OEau6QEFPa/MYNmwpV80Vb6+U+WbCikEkruRZ4em
sIEEeD/eoxMzwL7Pi5w8XZ5thNNsAZAacL976SjZ2vZMUv+rtAlQwm1LHm4XEhuTZRHqRE7P9O0K
3BhgBiz+XXEDdN6uV61lafBeOtRAL885IB47lznyPHXNlnN0A3dsdMVEwZv7e/gZTfcLyfFwT1HD
73pfgRCmuC/U4LZla1XP/MwcKiEu52cWuEPZbC/AKd6B/r4KaXL47EqBJb+KHOiWhMMH8k95HL/Z
kPe8Y+jomxbcUoM+mDhg35Xb2R0alBM6NZvLXkvnOdEDiuL5kxAhtwqAyuIa+x+5rSGCE9UfVCSP
dxmRrGu+37Fpirvh+Gv7w8+P1cHx8YI9/StdNL7vVE5DXFFvfRYVV+nxfKzYg+uJox5qQCTYipX0
TNsv7PmOyFLcHxrUBcZ7YacQX3vARc+RbV3bQHzfpf44nK8Pft4vJUjAUBJ+VVo54HQl959F+WPY
CYBRQy3eTyt910eSA//hdEH3OwauUHX/9sxYyCDcb1tdOJ+Qc7sWWQfTCeAd58GgICygwaK+gy0m
BFTJTN/xR9N6Y8xizfQTkpvNsdVZmJz6L1uZlzJE8YU/2xsQXNLWMj6oI3R91J0bR6qOTkquJ6+a
U22Zc8TS8Fzb7WB5iDlQC7lRhSw/enKbkUBCgAe2aX7IcW6LBn3bFOjVZYcFci2VTwAgDeZAUE7p
KZmNNW4fgg++IW9kjwUe17NJqIi/cbRm2WhpgpvjFAkVG+SNQlQXUIbMATk+pjDBFPVlZdjeKfor
9ccuo9aZFlZkDQnwwdm6DMpuBm1CfUiNA8KvWy9sG7posjJrYiCMAonMjyZuiYzaY7hY5t3QFwq1
VRiwbWYWQT/f6519fthCFEXgUrSQGpzOnIi1axoloGWYTy90bezO8XtO3/Bh0+Vhjnvlof8FSevD
EWsnaEXy7jR7SG38gFp4vCDvNkm7FdvSwOXvYmCDoyxFpyFZsMPawvYrpoinPdTlvlGo91VApM+d
MvWHIw/RsBLriosELe2MACO/d97y5cDf3238zdLPoyFUHgnxIPxtsPKfUDQh2/tC1YwGTeAqU4On
03OGU8h7LVZPkSUpynrKURVBUzEFkiWGG+4XVzM5sgCqiHcZ8p2e6TR4JzWeBB/mN942z5JuIwaA
56m9m94rRuj3AnLL5nqAIUWp26eEysI9smNbbndoOktOkS5y9Ykhd4sZLc02OkwshCHlojXU3NKj
L5eCfu9FLSToIkNbEtdxXrjIQ5cLSwY6e63qCSgpw/oeSYodDGu251MWb0X+Ar0he65ht9dRuaSK
BEzITBgXbYgqyRO+lPCHY8cn6E6bvz2trc2khbs8Pe9gKyliE/qUQwmJhpVEuafLftmn7odHD1g8
lurE0s4aOs/axZ5zLpZARbhmTLvoX2h9vN4utAUI5F4yO/fE8PkiQUnWWWPx4nwOkGgdtRQib8Ha
hgR7QJiwCYbEkWDQLb6Kgu+QSu8sKhuUUGzGakLVsMmcFs8h1DncKm5Qxhv+Q7/CfXoNzvJugcrJ
mde8VXkx9MW09chU9MM5cp+C1BkyJTJKN3KdEsULvOhj35zqLNgn1r4v4HzThn78BEv+Pb69feVa
gnp9++dqkN/a1Vywxay4r6ejG00HzdxcM9URm/wXzlCeuwZ+UIT1pz22noqJ4Qf5mh/0K4W/jfpb
wjROGjaa9xnzJgP9poTA0783fGT8hyy/YFMStgps2akF+pvpo3bQsU/pkX1QduNm9Hh9aWEMg87x
wr6TgyhNUdA8F+u5fB/4gnEAOjGpsJnB7cMiQnAxOmEeZei/QK1xp/TJ0Sh7UTd8OFDbTAtfqFEp
dZGo8FclsmcqA1UjTD+ZP2hX+NEC+Ze750P3mnIzaL32UPCkqIZjDCSe9C4416JH6iqzUvG0DrxU
+Wr+ysNhd8Mnguma3zQHmBbsaOVQU/gS+VZY9+CZRABMtRGeh5giAvcejXL+AA8NfTkO27leSIxY
Qra5yXuX2lyIxhpyZIHFRKM2opklQYs9e9lBrGTQteSUlNRuSzHrHz+ynAMq5Dfp7lWqARAcYPwt
svxc7LNlU1XWDwpTP4zkcI+4FBwAqCkA5chaHYgs3QY72ePv4POKQKC2iXFFAarvMdAy/bO9iZGF
lNXNgUav5bDUw2H5mf6YNmfK2bqgOuWC4kLfpSa3Muocfsr8grI5ZN+En+iophsqAsHo4j5AwlcC
rm1fPmHQ0WDEFfat4rErKPDn93QamQSZhyPHaqFm3XMgrGO9oIBbhmM1msDq81Q6rGVPIhTMaHWk
0RDzbhYDeiCztr9PWNaEHS6Bm4TzG49hxoC7oxu8191SGqyYHgeG10c8khUEfX2ZJ6M1u51NtKz7
kPJu5zWhN7Gr27/4rN9Xg1tK8Gy00YbHVp9iaLuBtyYbqcaSjmGKbyspc462H5n3cc6Sdr5mck0K
iJIJQq8exqYkZESHCAcR+EeJrB2Kwrow79lajOG2SUvhDZxwUjabu02l6Fqd6F/9oo/q9tHk2FLZ
95rFFWNdKHOude2dt9Flia/WPqwvTHj7OVPxjmY+qsIBY22ICWzwURDAAqzDlQwZbq+vOrPo4qKE
HAJcx6j6N+UEu2Qv4Ndl3/ZkQD4U8N3hZOhgy73T3E5QKqNeqdgRhuVkp6ip3Q5WlIxBI4j58u3D
9A+PC5GpoA7LsnOQaqFBFr9ggu0smjWL2F98C/9NqJbKkfvpXHT76ysJ+/YWVptYGdAhNeUH3Tom
RtmEqrZ6NMmM1U3uwZS9UQJjnw4T5c8sbjXeuMds1Y9F5sJM34/5CNm4uDcnczwcNKKpYCQypBoh
t7+t6mcuyOcDTeP6pQseIMbVioZHM4ZexgIAo4FdLOLCjBpq0migEnTRz9YH9lwMga1i5ueIeFCT
SUzrCXhgvdMNJ4Qhk1mh648C7nlvk9pRLmvZa+4wyqSDI+HBiKpEjc3YtPbj1KlDXO2qIW63IdGD
6xQgsdqFYEDlQw268Cmhp3dRnyfU/hRxM1m4e/nS0TUHiq+XaLibRSkvxJmyvd7nu6Yp/qiJVdJP
M8thNSGOtpIkEITsFP9tMfSFgkdAqGADCXaF6odEFGg+ULdYOsUxilDo0pM2ARbkmWO2ZSvLbc88
GErElsxj/1N1U/MjDaBg1mb1MS+boaWq07E7VUIVXAqF+BaFOvrOxQjeNUXVAeNlwLbUmi5c62bc
KQwn3BRbAXLtrkUfMNariJVBn+BhjcdSWkpklHl1svedNdCfiytFIphcsyrAo9pM85kRqUO/Kx2l
sI/8fQqjOL+DVTZo0x+0VoZ96j9xgFxibr/j1/a6X5evn24zp48o2a4B2VCw8mjqd3nc2mDd66C8
jsdnyha3TlEnz+eAOxpSL4eNdxNcDFShJCpojluNH14B0dm6wnAN2VNIQJmHoR7iZ6E6HrZpxV6n
T8ucLAJN3ODaiKSJ1qUfyJ3a6+npd+Nfo6cdQBE8dKpXLdskYCp9TUKjDX5NMhQZbgiFiz4yw/U2
2Z50SBVK1+2kxUEIYykeuugqsugjYtTdxLbi7f16R1Z5MlLzyZSiLN4u2y2Gx1b6nasazATSYiLs
dR4b2YifnDnBjhqfh26WmU1ffA84Wddpu6dNOtDvIlcChlb7uAfpQllcSuiFW7CxWBH+vhhkTFyz
7qt/Pi9jHqgf2IPYljkFLquArvzDZBkyO1FNEf1kutq2TDFBG4HqM2PaColx2bLysWV8c7mnRIqS
fVL+hEzrLqMli2Ks3HlADv0LrXnczzDv72LXcbw+H4wtLrGLnE/K+uqHM4Y8cZZJPmWGLOndiPUf
RnWfbyaCMFQkHvku8w3ESc2AOl39KLaybN/1zpeXB45KhKgE280rsFbYgoph3FasICL+mKbXxjtM
4cbbHS9q/G1SUdVPHwQGUDOshJkq4vvx9ovUTH9LVZHiAyqxbC7bSY51Etd9O/BRIQwmbXoTi41p
vOpOTF8nxnlZt1rmqjSWPYlJwhKZxuw1iwPNgpp9c6FWpbDgFuLbzon3MlbhRw9NsyIo6T+a6ViV
dbLy4aYJ1qlbFHXs1mHX2DbU90rS+wBDFcJdIZBg8e6K+uI8JmXu0wGT6pubWvLmZTxKC6F7UcFW
0kKBFhOCY0eTwLK2eOL9xzfH7TP+XoiQhz7yDcGbdRx8SrHxKedlf3OmkBz2wyTLWtfqwMAlI+sX
YHMkRLOlLK/xz4j+KQO1yrJ3rf/gPRMUxkBkR6tjjHMINQcsKFyKAXBRwQUPhH/jGiEpRKfN8J5Q
fglIj6FByDjhTJTB3Ih2HqiqZdYD1tLOndZfclKtKDgE3txQ8iC6HfhFYj70wlOviO33Ad5zpy9m
MJ8vvMTiPI0YVmFAQfXV5HhyK/iziLdp0uQLaos8SNYVhB/hNFThVVZZ4b0D3z1l2zquLx2+Nrbm
Zn5PjUcXBzCr1RyDPizQKBL7efhDIlZ+OBV8JqT0Z52+yt4rIo7g6ChH9JDDHB7RzlLF4OB89tNM
OJWMBKVR8kA7tQCvgRmhm9+Qsn6ywyG6KgcIkmFdPRnfxKfYJZvBZ3vWNC2DACV8cmV27eoQCtVu
Y8V+m7n1Ig05Ee3GJI2aEp7huguYfbZo6qzI+sVPZCrE+wV15sWiXd3pN9lNZG6wSbwTyno2f/lE
cJ0HPHI7T6YVVYiTfWKVtbRMiOI/LwjJWy2tWp5qQ/Q0dI5PZVvlt9yPggIebfe0Kq9cknWHWpHA
5Y76614MCyO2e0t7Jx6LXRwLBAqC/8zEwep4aM7lmPltrxZYZfdNdWVTIqlrFqTtdT0h+VGTtoRM
N8HWW0wUhmPbey/cb6r95j1B8z9famfRmnDwWe9fBUw8CZoedzStdbNpiFitaIDWpdQxUufq1Abl
uiCdF0pJDnfkVQBz5YtTvnUcfYG21xtV7L4A9fZ+2ckWHV7+fW8MAkcu5/Y+hUily7vjdzBNHvGc
1Y8v8nvSXjs5httVFqXhbQvh8k/2UAbFq5IB+dWCtjAR5hmR9IJzxliOOBVNVU6HF+2bFkUBbro0
C0U64rvNdtV0pCuOqUKQyqhV1LDRViyF3l3MgmMLaunVLADuI0ziZFgTftRh8x4FQwlVDASihBSC
Ow4ZikYK109sY7ggKhd/ZQzQgh1zD/6pSyiMNpGIl4PZuQJ2+bwtqPdMsw342JYykNpMjv4aiGuf
jVgX7ACpzQAA7oDNO9ywRXrl5qcO7AAH+6h8msBOaQdjUmBjZ7DnoRBKeVyhtUjh3YxWNTpCVAAZ
YFHW7Je9bOqJfrXLzgBWLFgXEfn1promduJAT/HkYckxDqmJmYiQ3oXU28FTdH8MHfCXjkSl6mk+
14pfEyfqjWfT3lP/p9edQjL16ZqxbLxoPrlIm1btYp2r/Us2d1IYKBM/kb1slgpXJmwOrKXmP91/
X/xkXSq6epTR3ZO5kR2A7/NVVLikMjIK3M146V5XkZN8c9gi3/zVcANQ3X13BwK3sP/QB+FkyKL+
T3RwDtKb6Zz8zA866Wanr2wLcVtxnWufpts+pZNYIZ6mS2ie5DlDQCq4uZCD6u2UZ/nRXtk034aI
agl7OMFEed9KxMBMr9ufI/Veyno2lgE1eXh3wWVnbx5+MeVhkDzPPq8HZUsLSRdKXAuPgGBa43cC
fRvquTA3+gZ/RGbLen+SvI7lrdriTadvb9X+zlneD9O6lHTqN5AA+1koo6CtlA4UNs7wSW+Zol9Y
5x+LCqXTSqXE4OTf7SkhytGz87tA0OvbJgWP+oDJVmHdVV5pxrsbkWB8YImMGp5YLp/TK7oNrD5Q
fFxYGT/d7aKb7MYZgBI9s2pUBm7zVcD6+cvwKvHWRugr6fgweyUwHRUdIz4yWNt3YiKquBHSRh5q
qTgL38BCrvxUivyAq/2klozM1D4FCV5KvT90nzzOUJ4H38DlgYTaBir2VenpI1oeSMOScZtmxhig
v+VIQ+9FM7VKFIJDwXIkmHGKji+MtvHeyq5uBfzY7t43Zb920pRxe7AA5hXXO6Qdte4Zwz18uYaH
5N0e7cW63flCzmYyRYL9+BFEV1m+Bh3yzZbP5yccoA/XEhq/uekZxWqMjbNEg+5ubwS19b5UvNGp
9DhslVYIUyX5Hz/Cp10gzUCe47iXyZ6THXGwWAG7T095DBfbKsy0MghPBBKaecMATGWtxcJlhr5y
6h8o931a6lmn4dVDkvU01hV7nJvOwj9yD8NX9QdOejIYMQfBz52yTERk0gqn4M7V2yV6zogvO8AP
srnNRRUXJmtYGiDs+j0N1QclYLw22BK5ph3tTvwByS42YrzFQAtJ3rLbGK8Pt7yyFLT4D+tncr2J
+OFR/Fe+S5gp4GatD0+lyriVQkhcFPEhZqrgeHfrAS+37wGNWOFA9gUQlleXt6xrR3dZCtB80FZg
MEyYCucsus7ijz0IoaSQNYI6H4PqSGtieCRgcs+A+soLuPr1oVxwMQRrJL8AH6Ne7eaDaIGcHD8r
5Y79KOSU3HCVBViYVX7rQfQa+JjLtWjxN1yesgJdGDSTO4mJMSSsHLUIuOMlcrLfEzvr/mYYGNFz
9YJEGC63YRnuiMnVizaw3wl3WkkkXIZV5sUADq6/w1GL2LR8++yrknGdIXz5kPSMm2jVvvL2Q8GZ
MUKwburxKWGCj6icQJaod8Xjl4kOTLD9wb6BqpJVq+uS1y1dcVcKX34S1Nhi0KJo3STrzNQr/owM
7zPwI1pWPKBFb1ciZJihm2rmKhB/YVb4zAMpJUE/X66zReC2WfsIGRLrqkBuMB+k5hlwpl0x4y4Z
ibbScvt050OTI/Q8jD8WhXV1499N4kh6TBPPjjskO8LmzbX1m35vmfsss3XgJ/aDkCxqiOlb2sLZ
5mG6QyyuB+SjZjlSfrcJRsKulpTSA3EauENCSbhmjfmRnQrdY0mS/vihp8yvwKx0qOTNrrpc/OFM
kFPlU0Fk9A79O6rNOMiVYEbiTIE36frwx63+kfcLCcsB6kqwOEklMlHmTRZxzVxN3V737xD56rD9
9p3pJW4bQ41sj2UQwBK6tHN96/t/ZbU8WWYGiOd0K56u3OHoxY0XZKV5ZFU6Kafg1rO22VzUlqIr
U4EgViC0ua0cL7bkedWEQD9mKuMVcE6855Xe53/UptpNlXWtq07X9djVlBTmYsixg31w/rjxTRbC
UrjN64qHluo+IWGCt/wkK3cUsDZ6G8IlQnRrt5KGOdIRWSCv6MQxQbGskiJQMEwZyNGW8e78uVga
MYeZmO0Ka15aMi5O4fvru0N7P2Ffyyz4UlpL9ANWSAUL1tu0RZ3NW0dbhqZvMN6XwT6PARuQAELq
luPrOR+TItoA//Z8vUMNZ5x9MwFyV850qrk/F3dI/K92DSdgn0+s6/+l5XnVxqZxtv+1s07OyJzb
WFp2+Z/8Ms8I/XqzCRpT4mdtfGddHumkv4M3PBMN/r0Bp9RX6w68GX/tHEsRaPVT2j5ApdAhtedl
XQq9OEqlh0Az29y61ZZRVbRD5j0AUVroNmZi1ssM0NCanDrUpgV8nyQE2G+02+fPjjpy2fJ2TGEW
hFV/HRxLdrXOHBUao0razRgLEKzCRBybOMXUIkMYjNZjl5fg3fHIPIpQkvohSl1AIFo+rY6sn2r/
iuIFwEX8fBemdibPzCj7gEuiySsO/wQIXstjq7sIpyqdZOBHLiiUKH1wYtf7rMHWSWvV5SSzldOI
BqBDFUuvvaGzj21LbXpKrTqNPp2GxdECU1QcpxiF6GX6tX8pJvvt9HGPsg4VBvYQooHDkjd7+YKl
tF/qca+QIQ+LOrKXZ7gz1Hly3oPeCXbcQNW2uLGCEb0nzJofpseKkfjYBpjn2ZRWHlEdUyGXUP5V
OdCnyS4CVEtQ1uvugyh1kU32JqPjI2W0LRPCswBbmpGsJ4iKpTUOPV4i4UxNuHBPXxjWjnHd7qtZ
9D3FZKUiiDs++kL7JzBuCPcVrYY+RkvNwnZxseXFMzYudvh9mlMYZ05FAppCz3BGQHWXD4loFyXi
UJ14xDSmZO7QYTcy8iWGEmaFx1RGevbvov1r9GLd77+1H7a2Q49PobFtviMB0q8U7dnEbTHixsVf
14+rufSrZl4cjo1n5BfHErSmtXTFe6MQRIuSscJSvJ2WB5DO5s5bQd4fPx7WjVhXh0S10nVsblam
nbDWlkNgsMiowE86n3Ztt8vGF1rhkXlnKAuHWYoEQ5VcoHebDkKUDQJR5rM3657/PTH1hekIAQWd
PBzaLtophw44aslvGfKUkV4SDeEgygGFq4i07593l5Sod4Jp9FanEA/ZMN/YVJTwrF09bI59bROZ
Tad+fs0MUV6GA18VPlbcPkAOE9TLPu8dNc9LDz9cT4AVXjOEOR4H/ZBxNAHSUkqxhNNPDGmefL3i
k4OM+se5wrzI7hJZNkc2Z+A0qAaCRDLbShIHef2Aut3GOsu8eT/BCg/m4qCr5Q65on577Up5I8Oy
E3HMJnR9aAFy4bsgFn+TNgpSrKpriS9rfjQU03qKf2DjY55UEJPlnr35QB5wqXA7kLfY04oB220i
Pxz/tLjqBijViUqzr7YS/c03XXG9tWywcejBOpwrqm17t2hQLoBnKkZblcOIJOTRVqW5UsrNQwj/
sHOOPeD1h2Hv2eekPfRXuX6Y9AamWvjJuY8l4ORmGxOOqaGPkxT8NlRUHORC2b8UwakGzWWeD+KO
ZLotBuJLVKkSqjQFFcA5Syx97xMPzB0Q9YJydgllHZspaRA3/auEWsf3oRDrWmvF/iGVEQj4r6Wi
HahU1QV4dzkKlvGolxPp/BtbWUWD49ubcBp+ZQyDOu3vy+DlsBst1hYxTD35XpZZHZ5bL7kzRjsD
Wv6ohX28MxO4Ufhx4FYLOy1M7B7otKSrj3whYK2nlbh5z0UDXp3eYyi6jU+S5tHJSnlE0upwAvoI
yEJzHoh6Qx+VxKwoYhoBBjuuo+wW5PWnx11M8crUDz457qAIpb9OTAj1NkgSSBKQ1L0fshEGOPEx
jak6eRA9et7SSOPLkLlrN7ADUygeNsVW/DxXBQxElzizXe1458PBJyPpj19qkOJa2uF+AZG+7l6Z
wB+aeuKED9ix1QwH3MuLTRGYLjeyvVJkUUJ1ugBpd4qjPMBKbqWGdfGpx3tdxbx0UMhU+P6tM81R
3taSqaYzjFaXoDZByuDUq8ssTQHZrpXQMxv5pGFLGvzQm5P5RIGNODgUXpONqsKemnBLyOL6XqIL
sK7tG3VSejM7RmQb7yj3EUvWTxtuQAn8+LPjb1H0fOBdS3wli334vIpwSd2bnSDScAn5DbUKRiIm
+YBKsZf12Mj5sOaO7YF6iO9+qEpYVcfi3GV7p5O/vAEz2dg0qfYhGWUFHftSkUuy8ij9I2rn5tdP
HpzprLSfvitlh9LS5ayVxOh+yQX7mAEP9cOSu8bX6VOBqECmf9yHwA/IjSTypQqgiCrmNfocumfT
T9+L3c6Rn8lfksAx2Dgc9OeltKI/7zHb3wnJ4y/Tm6h2OCDRm9aAQdhxCFOcK+UFRyXuWqpAtrs2
J5cB24QVJ2ggU94UNeDX/reZ5KMAtVE1CYrcy2ulvptCHhCw2WBOG+VP7fv65zeEIU8FlxfA5cbM
/VcE4lXMMJV9+k8q1946l4gfeJ63NtlvlnHRjLHCv43rpc4TUjoYGriylzTfaZRwXd9FhdF9mevJ
NAvvszGbgRG3X7qFh0xd2skl/i11eyl39wVx7X6uxZ3wfHzOl/JzvVTPiG4sNx5a/hr2/M5bPam7
2J4qBmlgitBCK9U0qkCiA+VL8Wu5mI/Qgs4nvZfWkx/JpuAflkEAvBIVGke7pOAnmALvvzsggDeG
v3x68bdb0w9JO9a8PyzTGcahd4bF4WFKlpjvZfTUKHiWXkzTtMgmDMfr5myXi3QUH6RmP+gO8u0O
13bLyMsLLldy8tHOc1r66gloMOi+v9HlrVZi66x267kUYCP1+qdlLot61tc5uMTuSxcxB0AtaeVw
wgzN0c8WWMWBCjz7o/Pph8P+SyIXt2uUsHweCE0e1j7AfXQltFd1ivkohBVFKISKP1e7GGxMR/Eu
e/GMOoti3/IjHVh24+aKVQXDGzRnoTvRzu53mEE2iPI4HnEAH99ZACvj8FFntgI41EPisGQk3iRE
b+ZYWS19Lb52r2y1he+1GGGs3ksUAwB6odfUFU+vFtRHDzfeKEInFAg8HBZCiGILKUvx1lVZ36Af
MUz/MF+t/MiVInZxTiQuBp4ifHhzzZFHMwft8NcMWIh+ZrInvXozW2Y6kQnL1qoOTR4jmuUCqrin
m1P7onBXWJ+qxmM9ZSbk2RuNvpPKOr88/UjQ/Og0TsBbF1YbTY+xWuLWmhJG/LlQg4sMZ0No02/+
oTU3F6sabWuxKL1NZsfwZaKcC2tNcBqYGTTWEsY/l91ypzRbkiXCr8/AEEOPi/OXWdMq2txDDnpD
MhYaD9fYDa89eNO5KgZiZk/Ad/AGWbhIV9mawdJBFzAw9VxzMfVGf7wl9FzqphJc2LtAfP6M+9Il
6ElCNSUxnDBxBy0cwBVT2gl2pSwbIjh5Ub/6NxiRZHlPoPb2gg6Xc7a9sje/FijYI/3RqMq75Upe
ezjXNFxZF44cMZyMeXYUsTAa4CZZHirrZHSpihBkkfpV6wK63AxH42uxBYl0F3JKUHWmNu0Rucej
wBiSn3fBSrfpF8c/9jySClpZvBwidkrE67xBS5HAjR6tgR6hCTEGeQY+5gEb4sojMOeQrFBLTUGd
Pdwqz90/L4tx6urdNUkH/VtS7vjACHzzedOrVjGhUlMEQTreAmsxb+sIQk20MPO1E4lb1Q2RWodJ
ZFkzdgAKJBZYZ4l61e+OMQKhKtHBUvdgEcjijDe9st2s5s9lkzJmYow/ES4Voej4hOZGQyWsVEZo
o1r6WY65MIK2EKVjNuBkod7B9elWpoLAonuantRmdrukwWFKZbyCiYKopcRGdeiyyieUL+UqrpgT
eOFglOxegt2MLlS4Kd4pPM0kcZTF9wUUcJe/29iihOPiA+VAAOzjSGuwJLG/3ASbCYxTclnF05vu
H1pd2zKQU7Mo2mUwfm1WTyKNaj2pyLzCDbSYa9tetvqYqvFC35qswRzqcoci4sEyapGSTWzZMCxo
kI3J9OFVtZx51Lp64eQj0n9ZQ22ReraxB7SDZEDFZDYEmVqcD81P3WvuT6E6EBHM2U62m1dQFQ97
xYS1SSbUxDvkgXsWP2IkY/rCoEEEbGiS/cya34aYYe78jPqINQ1aTLGykTpE6mTULeetRsAk54lA
oFmFA1g+kcrRAzeS/4OGCCvaMZDW0BHJX6f+Y5ykFnDP+9tF0SgcPD4lYrNgjxF1v7wo/YKF0Dwe
52wvrUkFa4j88yTOY5303mU7Qei/jyDQVUZWZ906CSyZbEtXugVvBcLFJ+ldh/BTcGwZw46OLyqQ
tj+23y9wk24fD4SDYZalCghptsFUnpFrf/ES3aXkjnzJqLONUwh3XYLOm6a+9KsIiWqdTpvnLaUc
KsaNg3rciCGX1rYbZPUKvvkwFjWZC3FqVh7lpejRMijZSc5LlS5Lr70ZqRnuSXLPkdtRD4TWAEfx
Ct2j16r33//gvzhf3Qu//rmnP2L8BkpT0+mGYcOPGgqi+uOL8a/11rnYCGzT+yURTG4k8OVuWevt
6FGZ3Vsy+fN00h+ZfyiDHCk2Mt6gMpYcpCDsz3vn+rc3pb6GkO4Iqe8Vxyb4V1i1eyVQk55v0Ft+
eRjGlqq9o3vKJ0M6KrsMyEtgI8sduq5F5LMIP8cYtXtb/8QlJAY5RnZVt+5LRFGmwJOSzeGEceYi
+sjLWPTFz9amEdTpTNQ9QmSxLlMUEX+tELjnFaEB8EMDD4XRIdnf0Y9ErFQo5fhwWVthPYPWTogd
t3C0bUStoB78g4h0iegUF9pEaWZCLo7YsMruMeuoOM3t8vZsK7DXXryvoL2QVdhIPReAF2xfYk/Y
umvXdI0Yp+HD1T8Pohi1AQtW0rQASCZhD0jd755GMChnngQYKN9LWlElEVq6IlnpxLYBxVeOgH19
z0WU/4vFbHs0HBMH36h8LX3TgTIheUNIqH7pLCRho1/4F7KOoEC1oVWeM3ePFwYEHjL0cLwZOWke
Ejd0PdS0vO/EpnIFPQy06Jo0rvANMhMI8dLUX6YIFps4+9Z1qnXpJyCh0mxT6jPSElGwFeSRp8Tc
a7nU9B/25ywjP8mEE7hCyW+3dfvYUinInMSN3BR7M0p5R68wAy8Ph+xmw2AUSBWKqzV3K8s362r2
WcrdjZT1ry/U0qwpW3FwbaMClhAoV3k64SAcrsKYJIqt4Rx6ojzSkuSQ1WkyBLM1TtaO1ewQmi3N
vz3aOnw4XK+7fOGcNS+Xk5a/B7g19CUoQ3gjmWdZHvZm9/J9T2utP/mZgKBQGN/ah1WRhv2mUYZ5
tLVcO9Ac281/0mcwCpN+4FPVKIv+FD2Moj6B9RKwJgEsT68dZVmwspzf2nxztaDeE/+U4WDgOz8g
d64znCaOiDeLnF1gxbwGnmE0ybEjMH5xOJ2srQo8tO5Qz4ti8uvXfes74tNxBbxZLoq6C7O4vjPc
HEYzkI2DpvyAfS0o1nrwbLIi9GdKC0/WhPJZPR0hQtUZwr+QABrjv9WdnWVGovRR1/aDmQeiFvRX
XGKTi0lDt5IELYWqaZ3cX8LcAwIWI20v1s/ER1RKai0Etds4D+d6dWWrvLnTx/o3s5edp/QiHypb
sVK1eCidaIrAO+JNkggVGDYM8VcYHJT6C5LusCRl5/cupAinHamgPsErkFSL+o+jZdb6ov1QOmCa
YMr3uHkCJO4EYAVD93MDHCTjyZkiSiy+N8VXLYEKdMiuNmG4GCDl0fZpQ7ofXqlsWx5QkxUozoXr
SUPlGa/2k7R950ne9fAM/yeBQQNUXLLquVKkJ9LnDGXpV9EwoMoEtPOwDQ2Sz1R7dtrVECOdOejE
5CLtCk0EO/mTh8JOs3R4+/hu5k2LN6kkUd1R4YRQEEi2lK928Yhggb6N4/qCJ3fqh2DvwJu9+L28
A78EY1V92inUQOOj7njwYcv1gIzaaIX8GEf08RWF1Y7D3yX68poffSHWjNSApV/1qQA/iYqKAw0k
jRKZoqEYItadC36nGdWoXveIy8YSMCuHKtjrTh4JqL9aCIvtgXahnsdfi95OIHo9DZqHvzzARrDL
VzkGg2cO+MqDWZ92AMuz129r4isyIwbQ6OPzfoeZ7X8sTdsn96bvXsVF0KtG/VIKsIADfPYTtu0y
uhzIpFc3uOLDjpKj/ArtZejgk0LtkwcWnmr3WAtYDviWZa0QIUgfPBBYBAKN+EQCrVQHv7ROiuC1
WRigWKJbcgq8WKxk9afqesnHH1ZmtZKUfpDMjBsrAMzM3KmOZhRZ6miLl0sBbBzeUDALWIk2B/JV
DvSU8hlyRXIPmbYFBEkS7HEfMBKmpfSIYuJo4DoGT35ejjen4HLYUAKEbUVp7hfijonEqR1s5pFK
SRum6MzoCWzxzpcnum3UU953gcQS5Xslrr4+TwRT5igkABeDlaHHomfyHXLozkAyduBXJpO5UX8a
SvZIuAfS5zz/vRn4n67T70aZFafEaavtzP7b2iN1lwHRHDBJda/7luyCktnSbZgKZEFj5/5amq4I
0qmRZ5LeNtz1X5D2RmBh8Hc0qrDX3om4A71VGOAdvQ3geT8NNSSQbIIQujNDtZls49MUVYCO//Rd
xzLoHXmnrHeLVY9YepJO49jdJkvjchjrlVPesF0+ZCdLIuFVWODoivYkHxEqx6XdtLahbiAjQEaA
lkAEb/Bc3jU+E438PuoCkeTZZu+6j4XONci0DyDn3SWz0G3JF7cGeFguokReEgtzMtTekV6cOrws
HcsPLCyHscdaXk62j4rmxNEpJvX3h5vF9JgOi/bIl5Zp9XGrL7J4+kOFhaOZpGQDLoT88jfrMhV+
nxHSBNOvWQnuUZ/c2Zogtnt3yf5SsHKLacx+We/nVxuNdWmfHPFMSQZMV1c7tvZn6F9hxHCOZovd
4xKJajme2SLhW3ymoh3mpzBnPgRRP1AN2uG4rTxn5mupr2qa8l7hUVU2FHLwnGodri+CbD4l8wA9
hjnCgMqgAg8dBbZdDGKluYCK+H2ghTQBHfocfSbfUSkOHWJJQXGg9HXaM4Mlvo5PZO+sFW60Waxo
2AGE8yWm7enVrdPY6ZsRePJ9ve4WxCKbA7zrK7CAGHNJGyx5iCiSsd6A0nEi2jdkEsQ2W0TWrCvt
NSvZtQ+b6ELXsT9yUYL4V1YqRwBOrTi3JGCMNh8uGtQsaAKO0VvQ9R1hcpPv4bImLAMeyeYSe6eF
wKu0iIi7fD50d0rXWAiSQZOyrdp/mONPnJB9pjU2k+95XrwJVyW0SDi2lCP6wiE4qDrKLncJJVV9
RLoMe8qraJVSmADG33iNY1pEn1R++5mdqvv1qD0PYlIltjWvt8At1kB7kqZ+rLXa/VNPHhAwarHS
pFbE+lpUzyf7E/MQNf8udPtFAMishHh8wWG4gtfWnT1Y1d+1WWHhyapR1p9X08ny2rCFDfyIUOB5
gEcVcLnG9dzEjNjtrY9JX5obweqg4tZILFm8QsEtcwGbvEc8/ye32jiCMZvbMBflpOz8+2dY9L27
qjDD/R4g+CdPlahZyPgzt8y2VDbvwWO3sj15KLHkqdIpRt4/s5tiPxrahX2ycdGyUGdeYZlK2R+h
QTVnfbBXhvpOJf349oKh4N3IkjTKtjk4W90S7KYid74tvFb7c3u4njrmPqmYyibYw+wKLmHdB07x
FYLuK5o1xEcdfphJ8P+ryhRO+6QvAA3UZOslt3bKewx9NwXi5KUP9Ytz69lazFCPjYwefUSYLuHS
PKR/ssO7hbqF684NODQAZYWX+4tfb0RrlZn9Kf6y5I2mnVGLU97BlyCNRJ//z/mKS4Hy+BoLbxby
2RYWzs5r5QqdtH/X64u/XSMzWRfgYwQLNN/e8ErR0EJ7nio1s766WGtzR/wo56R3PkDfvkkEbREo
U2Ys2PTDdh8+D+b0bRVtXv04MzUd1BKigv6D8G9Vs34vL2X0W0Znr66vKmpEPQ9HR8MxI0Ufsj/8
j1DLPBd3euGZZkH8k0OC/aVk+Rp5+KcW9Yj8IBrUugJuv/TNcXLLCWt4NaROUSkWY1Vg6l0a/EwV
rpAb3icifz/FmCZYcQPIXJwT6nXn1sMSgGmd2V9eV2ymSqCJ+HpZDOoA6KoOT9SkeXUmnwOcILmK
hwV5rhyy3ppr3zUVcKb6a7U8ZbzJFj/lbSO0cwZOcpjjUZ3txlvQFGak9NrDgYbKujWgYGZ9gPaN
YFMqkWaLJAqtlFUMtJcN1c+V6uuye7moU9VYn1miY1QnIQ5ooNiWUGLWS1n44EVgr2tnPGakcA7Y
yr3P6ZDQqmQw/TzU2CQAQeI2NqqbRFg0UIx65843PC1NuSQHwL7dgBHZppO6UjKeWLCnvLZjaaUR
+rqZIVMjkGaovNCQt3LVU3qfyw948zjn2X4r3WGFUsGgKZ23myaB0FhBiGV2ygpc2zl7Dy6nBHXy
YA1gUblOuKQVpa7YZDk8tyDQmg1Xv3hjSxokJNGmQDu09xVHneAaJFgisX5byeueAVEeq1IvK70X
QHj1i5A1hT7d5I9OjMnb87BYpqKOTMAQMiJBrn4ZWXjYPxHOK8gYz3QXUAE5Qulx2LSbUJGrMqlM
REjnQKqwg54TRvQhdbj4VXXJ4oFWvi/YTnw+H4i3td2SzQQxZkbHxJYgbQJt1YBUpUbYxiEoRSA2
gBca1IKGBVFJn2qyNMNHO0c9g/deWZuVMLnZLlRxVEj1ZVDT8CVt7B8Sxe0zFlC6jO7ajbKXIMbH
c4KSLZbu6bmDDna8lhfFgWtvx4g2pQ4TK+fGRW1o5hqaOkQkl27GSg4ysx2U5XWOs0L/KtBU2oaQ
x8S1ZSajBrrt6nPJQzE1xrDLByJtnvQpsbx+aiM0nlF7eoZFxxqBST4TEIFoByY4fiMYmiTQzUpu
Zo8PUgET0FkDyutL+zOAPCaNsXN+ZeqPDQM4yRGic+2kjB6+Qjcg3y3czNrfE8j0azY433gA7AWI
kFOHyv62UIWmeF8NvkNhcJebbXQeHD52mnwaVaoi8mC1Bi7p6jWLh/dn66KhgHZZsdnQcpdKn8bd
5zb9KLPQ/tAtXcx6KErQKMoq8qua+qeKpR1B8fQfqPRF5z7i4vMIMjKTwtquxcyOVpaWQjW/yi7Z
JO2Jy47vn0ZGJ6CjAAWCa/XI/Sj6j71ryLvDtkOvFbjQ6Rvfw/S/Hmn0TFmjCZPjGVFd7RPy7n7v
feYvh2V4w2+qedoSpkxNveZ8RDfnKyJoxbiZHyM87fuW798SduiV3chzNUcv0uIURxnFDciv0q0z
fdZm6aV6ZWlweLwJs5OxowOt915R6z77Ec3PgXD2bWVyNXfiVneO1lWd5m9s+DK79joC60PimChI
uyJuudjf4R/ufpSeYbO7m6xDP4SZwjI5MPrwFViwjCG150b+ASqPpCr+PWFYHiN5vBh8KOoRzXRa
QhgMkBoTflWx/FT7olMaYIoI7I6QPJLSO8R/9y0+CNZHQMRN3S1qPuWzek6cRQ4OPyr6/+L5AI/O
PZVAXhWDiduqq5L90nZM0rZ9fvOMNy4EXt8TjUV8DFiy1u+iSuC/P704Fb7mXR/UvUovvqmbJWpq
0z/YPQlU9XKwtQJOWgCz/LOhx4I82CQCc00dCTXa71lHVdWFtbkQ27/buLitvrjaBsFldp8fUJGK
02/NJItTLpp33I6PjLXIE+pkmP4LeNm3Rcd8jvPjkXTUlR3uVZLv0WfniB6fV71TclZ0JmruomkD
bltrdezBuw7O+UjO8pvvH5bSOkjlLrwXYqVk1OxkiBK8HU7xy/ibWaB6g2gm5lsyLUxvk80bd/Vr
Tg9zUc5Q/SR+fErEXIFqV9GRY4TzHHVHLISbOK6hfTSUiLe8gChzCHZYOsll9KxTfQ41IRqu0cvn
2LTWQfPVJwvO9AMuNyCxzhDknbJqypwRRENSByPkpnELM2jbzkoHDHC0u7ZvRStIxvSME2uG7YB6
egUN13p9nzKbjCXQh1GdKMbGIGHdWTbhmJ//qgHp+44lBqslcnOXoXRikJCYMqFpeQatQDswoHqT
9y17DwcHLwn9TEXpjAbKnryS1s31Z4SrxgScBlvTPV6GWRFuWFDkBIa9RzSuDCNVMQjgINN6fyqg
CgWHaVZudp/T6vUmNrdilqI4pPBpRbsXORUp6gIZfC/Q2GqbsYTJyG1VCHfXO8sLiwdBd9PAKuHe
bWXnHuvR5bF5r5e013vZ2bXYSCVUJBUfMnwMQ4ErlXDskguxnuAujBdeh4WYjSFQu13yc3RywcVR
BSfOTo5FU/PE1l3smx82RdM1HUu+wuN1FhY3PD2Qfm5v9FX42B+CtSGfJrrXu7EqFhcAE6GDbypp
eWsexKXO/ZTe20y3jLiWmM7J25ewgnb+4+n/Hl6Bt9SMl94zYl0gO1etl/5klytONPrzuoMnvTp9
5S2upbJDK7BGetVC/DXJQvOc543yVM7G5ewkONKAX8fF8Sstbhf3YolHTLJ120LlBBJsCsAyF4zk
vSnq3DJnEkpCC8SimBAevWpLoZulzm0A6q+gAcsqCCCIOiKcf0CtEvQN0p+1Ubl95N/sC9JveNEY
iOaam25Bdi3cI2VQzLA/XIvBzh9l1jDSspn4Lqc3Ppzktp0ZLFgGYx5UwPi7Q9RDb+syaEYHJlOo
JGZFjQn2fo2ZTMwb29yzpBtGcHUIQ7XdP7jb9cgERaI/NPbKd4k1TvNRwl78Dhd6CRjBrfDEavcl
6Qxypvb7fzIhwui3LAyrw0B5Is/BCz3dJSffE5pRwSwXKRj0B4/UtQJ8sDTmjZZHGIrNn/b/qSns
Czk7spZ2YWHrcDYipVTlTSLpK7PJ+8fGIZkWLEmyrRf78NvIjTqdwEWNb7EYU3DI0o9i79rlBbnQ
3GpuDacqzM4Cry5Gl7oA4qapwNbFTMjMBg8gbxn216xK0Mw3Ge1o9xKTgjradPw9V3o5KCpGujfS
x2tR1q6z70HuEGQ+QB6vEvRqNcpYY94K8lcUAV7Sj3C/Dl9r3g+kYYAdwIQtkwhPyBMqQs8uxZlT
bB9AamsFSVn+drj0E3L0HwRu4CRe3+/eTdbAV6XXuvpKCizcwo88mODmI6PfaA1NkDtOtoMjqUxF
ezJbKi88BvQSXAxRieDxmt+ku7vpIAh0dblsQ79sdzhZqSeGy3h8Bh6Mew2KMrkw5VRjnh/mLBUJ
LdMj7wSVhHwBc8V3KrSrok/HBgTr9KGDVSNNtm0tnUaaiYfRytXD7PM5j94Fz0TZHG8Ap2zCpmSJ
PQMLZ46Ri70L089NQPfBC3k3VGCssc3yP3cscEaksCYfECCzM7gxv0VBkj4X8+H9WecQdWTe8ADv
4JPuG32OGOBGg8jyaqYj7xyBWAwoDYxq0EA8xD1tO31TejnKU/g0jQvxxHJ8WhJwgt5blGsCdG/5
jzVhUmyz8z8A2i89XV/xZiOdNuaIli46JI7w5XGRXfUVwNzTYF5p3CXtVfvgPX2CiaFGWWZbVJei
lge3Um1JWplMLG9jYLBRKBgCo2g6F+MCpn3jKZxoHdhGtiYOdSa4WXOoZGRwqAvmzNH2GI6Gskpu
itFtbPWO+4YGDchcni2qza5c/kej9OFB7iaHlVMEKzyBK/Nb3x9MgrPAK47o62pG5NZ7zaT5pHYt
t1Et36z3xM+z/a77hyGYaA5YqkI0cpvFr9MQ/hY+TJ6jPv4YGHCdE7ICX88hHkcKHMXfMATnFJGl
N5WT1IERQ4JW/TcbkGIA1FIQlb94v8IcqGextCtTIM2YhCdj+dZird6XQb7dZDdxZ6TtMGmtWWd3
FeBfp2BzML0d/0u32v1v6PPse1kzDphLOKxyGz7X/5F8IBwVX0X3YI33m7mKQWnO5hws8bL1ML9r
bbBqGUxlKMb98gzw2wXqHHy/Y1Z6jcZNmdEkljccbh3lB3+3Et0RwoA60Sf0QmRrb8KLd/MqwN3k
P+sEAE+dgjLqr7mv/q9ec9m4L0ARC57u/x+bF++nyyabL/aykZjkmQrHWO0574nviF6iEwezbk7b
c9Q/Z2aqUqQbXA2zu8Mf4PSY2UQHgeI5bFY/4LjHAj8gk5If5ai0VJqQec8zk9mnfyFABZdtUNSl
1o75+MBBsGwwoY7t3dWkqfzzsrUH71n/MFECyC4MyVi+uQp1jzCq9YlaTKDAZAAfb0qQG67ScAZa
Pl+JjLdnJuCTzapgnJPh6dI49AowLcdlbDZpZoV1qpFTmGHjewcw10rcK3EWI4renz6KcC/FrptW
zPj4jxrWBbR5k7zsb8TwGRJsxpn4rrWGV73+b/F3DWDfPIN42vISVceykLGAWFR8uOpZxAuPxmTL
hBx7LIqnDJk9V8QU5vsOfXIwDdc+BdPXd/nvJXJZNWEDEo78Kc3QLBcZnesr0kCepUCioE+X+O6u
GUeIBf2IsMXobBktpwG5SczeXgZNjr7YOip6fb22ewmAD3bR9RYIRvuMFQICJAgKoDXmr+JIE3vi
l+rM20xvN8OmVSZ9ezTRNocCZ4ilBbPk32JY0jaHO+kuTmHyMDsUCkAtKzGQBod/qGc+1Jgjbv1u
Z34oJAqs/B/HpMV5NDW8RKKu7jAk7Ps6kyxz7YlKsrwJQfa1XEVp+eKbF0PdjBdnyvG4PYENumuR
H5Z5o3yiFFSiLCbrq0MhHMYvmAEnUHYw2lyhm5HrPZDYP/NCCwoqWXAaF0vlAvguFr1BQVjVxWo0
9VECoZl8DYBJY5qP9Pe4mG9n9tNnL4ZZ0p94pNi981cy/Wef56QE4mhVUQRWhu37aHdb61HOa37R
+esYWVr+4ymKUNeaUMN7kOsqA+V6A1+m6hjWUFvcJLmMS27SR8GnPsWCEsL4eTIEKRpBBmmfp2mu
r+tqF3GPCXfvHxOtv8cXZbOgXriwf+xQ7woVdKoZK/SzwndS2VJY5Uwi592WeuF+HzmSXv3wPkY4
2xLtrN8HIvBW73J73z6cS52hIdIeo2mi8zOZ3NIJOxuo0C818qTaedjOAJiHIhi4cN3G0inx6YpT
tDmhpOFwAHeAN4LaDOrPkXBmzPexLcJT6ySrkWH53ufzE9BooQph80vpRhVEMYFYg99dMecrLv7U
EBXzrSgOzX5HZ5IGYCDhVSo30sZfy/gwB4p4KKaEEOdnTN7MzOtwkAbEkpREAn1htQIJIbFpjvAX
EuO+97zy/ZRcCol91UZyn+QjgWRn0YIzHQY8U2A0nNebE5qWDGOXnM384iDZlB2uR2/CpwEVEPL7
0OqELad7LcC0vccv31OX05/gaRQE4Y53fueSvyxXSoAYSpGneDnaVs3wCR9MrhDXI0gY0uh/x74l
wzQ4YNPCU2ZHfd/bgCCLwukbrekSN6AZXYZMwTVIoZeW6jIIX+RVLQTh1o3rxlYj8oWYZoKDgp+5
8PxigmXC7G75CBfsDEjECmolY/g/0gB1UwwUFWAQ9aJj6E5Hc/91buy9J2tNmiWK3BvVCrwF1jAD
RfARxi9e4dYvJ+lph3NJdfqU3wdW/CGi4cCdKML8vWN81ZXCX66m9Cgybq1hniNcJJxOMQd74VYT
0JTRJ8UqPrfIqjHhnREBfAGM4yElZvVQIO4kC/UE53xGiy2tl4W0I4iMRiw+TiuWMxFQ8u7vMCfn
k/HxyQjdnMs/3pMdpffJwKqnV22ff/RDxUQCE0fXvHsee50oKGwK/lXjnW4YJBjCLJxkMmlUvkKB
gIK8yebk/zZWQ1hMDP8pY0SfBOzpOvJlW/vaC4tvm5PNl28ZqMaqji8qkWXtOEFSxKoc864unfku
HMfvUGMklQF7h0ztu0Fmvshr8drAc6U8im+tGm8D/JMqp9jxFZqr/cB/q/T6480DWZ0hBPuS92zR
g8mrY9zkWOoE8QnzDmhxYVfyY1rIFWGZQRkQMJrD9Nt9+5PqZuyp62yyafNiQKpaD+3u3L8FwcaS
oqmeMRCIu2bBk9iPsNaQJD5/eJUSBWmt2DSeZYZ98G42jX1Vqc/+bOUrnxdV8GvQikEo9lJ9stXp
C78S7XXMOYalcR4bbuilkzGoiLb+nxkEdN4fwEq+21PAUlNaPTa+bcYNv+5aUuWTXgtDnxxIPluG
NoXgW6MqjX7Llk6qIEZLcybnMvOdypp4d4yddN4OkiqLPCv6eS0AxiV21hEJnCWGDc85UrlzF897
9DLf/ygMTmh5YKOuB1y+gAJUAU0lPt84oq89QChLSE4PPUBGwwYZf3FELKHe+r23q4H9GjeZcy3e
wspdNU7335KpcYPjiSGwoAjqIf/ste1InlWBU0aIWYfnUmjITiGqHMA9liLL8Y9aO4r4HkvRO0x5
bPPy2qwofoS+aLgtgRc56HuKP/kN0YU31bworEEzJo9NmI2JJ+Gfl8mha4yY+Km4CaY1+i8f40JR
pozozU/pN/uyzm9oiHN+C5v3zDmsODowQdVaVx2kcIFn1N8X1Qv4/kiMnpc4zpUcFr4V3PTDURCJ
FZ8rexAXx6yqzFyWhhQgIpTB/IlB9dWpuMXj+cR+SDeG+Zyhn4bCKfwrVNLxuK/URX4x7WPuNS3s
4PLgzKBdFdjsX8zy+cwks0wyzcb+6pVjeXOD6aVCYmSHtpCHroTwobofk+1R08K0CYReoIKo63pG
g6hFCXGNx2Sh3/TXJA8WNh2lns7/qqfngZqsDIPy0a9VtX+a4PgxYKCfmZEa6o+pmbL16j22htuq
IPp7MdPD1DcUqhYfZzGTezojqtAemgpUdKGhWSoS8bvuazQN7bQr0TULh/ijWzSg+TGgQJIy0ppM
J8s0hnH8IMnKiyT3Wb0n0lOSyVXSQJtk2A9mTLigIh42GXEw0VW5jn+l2pOJQixDUkfF36rIi6Vh
7vVABvhvhcD4MT1Ts2y1OXJiJ/FtMg77odV9oZtXvqGOXjWJvKsk+tjstBvg2VF9kHFra9UB+o5z
tqUKcWdfG63+2YNJW6ixfZ6NXsRj+uY+qXJvdN4X6G9nFUlO5xDk3kwmHorQbzRLxfkbqi95HTVX
cJq6vz0YhSLc+w+DmhSnIIj2zHST587s2tQqbScFoMnhz2om48oST4bxB7WfVsomR94PlnDepi3g
GldrGOb3QaHjsEanZy6rYbzOmwqH6kfE3ZMwo8Zv6QYFuMORCPxCdCjq7ITN6WJXph3I7exbGJeg
XSGthMywsDxbhzYjsaRuQWsvxWl7w8vHu/BdUbgEZ9bHebMDTWGLDa4aqodt5hSV9LA8jjgh3OFS
IYVFjITgYPwPvyh8y7+tLdqdpBv6Y5dYu5oPgfym2nP+89ueztLIZa67QYcluyHn8qc2fVgcIIIr
6MvmsYODGNEFS0bcSDTbJ/ZxQvMgbc+ZVViV5LaHzPcM2u0x+RWPaIXfY9Z6mRnQeihzfKvTURXA
x0ENCUZvfd4RdUPwYa1ALRN8CNXQWKgbGW+y/TKOMW6DEMfezoRHP+EL4MjILX8vPnvNg5MI/Fhn
dvB0vUXpzmMbAxm8npzQGRUT1PWaBg5HmqVwcjWei2vLQ2/H7LjcHaWByejKSmmYAzBXCY5xchau
vEJsDz5X8uuFebhZi41i5qnRu9zIVcfphtVgmso7Sr37vcS+Lv3YA/mFJ/oDfewtffMn5tQBFUNX
AAyfIsHNTDx4daBckMrhGKX5CDFtKW4naMsM94OHjR8Tmav6wJwPoMhIOkdt9+AwGB2Kv1ez1k1F
BL/cU3xpOBZ+nM1k7SMZ8hLySlvMdAeozNjrT4zI9tdPlB1yM8HMnvkb3Cil3ZF45qylD34hM6oD
nsyb4QZf/gwtHls4zjElYM63h7GnNnC1ZuFqJA5m7LqAB8yhUHiCj+2GLnnMVuVsQvbw1Bnh8vHV
2pcPw7BUJjiDUZ4MjuClkGFVnMsiEm6RN8ZP+mxY4lvAlnrNgJKKtnOdVhzbtjKRf4XZLT8Oz0mc
Nr0p03h+s9q7MJJQkuIzTIPIznki3eYe4h7e8SISk4npKEnfRSw5p6wLlKc1ar0bAzxoWKJqxaTO
Whrkf1GsLrxun/l4PiFbyB46pqLOOANyu0BykKLb0qYO231a8HfFd9A+A1VaZuLHC+6odbmRCknh
sdz+ETDdze/SMl8Beu8sYNg5a8y8XpbH2fOvJiEKlVUPR5l6cyWbRZn5gYUxXVfDIyYPF5iSi1zq
SEwS2oYH7X05PutAKtEzsbAXLztG2VYiWHYcsDded/N+zb5ucZvAQNYuB69tCsHpWfo4dRP37W1V
9LI9nX2yo4qVvF62U/vutRhbNj1JNxe6i/H0USg7UkYrpTWUUO/XYUjBvQts71ivsvg6jOMk5QeW
D9CUekDRxZs/iGOTw49Inc+BlRt+Tdd6dB8konw1QtP8/abM74E3lDKngjC7mcd2wbnhB2my0uUJ
k7ugt4Fy7LjOdFacSvhsXXe4GuCumeN9WXQyJP7t8QAZ8j27FoFnTdUGEQeK2euoArR5VT4LFsZ1
WZVRFNXmeI8PTDHQOFEAkx2EQwAOKAeUlx5sXsTGp5J93wLM7e+yqqEZVGPa8auvmk/eipOj9PPj
XtVhw9OEDDda+F6W8ErgQLYAm5E5DR7jssZP1wX+Lsb47jpBayZf7pqO0UkHcgcaGk5kPkvevJ7y
/GtOYiameARAuDsgVufYqgCCMhvzNM6Za9+h3rs50ycajJR0CvTjbH+vhmqqEPPxXYoFc4a4/Lr5
QLKkdmQJvYZ1MICiviAtOe6DwfzJKQrW9yxSdcpFJnK+gtXmMn0KaBtjKJ42WJrZ9HLPWZC89EcM
T18MBHlQliA9b6jEXZqYUdE81MbpT3M6u3UwPhooJyrI0Qlo/pWu3baTzBLd1Sf/t/gQDP98p4gi
PX7rqXlp3dyzgyVZnUi8r63WX5dXVFMvWi9dpJNfk2LOiYOpGmsvd9NimfwXgIT/ax0OnG06pq0g
PicJHl7LfwiQqEIA2ENuPwjTLzqO+kzTroryopQTDCZgOmhjYxZCO0knhTD5qZyRbHCVVfnfsjZE
Q2l5XS2NxyUj2NwYZBGPbZFtvPWuKmr97h8hUjMaM1741uV6h5b+BX5FpZRSnbijXvfEyhTLLG6V
BTFSpttmDBmdUR7bDSCxXYpNZG2Jl2TcPuE/q6QLr8LqumYF+0ObGW5GiEqGrWphVfKZvqr/26iI
vkQCpc4iNQEMVB3rVNP2PffWMbX8a/XiQGpEdGuJo2EpKMaJSWagZd3KgsUkd+tDgq9n7Y+3HhRg
xaYIkVlCM42rvOD3i8MHze0MfPvST7ESaIRO0cCclyJr8MLwHT9hyuLb9I4O7mbVX3rsPUwbPVzQ
A5m9OCP0a0sMapdNjUKR0ZzwQVP1Joqu26M9lltrtFZCDbBm/W9/XXtlHIh36tAs6dwkEpXi8pCV
2MO51/xJmHKwsTO9fhtEj2p74J6vdMnH1n/ghwYbxcyG05FvxRR/hVW94TnLIAJ7HsVTbLlAElKb
shh5TFCkDl0MUB7rIPlpzRIFUCND2rw8TaKxNFyZkVA5ZeBmo0dDhuVHk1+GcoPd2RqIIiCpyEHg
gg5cVMNinfS/IhK+rdhz1OxQPj2lWvQ7u1EcCkPPPZzyIJiVyyr//LkHNS3MTXqT0PfYnuE6u9Kb
aoqwnvW0oV7FvhZuVgBBfPEMZwlcbfe5ROeN+EAvEfVtjNBivYNxJNq8hsTsHdhY0Au6E2Y9kzoE
3goH/xQ1ZKZmwn4PAzmz/76qYZ2+x+yxfMGfYR5X3BGn5uBnfnorY2MfOp9uU/6unGNBZ1rfNbyB
PVlV44J963PFBO57QEVKIooxU4463AQqPaWngRZYBMzkg2gEiTpn1HLzF+4KEpeYihfVXBgOCiHR
7U3HIpL/sJFG2oINLyBK/5wDRp+X73Ccm0qH62gpWYOVBTw2S940G/oLhNcx/gP/cEV1xyRBdp5T
AbRuSmOk3QQc8bqEDzacd46UmnekH+ANrjbjelyq9oYlvhs4mbAkCGVAwvuXVBASmVaSXNZR3Fpt
XHtIZo+DMUJ6Fo3038UCxLINJX70EyI9ueld2dMNJVL3iDNxOSKK+dEZJcwaCC8MTWv8y9Gq96XR
ncgMNmy+BvNgf3sYg7J+nC+9olGu5xDl9uEsX0dNhNAv/Uuzt0poenXmgHZQopBLs6PLIwKK2oHQ
QUyQERvwrMtKulfZCHaEw+siQ4f2hHUejlb+af1S/WqlREFNsBVegOlGTfdgq5LiKMg5Lse1FtNe
BHKCj/xBG7/Xp/iUVGcKXrj2ykGcLXJ35S54Z/AnbEgJIbH4kpXGiqVXQD+f2L0zVLS41zaNE5pB
pVcMDd/hT1zMr0tllnpxtgOb5swVbBUNq22FsI7P1Akd06UliaXlUk1lV6DThc0M4Y522KUNmiTW
5I5DR8AKwmnFED1gx9+nZcGpaIHIGN88kuHjMgKTyX7w/5GfClQyF0lfKhZVG4nFLB7yWO+WBZsM
YokGGOLGQLr+ffmvjPN0BwO1QXIxRDAiBbgseBzG5N2zq91vB1YH7XrBPtl+1KzHaa7prTQGTMfz
J0D224FY/V4c2aDZHP1VCaWpsA7RPgOdcSxPBjYiZV8lA/RABJIdYf4ae/9IJnGPad2dWlhVUrv+
i6+AIEE1kDLgjv0qUPSYwRTkmNaB3fqoGvSVPOEFsgU1Mr1l8+bVyDmLJb7iXnfkv0LR+agPYXCp
5aXxBOeMKOcnhLZocPCDnVLNSzh/emC/0FfhCv1VijvImH76VrVKYjumCZVyipajMZXSTq3KDGp4
GXmB48Q65V2uheT3UGGpnNQ/jKBFIPGYDh8GKAFZ+cuWcGpe/oXCelK5Ol9W+8RQLhw/JdcRWE7f
DlmuandeeO4jT7g4WyOl9XMhXVIxjZ415MZmRy9VaiFjVwHu/wu2ZM0OMJ/YcRm6/+VPXcSOK40s
z3QGmm/cdcurM25xdvRIquBafP6bvt+v0aFwa9iSgpDrBl4O/kUC4rIRAo82cfANNodCpnwYtIqT
Mq4jsAGn9JCcEMn9aJg39hpghR58+euM766H+poUUtQB7XwFoA6LndsoGFPPOjqDDvycEJ1st7Bo
zGiOmHagju5sAfrZlYbw2Y4dT5kox8gscDpxI7Ikb7GLH4eI6DGEr1GiLqsnQDaWEleFS9F4xnXr
98EtKnhYhA/5EJmYWQBbq3JmjJSCHJj/iZ1n0EaP33OqYfmeWDthEMrYndqTv9v0QTfTtWqXkz6P
hUlPJRfiLa/1dSdagdOEeTfkhOjclsUdxhjOU/ZQYLyEjjeywKDLaww+Qd5Edh3pR2jN4g0pZZhD
w52lUGQtu7qSgw3OjwChAEghWQdqxkqxxQswc7W97GJNwfof2Xc0UWLL/XNekBm7hjK2gRRaKGEZ
TVC65gpRuG5tZQI6N6jJYYOhMTSRNO0EWMhIkLO3uwupGHNYejOW9uyKFyleJyLh4jK5o+Bx+OUk
pf9Kx6ErwAublPQqM/vKKnjAmTkqnpaKe3TlDieup1ruT1CFB+IFtHZj078vW1MTQZR/6YUKMbtD
WCaFhhCGRPqj0k/j/ErVU0FWL4m9oPky0NMAWi5Qoq3kMZe0gXxeznKVhPtvEy2P6NJcriclEn7k
p3cCwM5reuDos0cGTtTU2frnn/R9X/gAbI6ObFEhCJJWOYcX2WeFWmYlibbCqguhfxMMK8g5IkAu
DhPX0BiM3MRPrIY2Oa8MEkt7FaBiRBqprVbcJy7gFVCPyzRIA2uRjaEp8X8QQHPp9TM6wYgUYXuU
AKjmtRp8NMQGdg/99vkrDNZ83oxzq6/O2F0LGFo5oGfDqTQ9kDixL+n+0EKHEMIeK4rS5tlaKUcK
CKqn/pwOiOX4rMjh6BEosbATTA92fQNinwaAWLHJS2NGH6KLdtmZe5kQogz1/tHepskPDAgKE+cQ
4d/6jc5HoRpS12QaI8QAAFEs/25+fyPAKiOZlzdi96NHGGrbClf7pJDA1YycqrXhV5iawJHJ7i9f
GgIWedPfChZtoPnbw+FMkJCYEkzOFXmGZ2kg9TTm9OyMe6EWGUlzm8v1V3GGHWVytb+v3AGI+bYt
oZ07l9lYzq+rAwxixQZzuNEIBTr2tKoCcxQNBW/LSE4j6sWi1lQkhxoZZhGNYdga5Y4EXy7vz2AZ
WTaxKl5V8G1cvPerMbMhXzaMxzU125AofPSz0I+g8RHAfiatC7lu/J9XdnsX7U8XaA9lZZmflQBO
PNz7RbakVw9gFJ+qLxMxw6ZsimGa/yAvvUg5MM3Z1a+3Bi/209dD4QnpgUGlFFCnf5dbjn6xD4Fi
cxwYVsXu2PTYVvRys43ml5Txq444Mj2RwrOr7Pnu9s4rc9dDeXhTR+yalgrZuYlBfVLTFfafBo43
cw+HZinveEJdTC/M0hsMwYMX2/iSW2KeFmN+v7tX9uo6QWYksefoHvcu6wMHmqcOkWUoMLvk66la
83QhgP3RVh1XXFxx7tEgfun/+KbwJgmsK0az6r6abiXQxObQ98Ycx7WReAxKjFfY4JiGXOZ7te/R
O3OOjOPPicU5Iq2E/W8c3jAGOoq0SklXr+sYkR7Fu8CuTyM5d5SLGsmQeEF1rMi0WSQy4QiL54N/
iF0dvnkgRgWcDpuKiwACfWuHg1rEuI/iOb1wuE/0qvEEUDRrzoiwbC3QYeDc0GV3TOvqYYx3e3/2
k9HJW8jzNJMEcQPZJwOOcFc/kdAKShLLgRj7o7LBt9tQkdBiPXFcHp88xVmJksnb1I8dlPSbe7g6
E1SujkW+NgHJ1gHRADDS+1YPDuzwHiUqnAZqY2WM0sqqkIANND/bNzLbuNUpzYvOy9mQZ0h3FDM3
p53bON0R8k96pr9XmE1+AeqRgSutz3TdsFCpkUoFopNnHe1AjOoEIjQ7Y4d1TA2B2O3eWuCjIqK3
MG2YA6J9fWE554X3gOlV9DudGwBWNrurCQK4a2pK2+QjYmRrzRnawzSdxZptmq5KD7TbZruyR9Ui
Z5uvKvLY+Z/Jxr7i8dgfMgJKcGXPICA2Q/+U9ifxTQG3dQSu2+Bloydr3BWXgvPhOk6CwINTjHvq
HNKvkL1sI6FCASH8d3uilHcP0uUMrn6XWM2DJtS7DcVP1vIP6qoexIfBD3NkToDbpVMo6PZIeNoA
uCPcRiUDyrMVf2pWauupU1zBNI4WR6WLq+oQUwhr7JI6UPj7aIt2tEfOHCmIegMP6UcNaR+ED/hR
qWGP5tLcnHe5V9P0kumHXgSMOZ+Puy/d9+1Y5lw2A/iTVPakREHEsxATuqc5TpvOzbuScodt2QK9
2ruxLH57UY6jo8v6dsvz5LHchQ3mGbVMEjXuCdd1ayS1FwrX9W45dFw2PtEZ89BstkBuz+nNvxg0
u/LLjLIci614UgiYw97rUXF/3hXfWf9f0mi5D1REt1eU/r0RGduOizqlYtHE9IGecFm55I+eIcxi
pdyBaPD6ErKPvH4Pc5mWubhUG6+w+5/8rZOndiE+7Bld3Efn+I7QfnUUqgAKPzbUm3b3WG57gHsV
DAlgxlpVPqvxCCK7wO9dowENnOBTIO2XfTjuITtBVx7K12TImPSrmdX1/nkmvQYH95+MZnIrfqtV
U2CwRQvwAw4wYt5Rdhn4fuD94DPJpjIgIsVfRY2CdjFJLe42gR04mKbhieudu6RJbgFuGXZ12OrA
7dLvjvryQnX1cqNG1n6ky3oHpqTMGup8Fa1V9izXujt7BWIq7KfIWi9s+03RzdOjQirO9ipV1go0
CoDFUxT76g/giSoVs9svuUri4lOz0ZLUQS6hMA6+4ryj/Jis8InTvBn5Ngs0coE/KBIczCtHNMdD
XH5FvSv3U0k3scD7TkP65PYri1ulZnZHybIoeAJKm36rYN2rMJYXCS6zHxJHJGp+ryTDdCKhYCuT
IQFBWOfetfK4aHZzcki8yXcIPEigNRzLRQqtloASHWo3k6d0xeWR+63IJNxrSqqpcx6KSG6izR6E
9uINu7ICPSALmqQASZjua5NHCftO+vEtlzp+kdyf1/dDYLK97ucw+cv1h/oXerX4yVE6LwlQAukg
dGrI9ROt2GVYmeF/AEE9JhZg5AHNpVQFtn5CEsWCISNkDghVF/tUeIxIortyP4pMAr+3qKJjmylY
e+/MDJKzMwA4Zldpt36f67ieZDOpm2Vfpx8jKxp1doq+pkH5HzL71ZSL2X5/dIdp1byfZCDRu3ib
1Nv6eHENcfcsIWVLeXOEuoQRmZ8RtX1ZqTuVBLH2C/jI3K1ah82mhaZVBxiP1gHj42UpnlDRyqI0
yyNaTZN+3zoaJD62vEza/o96eE55SwmUwuMznyyCP8GP71ln2R7HQ6IcOVRGgL6JTeD+QQkzXEtr
W97ww3oJ2dVnd/GyiBph6YNcUDBPC84m2f9BCxnajIqcpGXSYYf+3fRTynXBpvKLyST/Kqk5QkBm
o6EeFrLaUn+6EShMt6uSQvi+EuR17XJF5CiCJobX2Tq2UATs5OEosGarpWJIy2MyBF2bk3xw4rS/
1ldR8Oy2ha20WghQ6Ge05mTpnAD1smQ017az/UDudGYuUqZUBnGn4GGWknuRSAB2fhL6boHcxv+f
L31pRBj0jnECFtUjqsdbQp4qrzBy12O+LK1hw5CNgZPJDkqEvwIKRzDQq0GVv6HvEE0N6LwKQ0U2
HE86IhilgZBRig7ONu2iKZIjo/b/ZGA8GZ6Ocyw5VxzTdjmy9Saw+l8DttptUecNqj2M7296trbS
WkzzaY9WE8XGpnX/wWL5NdUDSV1i9gcyRI+40IHEhezDaSzZJ1lE+B0YeAKXDpdZNgmqGbdxRZbT
Mxm8YCnWCV0OJ1hQtRqjEeoHi1MfPnJDCIGNuSmWA/cQbUxbuk8Aj8114iAoya1DMflBfbJ6uXkl
ZVIuP8fvccaRS2G7ijbT9Za+d4UzlBWETzhlQESI1HOimuSCQZdht6ws+lerBpVTR3+c+yIvs6H2
/aI6w7w+3JpoHPA9g0Ea8zVNHbXQYl7J32os+OWtwEhd8W36TcZqqJFLb19wlokfZldNPWPN8eZq
NtTIyS/WjCsIxAIjn+6rnHzoKSVibLwVoueHX8Eb4Pr/sQ09co8fXK4seRUBJp3nuAEx1Ha7Nogp
h5WLlH58ac26g8wFDEdnYwKV50V5nAvmZ4H3pNB+CD/ftbvukuD/xnRSUQBbPUs4hXoaDb7XYQd0
Zvt0a80pbpalNRT6zRF+vQojW4zaDFVWGZ9W9rEGaLPSMpPpteUAy5f+IcFRwT0mLKf+5GuwECu4
IAsZX4z2m8uel8WLTp3oJ2+FpRJUkSGfdvrB6p7HTMh64ln2Sto2o8opMJYUZjw1HDB8VSMk/RbS
3VfRkYO4IZtQUst5XLZaM62JIGx9yLRaVF9Ze4FWBGvU+/MtRvgLscp/TXI02j117swOI3vcHAot
dvhkTWUXlJTpCx7qp5GwF6lfjgpOslNEnEqhC1k0G0hgvLzjZT15SYSg3NGrWZ+xnMmfWEN9OsOo
pUm2+Js1sWWwsjyze6CdpwZU3B9ZsaoWm5RpwDjWGjJp8GLXHvYozTJ3EjIj1XeHNnoIm82fOsyb
JStYPuaJrYrrXuxVO5yFzPMxkzb7s54jF57/vKkk26RRobbrSKAevU3vFTEovzVpI8P4srJuHYdg
r2N7/+kZOZekMX5o9MeG3Wk1iX5cC/taWeDXL9hRHFETe8AWn7SnLYpomI1xIb3tg6DxOUx+FYnn
0oOjqj6tIu+WoTPyHwmjjAZLJyLJjjeVgNdtIkjn0g7q8bpIi3VTvWMwLl72G4YBcsSumPUQhy8z
Hlz2PhsSET8xdseUYDZGgkbo9r1IVCCGunp+91i8UST5ZnJgPdYesKRJF6hWKMqsoJPLGTc8E+n4
bMv5jvM2+nFuU2UeikAHQA3ljN4czABsemQ16GUIS8REOzPaqmC/RdkbyL6uyhspf0XF/8mq0g2x
zwab84Kh85lwKodi6RH5ewLtUmYwYbSYuPJum0PTJ4XJd2XdPn+pE4k6g3oy4QRbyejekxeK2EUN
Bx2yT0dvcXnlfBDJaXCAXg8NkoCB8U5JCJnq8Dyd0DZuS7+x1DzW++ofc/FcIOdWJ/EkjZRZmyNa
NsGbRCNGSAsrZdoiH4ldyzqrAEPcZjBQjIZ0OmotebEhcNCKEY0j73Vmr9+BfbPrlhDNoXiMwspw
wuU6RwaWzlNpFy2ofIgoKRlKHtkxCNJiIl+qjRTz0wRvAygE/nj5el5VJDoMtXy2xUiiMUOlVjFh
hP5c7cCkWCpOXm4PSJfS2XzXPwgc3beihN/IclnmHZVDksXFN7kzApbMZLOJbSy/4waSazBbv97z
M6/poRvNRMWl1mYIijpIMSfHbCkbjR27VeTr/wM44ezHoIP/C8V/7Oos6h3Nt4wEEpZOOhO43Dym
T6BP8o9cwwFRTQpI6JzabSXnWBWyMVhDatJEmPrYi4RwTXVFSTCP0TZnskFtb+jreqexK38IPkiI
UbPIFd68chn9jlluuXpJidFWaMidysI0ems3awTB21+J+0E7ikF2xnhqBiK7ccKJsNDmtg4cbNHq
8IF6QOYIB+6YY51GXU4LPAKiLIAGe47aYTlr7AjpEYMwe53lLPWh9h6yV88SB4UKkjiBwUpmYT1z
WQb3qiBoqDCY5E105Fo99z2VZv0JM8kLPD0XVR7RUui0A3J8lLL4RsuMiox8OrMnRt5j47ZHxwBN
dol6W+xX0DD4pXbxbQAZpRB4r90/FzM9kSqD2pyanY4yaAzJRVvVUjBOsMzC5ph5gj3z0J4Qo8/h
C9A75ngWbqmDyHngXZRI9xYe4a+a9RJYRl0lugi+shV8JNUVb2kLdTLt8K0eBLRoi/kjRQlZXo84
yqHEkTGfmzlQQKRTgSANfTBhy2XvqPfF8Wqdnp/ZRO7hTWYNJYAt6L7Dn43sIrpKzMWBvfwBrR33
6HfWhxihEsXLA2me8VqN9UpxE4k+VVYxdl5Fvmcrkp4VX34Dou9UAKCdPcHnntJd5CRlyx/CkgH3
7jUX5q0OkR7KuImtqY1nzRd5ceX3+wZAac+CG8hTRG/FGXGcazaR0gSUxgcTeUrFa8Sb4QOVfid+
PgLG7+xChABeTK3NebSejxw2iDl9k5igOPqDW+JqjIfHVjZLZIrL+tIDWX7W01+hQkwefkq0ev6h
FgiNQpc+h8lOVypJH0shmhPKVH9rnxIXRQ1A6pEsvV9pXnoDBhb3P9okM+cM4TMSsZEigMkBlB+f
cdekHwTOJ/gyNlIJO+biQ7C37PdgyKz6/VugPCWuD8FaHS7g0yxc3rdU3AV18rVGQReLPJEFiiu8
dPJNE4S2eZLrrqPT3EhgFYdiEnbmE0ISV7fFC/kcXunhcyUIh6+ym5Gy0ONqkVsrgrY84YaA8Nz6
sDklgD99cVqDPiIU5byaOynlOqMwWnb9EI+yClSdL3VErHEkQQyfB11RgDAYddgACDRLKDjxqzTo
Q9zRgd0UbtoyDl7jGbU+20nDPBH60cqsJ8W1z/0M55MciAQcYRoHcKP44xOmFNfKbx/NU/oo6J86
S3FwPtiOfFY6XL7M6oGUxScv5v+7s4GAtJa2Td3BuAgzwT1re7RSl6knGaH8TzfGO9FcdoP105r0
3o9tT/K4SxHr9LUgQRMvPWKHcePZI2UfcyvxblFYKPbyXpA8sewmUX/TCGdVsNJgaocnVBOTXRsv
hsWDoOuPid3xbxKyjFoFfLL1rya5h8XZS7q5pb6FdkbMAhMdESzyR6ZKwZNrt78CWUFnfyxxeGrN
/HtcpoaPaE9DT0VneoZmQbmovSh+9G2bx5hRTTSoE18CX3x7ucF1E0cZFZC8dFIJLF1lnKvsfHXn
W4BDqq5Gg5cJfAWFHuv84EX3dPFgiBi6jFi2zek97iexL1j4+YZjCo0BxI0FqdumsI6UtFJ/N/54
RdkStIXZzpFuaIynHF0Rt+s+2ozmhpJO67zLqBfrJp8IeBfN2FXFHpoLXEe8ODYUQLuKRXrTS0XH
T8dg7vMoHSs3fPKlptDalhvfSEnx993AG3mRHASwo0W9TuCPIos1jpebGpSh7C7ROuqcmj6D1Y27
o9SXCNHJWqxx2XF+pO9ufpjMvj5yJufKSTUta356UX5hrmQLcHcdvFJEnPGAhh5iybtbhGaAH7Yu
4KW4S/xVph7y/lZM7YqQPAC36aV2g9it9DivoPU2MX2ZsjF4xbBBVVqQw/ATA0TrU1SD6gxD23I7
XYhx7rVk/j/hLjWznTIYco9ffIsFhNlVhglBR2Q/pxQCkeGeb+0CCDgHg8sB+vrkLSk80w8PRl7K
xRhL6vZa6aPUaPA9WLFGLz2k/MDeemeb8POTxW4scPtnGJMyd2Ckw5ZELvhhnTStF3gufNya9evz
eIBtfB/lPwLu8pSq93Zrv42rQxopEpeAUT/U1OluS1z3rFJ8IINE4fzcykn9C2sIfGE/5f59ZLyd
uWCm1m7N+ICwkSJteJCTtblnW2rlfxco61Owhl+YtCQiSj6EOFQCZsOIk9rEBd4+o/E9/pZCeeXk
Sg5hLaKa2cpscWZ1miV3TIvRqMRAFboa+f3IzKZTeF2sa+GtMvHUIUAInIMEdZZqEyanF5kCjxXI
xULFN58JuV+Bxcpgt1FvRI3YFmaT5bBBH2/nt9qjw6PRSUNuTQ8S77cHT8Nm2klmwibA2DDGYRxR
3K2ParkShESpm4LeKZzcvIA7vFhMM+odA8StKmMySC4vbrgPsLKNpsFXUyTdhs5su8k/oZDqYgNw
osdaacqgdPFeJb8TIQQ2it6EGDXJlHaXh8J/ZogQmDyTK2S2d2fDQLPgbC7eGmPdC/bTgHGQ62ce
hROcOn63/yTFbzsP9ld1/wFcfjc1j+tz33389+jOnyzK9lpLUHmGiHE3b2igbzM9weMKc93LKBnz
eTEv8/MpR/363f/6DtB9RGaaECO6pBZbgOw/NFdH4WHlD1RqJ0ICHkyRu4ijjm1zk8o1EAw0Owwo
m0Euvvxw86noxHhk4nV6nteYXjZfFstTyNUOPkFQXJrfvNhraHQVLpYoEkjIgEtRNhu81I0vTVKz
g1qtvwoWeTE5h8ZgZPPdxMOWiER0HU5qENozBL8y+IXjLCNj4m+uobqmJTPAL1OK/5lKeVA0fgnD
qWkafYUFYX9Bp50wm3RS815EaMhjvYUNxPvAD2ntYaYKiqlnzpugLn1YqPjSQnahnxtEMQHf4H8g
FrLeIXfaq4KCKE3SSGetB3czW2gOn1RkPmRsclpTCBmr2ua0ZxaMXZgLA5Fv1Ne3HDoAJJGCR29u
NX4Vc5y7oDHjZNEqyRh8QohSDgSzbKdQxpoCoZ1xaReM2IzT66kQpkjOiUC+88GB/wDzZb//QeLg
ESMjkpIKb341QuA1obuWGn/R8GbfK4zNk+dW+DbZTXe0ZZdKPQMgfWOY01a7w/cd/I5YV3qnzsEk
++8ufxKHY1DLcxM4K9ORv1Za61t2XLR+E1Rv7meT1876bN7THBnl1dMFbu8aPm9+AVypKM/hxCj2
Z4W0PEbkpOgJpnY6YDWKOzSDJcC2IeGRy4nU4OjYwRTOqMlkT/nCqt0zYcuh21OE9PfKdXhfSxOZ
pAmc1mQy3eWFTT4YS34gdEeVRnaxnJyECLJSn0NVSeS4miTb7763uQLptsMlhFAmSTgmDjDuh7Wd
ZWIAsKQa328ZrJJbJkN4sA/ppBKOoGXzTdNaA208M+x7At9A14tXLXgfGw7+g4ZiUd7Ow+5k0lX7
KIjt0jH0rIp5QrJjotii/kKlXaWVDNt+6yXpQ7EsXKaxbFAuOQ/tXT2qZV7SiyC9sGG1N+Jvwa25
PLNLJX9aXXlieqJwrC/KZFLy+ip6//4xYrzBzbcWzX9b17rHQKFPhQEiAe1WWXwN2Xp58sVQbIdF
+/lTKJ7w61P1Nv+Bc384WMvf9ezX8gMcZ+STyHWl0cdFLmf89w4ihiZH2bAQ4A/62foJEBFvu1sk
onItts3G5nLcV4j9qyndrqheDiBGCBHyawtf+c2R3nRsdZPiLW2Mr8JH0NxXyezRNlcPgJnmXbHb
DUDHaE7UmLx+RB4rWlN4P1Qe9BunKwGY9Q/bjtMGWolALUDz4lkDxM+qF/v34AZ1UwIbsCIcFJrr
c+dQ7fbN98lu8DXsy7TKxMS4H+RxXS6B3x77MLGaNYMacBz6xNKhMUGPOetnh73CFtuaAqMWexyT
xj+dDpygD5LpBWfb/yB727cPZ5sRgP2ATqIIVBvEIxM27ZhQyptGdD+aYZZQEK5PwPrV+f0YuShq
lzILJ8jN46tCcqcmRHo78TKQqE2kShrz3Mczk38vBxBoJYLKY5E//ZxwI+jdTqsDfr4WkjnpBn1W
veaU2WXj+ZBrFrdNvdBuuUsGR+QDPgKFsdv+DeTEAedMKTT2JCl4aUMmpleQzSoT/97tRp++f4rT
aMKxXVRvDaCi5oPS23qe6lMB7YR0VPdc4+frkygmkFhChlo/3CvaIVrcrRwMLmkqCHNIxMRGW74B
+bOBuDtC7aQQUweHgZzjJ63f+7p/A+kE4st5G0rQddTD2+OubQMTGMTQNjx1Pf6ksBh+qcpl6qKS
lYkugC8jKtCtERcTMzdywq7L4lfOQdR3/UVmSi2gDwz8dYSncPjeRK38q8BA7CbS+0G0r1iqtKie
Zw+NkMGOJM55JTNTOzVeMC7+XW/R2VGsG0huWs5V7UFa5pA8+X3g1riD8kZO9ZXJPSPPxtq9bgkw
xUOYk9yBnM5ZnE+fy5Ly5TPrMhS//QNG1slzwcvG1gFo3h1fcz5c1IFPjgVHKRSjPtzh+k5NbPfK
SmVisNP9ETGfe3Bd6rP0KSn7U2lKwdgPT1hloRGnoUAUBiH5wLp335SmUOcFzTWASGwX5+p2DjUh
VztXDLHlKqdgKmGcv6eDOuqcgA4t5gIk7JtsyVe3ZXWSEiy1VZxSkqHMWU3CIN7yEB1/3b39Vmf0
aE8BMrvsLCY0cys78Bea8t9pXP7yRg0ArZtbjlL6bNi2skg//JA+6ujWRdmQb+B9rfBR/g1g/mOw
XDcyUtVlynT0cOxSi1JnIGqktPnFnO8KjAz71JfPdO3D/igELFqI+WkmAxa/0vRl+QrEkccJz8BA
7LJKUwNo5GMzxQHpmC8TWBs9Yd19rUgwURlxfUcv71IfYke0LxszrxfTH+jbFQT0avEzj3c6lTK1
PAGuext36d5lc6w6flGPPMlZ7LeqIEOw7LTLdMzTgIDurUGfsxemRUfUe7pHlnlPTTJpxJhkhavw
B5x2uNLEt/bFCTj+xccdXJQ/7Qdx6btVFGekzkziUs64ZXhirLl8ijFyHWsR/aUTzwgHiojNJ144
p0Py8teYejKW7lY4vmyqxBGQ8Kw3KCusmyl+kplsPg+Ln409JZR+0Ug5TNpKpzkTYvhzmCELxyYu
Gz2XYbWvaWjfPSqKJ0FpSDHht1HxnwXWv4OhUMdtO8IIesV96l6YvhQcg4jdCKpyJsud2utV7dcJ
qtopx5rQ7LEmqiULLJaA6MrTOX5X4G0th8h3cU1D31as7RNyEzwqpCgRZyY+e3SqtebgA1n0nHl8
qlS4Tc/sH+YdBtEOYOm/5TiqCi5QUinoULz3XOPdeKyeMEebuVCHpv2BMaROC1hTzlV0RjzTdEz6
g0jzmh3N57rcaFzpvSkmpSi1czqmbK01AMGWsJSUuIWxStrBMz9HRIWySeF1RpVDSA0iNdJpxmwQ
TuqzdVjx96yejV2wBzJ6siS1aZaARPPn3zSDS44aUTErP56GG7fdvKRcf7SF8AlNm/AmpG3RFm4H
rkuTMdWhqRP90hzHVAr6FX8nVC/ilDX+59yttADDbcQniJynrLhRQI53HDmdtB3HVSwVyN5moA6/
D/SgmD9RhsJYva5jcSmEcvtcyLfF6hncxGG6pVyWbVhNNyHb/vKyuN8jHbpiJwfA0u/ARgBLrldS
jgOXEvms5rW95kWUKbMAU/4y6+ZqWwkc+BgbwWn0dyFvIA7ZlsQv2/wohM+IQuvXxR9RitUz4iM/
M+OlrfX56c8PdZLuOxMVUshaBoRU5Oq5bnfuFzpDVAG6dvMV9gyrOlNoRul4stZC2MvQRJvxiWZ6
aD4+w9uyS4gqh0RDv9aAYPNrH2042ALSH4ZHDYcK3Ee8O0WOT+o96KpgutJhmhYMu759AVL4gCfb
lCySxyroLuz2Hqq/Dg3FcimEjp1W6Ny8GNLB+B+80WLO/JyMIHtkdz5uiP9WTDGdPUA4GFF0jr7J
WqkQSGsGi8BE5WqepDoNRAPExBPf/GaRPja9t/KRjAqqk2/roRr38I2cGPt0RkwH54opfqwFUgob
19UgKz8NY95tY7Hmz3EDQB2h1jTN7Bvaip/lEEXmhrdYJK2AxAK8YyjuTvWR8Tp6kOMegZm8Y/7k
RaPagTV0mysajCqN6cjBJG0d87KovPUqX2FSwzLHooURQhSQ/ScC/f1+6TZWkThbjhidrMNwp8ta
cd23517FIti5klLppwC0zEWHnZ4qYpvaLxXwhLIs6RN9TqSnnaMPkZBfi9Qo9G8ftx7jVsHPAs6K
JQCw86L2sVPtaluJ9qt5KtnUALWFH4NYk9u4iZVDdLzJwNH0RuCogBWyNwM0srUy/aYLxrad6ena
u1aUyCLE0OFHL74A7NaQ6XizsBl7fHujl0sOXdfEbzwrqlj8MhFnRiyzXKcSBUTFYQ3+9v4Iv5XR
4HVqdMxIFc9R4BMwvt6bJiQgZof48f90mwsVhIfrEn8immrGCHd7cOWuPB2yvtHOLhBgP5NcrJ9N
aFMKLgEiYyXGnYGsvx/AiqLK4KhBirzxHxHkjwCkIIa/ZQNCERzCcHC+cTSiT1ZSnWScM6XfHtAD
rBAQi/PVlbIdZPBI38Zw4k7aBhOJKECFBVcKSfv5x4fdYO475TeN+xBLRHCwCGy1AfqfyP6DNYqr
QtjaUHPxR8AWIA9OjoHpjubx5qVst+IUlS9sTPa2Ag7G4siswFnmhL9Iv0N4afSRZ2rfcu6/mAqH
wgsz6qv6ao+iEY3WypQ+TgJuNk3H8rTdJRb3adu7VM40aCeszF6eN823cJyvHY+P9xf2yiLi/WPA
A/4aHgvd1HEOWKzkQvqpLN4gHLqtYqf7EzK5gW1d7mhMqIXEOKFsmRFScGdj3jyNwJmd/i0z1ub0
WUvEEch9fWt8MNMEIUBxe8mMPNrmAE1if+nAU/rDek/Zy7+R8GXITdjwWRR1WzjkAXeAP2HLwXzY
Yxbwtje2/+VrUd4SirSBNb5MkUUPcTqbx6IiAGqIL3wEuwXXssqeJac2YxgDfbe6pjb1uQ837+kU
N5t22yKLGm0/3Rj8AfNF+TXL2TuCQDfUQfg6oaLSbD2rMSYS5RWvlD8Dvydi7pcBd+VQ9Run+pX9
0IBeZvNmCrGsVCWi/WSJY0YbF8azqY/bM/5jPnKSBxtdD+LKmSxEqJyhIAXIfBzibWc0/YVfmPf6
1fgINuNbBkvBBTouBYOa4BGt7g0yza+5tEbhAqmGaO2vhZJ86A/+hAPQhrKOVfXECYpNrdiU+QnJ
ec4f+MtTgr7FV+F0ZBkudWP3Ut3xhKOLQh6xhX7vQHTP/LNMQwuO4hrYlmRBSJwc/6p+BydTE48n
3X1jZCeO+ADK6n0r+gocG1Cn6JtbXOp68oWHjoyCSBRCYG1BSM4ev+ceDMpmIjA/gWVdmbSPex3c
fJ6CquGyp9JSjMumZEY5ctS92T58xKJMhkDw+8tuXOsTMcZ1j7lIxwlxkYIqRKs4yXmoxwiNufMt
Ok4NdPTyX4QPXuJQe79qyX5JXrka0dnQ4M0c5toUwXMhGGhPn7mfDnykJFHN/WT3DgdataByuzZZ
JUKyKUZjPkZ0MkfF6GziHLam5zTbqFgeXSwiOD4O/BkGRAT+SURTuhFOvcFO3rwCO1tkxvDhPw3L
IA7/v/SDfl9D0x3aG2NRJ9UqjCOnccIGZc8rKOtsIAGHS/pjaVOsojrftY8CaNfuISIs56M0mgDz
KrrldlsAzI0uGHJ+tFlQt1ng9Fs+AgLaBIJaRcfDUFeoljGpK8VCib+ByPn0jHKy3IXuFjYz+oCi
wx3l6uhwtYXVj+G0mI7HwKonHsrTXupSKxHb5Gh3gOsxrafah2Ze3vz29TjO9saWSWSS3xM4KI3O
cqVTslScZjzWte3VvAfQkahHf629KFtnM+YjIUZqc1Q1Rj0GPOBoNX0oJWn7jKM7PgzUUtAfwF27
ihAYYMvJIPalFTlAqBCLdIb4oIPzs3t0sFgDzjv5TLTQvCXFrMdpKdUnayR2GfQxUW5TWqY0SZaI
0s1Zvfw2FMaGWyLxXL9h45CDkYpzcH8+WL/cwz8udjutHli32otzhhUkrrtX+pUnaQH0L13t4BRO
CeTVOEb43zhVbpqlSYv6aHHDAOq4mEU94HGy4Yq7SbA4M+Z7l3FSW5Ed1VbraONrq/TI84cG2tSR
JGdiHzrbse/RWS2h08GwWCblCugEKMARcYvEdSL8uF60W9mv6sWCEXvpoPB8YtrZs59S0au7PqK+
CJLbQC5mR3cx+Y4eEwvWS4/nlwMh2eM8ZyBkuxcc34Oq25kTFVdwShq6UQIg3s/iupTGfqR9Q8Pk
2X3puWDsneJb2UniT+pALS8j9vM6cnSZFfHKJoT8PEsAsyFQHtW7F1fp05EJB4v4XQhu2KNr3o8K
R8wJnbaO39/o9gCqBH8rvsy5QJFyE2OoQWP/E+KZoxpOrxkvfq71IoY/DRjO3eSSFo5QTWUO9+M9
FjmZ023q/0x0z7++1auftVTJjxr27mss/QTV8IbP4t/+sLuuhecCnjvV2vePy6g1OU6PlTilmGAR
szpBuvKx2oSCCMo4SnwvnzjIh7xnJ3ig8REd7w/Tr8kVJTWczukkGDl9nr3PEBex1tQV0LkbGrl6
VABkogh042xRyyJ1WsnhkQ3P1Eu0sXYnYCAkK7moGzddl7zaxiGlEKnFPXEDBnFZT8qw3EQMvJUH
kVKwq1rAD+XLTtBrRaK/M21cwuwSWLsnwP0MS7e7SVakbFwzhrhjO1TB6NiBMaA70JZVMcINBN1u
QUTwbBKLgpeQFoYEcKAfNOY3rY190SQ+Da2m5ngMB4/y4Is2RTeVC7Nxz6dsbDzWl2B6JMqBCEMP
78zd0wj9a62BG5QLZfKeZrRhcNVbOhkYuaktAkE2CVuJ7ANfH5G321j20qrtLDR1n89YF5C3o0l8
wlILHHllFIdkn/Tpex9o+IfxsgLvatIaoWBW80jy8gAq4cL/GbvSKUK4qWRREO2w/ubywVvWApBl
kTnga4AdmkuFMynIIQMKFm9ooKZESk1Z8GMiRYnv/Rip0go/U3lSgUIw9BnBgUPxDexngmOk+m2T
0JOEKDPueDWiCIKI0v3+ixHZ1j+6i083RsafsKg7qkKHBr/nYliGxSOJe7Mx953DGkJkSe8r2iZA
2a6rIlp1KWrNDRdNmxZjiHnoEOjWyAFDc8jZcl0bsu7aJa1Q49Z6G1dJ7vIQFl3pVal8zAbwPlPK
nOxYVgUF5e6nHACNDhQbRodg1zbVB/Dtlve+Bhb2t8mt6tT89A2QLPYq1patQJS5zNkMAVPzeDRr
f/zH6zyhIQwGlo0fFhmaaePWlMfH5xjs2QFy5VBBbA3drtXAMu4skY6MV/znRnPIECyaDIuUEpZl
xsdvo+1BQ8LfqFOKOuvNvMqfNgM/tCYn6uXNBsPIqF9Rv7Orok+q2LmHFUOSe2PKn0JufTijA5Aq
U80y+fz8oFpcC3K0hDsMpz64LKB3C3LUisvrxTKyzyyDIy7QNlxnAs9gjEhFz1gpJUH2YN84GC7w
wIDo4k3MmMpODQt1HfdZByEXEflPwrBtvPjK+MrSvxUzRD9EU/VCN5pL9bppdDPbl7s/wk7m6j8b
NVTy3tiLLCPviqRCGWr8yYGSbYgtYOwXV9KVhQfgOv5jdqfmuImAianhwhWlIHjmF1nBk6DdTXqk
wKttCtuH9sS5DpkpElXi4uAUHQmPr3O6blf6DPtbHs0WYK4/Nk5NWMygDFjxdgDP1Kt5QCKf4XVe
dj58ym8WVNgJaAiBfsPGXDr4axTIdnK2kHFaXCErFlGgrJO1lJXEjrFmlHEgtb1A8CKp2Auuq1Zh
Au0IKM0ws73h+kALv4hmXOCTe2YSWayZ9CsfyAxAlRjLkrqQsjPgGg1NSABET+byeYdTpE21GgNr
g5/Gm/PWgvzokmMn+GULERU+KzFl30viHcdKnsRcjPwJEdP7ItD9gY7qJgvefvYzQiRvIquNo1tc
0fmBXAjlQrBT3siv6MVGWL2gyR/YkJ4U7ks7znSwxV1c/r39AzH1yFXQzN/sUgGX/rnwMl9uidST
A+x0PJvcTyRy8Vb1i7evvs/4OsDvW6Tup05ATY48KlOuJEbZsjQP0U4Avz14s5TiK+yJJHTF+1h5
fIQJwUDrsEif4Lmg8RJoPnZb4xxpNxJ9uM81trdWpcaVPqOiIXVmoC2Znq0e2Zl5SRWoSHBa1Olx
4v3iRmhHCUmt6+kmG0hwvYkjfbvBVgTwEk09PuMw4zmXUW3MlO51N3RJ8zlVnNYsjcFH2XF0yDWt
HsiIktQ1etGfxPr2VDdwdNbUyD9X3I9G97AbxNyhDMtbqVZKqgCsXvT4+u4RXRsZO+QN++wkp2Kq
/Cbs7Rvqb+KfBS5kyN+id6B98busPEl/GHw52fgQrCJINzS1Fpzgsbrq6+xm2VspEgFdLxv3oEzk
b1oC5VmCVmtTq/BSuRIkzabL8BCejfyTcVKbqvq2L9pB/Efc8vEyYr/t0qhmiNakg3/CCmfjDY4P
v7LPKU1s1OMSyUMNQFKvZB5tVflba8FbDIr8cC7uyIGYs+ciwlQHZNrTza/oBPuQ+w72Kg2nWtuS
L3V0rZ04mRyb6UF1ys0jkNsptgX9WSDBTo980fGlJhak0YN0lQrcd40LiPW5IR/JrMPsnySwip84
04MHmFunII7Yp0knlQIE+o/fSmSLSuobq5HQECLglowZABRgLJUr8HKy58So0FCWqKvezxsN40MA
Yt2vb/Se3CisBp/bMMi4wUakfjnNswu8gWD+oKJxYxHliSex6OPTxfDPGJ7D4IrN3G7B9PcFpJT9
MJbZl5KJ3z7CGgmxBCUr8CagElxmmhD+wOyvljWqjdzDiUMdhyaUCEfBmrMaetU/yx7O0CMcQvmU
Zxx/LRKGewXP6abEGHOc+M+oYu/MgEG33SoRraYwDXJxpVnQRdz+9KPpaY7Qkdi9/Cw0UAX3BOYo
HHkG0wbg9IyPg6PoTylN12HLOfyLudfk9IkGXneBkers8McEiRLDu/11PFzpypXzmZOUl3+znSQU
J40dZ9zV7ZMzHAclLDSdDetmdhOD0mc/ET7NpsoMJTRfeKAkGJ3xDdIhVvs68vGH7H/wvWmgbDHS
GJ7EneJx6P3RUxvFMAq7dmEIamyjY6kAiL9fMdTNb4GQlZ9B6uoPscZqN4fs8LU7LmEucR2k/6vw
ALMRa+5pCpaLdm0lMUwLBThDv9LG5na3NbeQe53rPDi1eM+1C3qXda5y4nji6CYGyPgjI7ckrw6T
CE32ZvytMekSilUof9ET0J/RNZODM/G+/aNHXKeiS3Gci07i6TmV+rP+dw9Q9d3B+ODUZ/fX6Kh+
AcAs0g4U1PieNiggkdRxXI18SZi+/cuHXkV3zu+kYHxlMziJqAcCncUwdZy2aMvFUAnN7u0Nlnul
Y0WSs+iNqgg+E3WgTMVlM6BJwmmH2lWZmzFVE3im8YOX7MajUkB8kvleNlEkwfHOkFA4Ys2UXBaK
E8xCsvK63WeqgBZTeqJSZ+maNGbjq9Vzazcd2kaoBNSyGemP5Idr6nmZGX2hhwl2ClGf/Nk3IYtA
NhHpgHE+lvzp93MO4BGiOXYIVMP0Nag+LfD3d5sTgcdnzox+WpNPSywUONGMixG/9ghLJ/1jIwpr
gxAoXxGCQHYcwxdlwkwji8HV/TAt3REBfUmd7NPX/fqtSeoMfYFg2aVL3rHoPON+fT1b0HUqBlft
W40/K2uo2CfK4MGal25zW7IFD3i+5Z8x+F/sAM2/Dz3gQ1Ip5I7z7wTIQXh0rDjvI8WADAStmZrs
tuhYm+Tj3RyXCxN8SHBklo74YKuLGX5/utNNsz9U22YQfdfXFZi+gSqyy7O6djJi/VNGxDaNT88d
WO8/RDA0MjJ9q2XYE8r7U+MgIVpMLqPUQ2ROtlkJEYMHcJbax3d3LDLASokCmaa5lycsMGveM5MG
POqUYRKQMH5Eb0jZ3huva32Gfdr3AEU61Hj1wS3YOg+A7Y5rMILZ6Nji1TQN8EZgdHDmQtxyVTMU
x3xUckSzWeh785NeWL0jsrNmMo1ZrYSBa8afT3GLE5IyZyrZX81RHLjjPsxvuLS2QWlzCRI3U059
c9rYX7NpRGuSPxGYQQgFvN2B/ihFoczDwNVC8MjpvFcswp5Lr22DlYMj5hiQtM9gCc8LH4HkV++d
PfsQoWCrzG6kqgQNCTNi6S+PnnRB0hFAj1S6wl29IGi0xhE38Cw/+jEOtKhIKG6nu5EQPMopOUJH
hbHpziHBa5ZQ8udsQHZXQQBk10wcM9YqSSg7o9ryBxUXBxb1mSJE2R7aVmps5beNAVF5Gyk+RKIo
yOaFfpXgYBbQ39XZMpbpWefbvXjW7rsP9NejgMCN5rmc7dUCI3f4sgCLAYe6C6BA+RWFU3gQHttJ
vXZ/FJ0aVC+tiYncoXuaPCabX6OYyY6WKtHVwMmvj+6ZaAQzefgnVTnXTo1+c3ReKfysq3zOg/FZ
yEt+6GPyBQie19WXZo9HLfZFjv3TdSY3c+0pgZBH9rYd+R698zbupJX9LQ9o9yI0Fsbb+eHrJBXY
SSgXpIrPmQMFokNfm39c3vHME2UOqj0JT60LbieuK+3GX/enz/A0f+jLyny3u3ZT/r4BKQEwRk1D
PgIV89doDAAsLSSiYNX3ruWFaAJg7sDlpImsgS39aN0EO11HXjeh/75CsTNYgMo1tFFIAUGFHpBz
2bfL+Dg581gTnKXxYF4XnZi1CNnVUafTZtumh9h6haiAlU7FX9AnHyT9ysju39N78wyGAnLMb+np
OtDId/I2nCe+43vbdOOLXj97D+/5dZ8gs6ed9J7KIIw3FrBDcKYrFB1dpVIjnSLCEsn5z2WYxHuQ
I8DUthI8cajhElYndWM8OR4sIZ3ITO1MEqT5qOBKbzMIssR4N1oJtr/PKTPa07H5MVVkln5G+LeZ
1G8YeOYOxbqil/ZvECEBlQSHbVOb0CScuuXVcac23D1XRKR7wi5fxE8eDsR2ZsxJrE9OQPGJlG6c
aicAoJsd9StMXvJC92VVklII4ATdEPAFyZDrrYJNHq4r+tWwxbDv2ZxG/L4inpU0/oxtDIShW/Ys
xb6V0x80SqUJVH8524e/rkY5g4ificg5HLwIU9By6cnSjXxjDrkzYqrhFSmDwm+hxSf4nnKIZ5xl
C2ubaYBayne6FXgzzI+Sk5LBRKpN+23OjLU+5UU/WHnpzyNxlZBQsQs/aYTIXrCEKc7VWkFFLe4D
AJ8d+uvOmdngjYK8YEeKos5ReFzjm31vmFBfcVhJFAQhNuV51n/HDlI/TM3KxOcKWESY0kWU2crD
WwhVzCNIHu/iQVNsWzgxw3GzUpw386L86ZxLuJ1vcgEDJHYnaIVwpNVq5OPbcsCIAjLZbwjxLPnj
EOle5vGkI8wBSqjMSmdwejF8QphkWGbPyL7FRJ5KTfRNF2ZqagF2Dqk66e1f54MgSyQQu9hG80pT
KB0CJSrnL9Hh6p/v4FYyHGlAGKaIa+6Amfvz15fHLjL+O1qwQzw49zVviOgoIgDn5yDDLt1dzYNw
C92tAQdaHXEzVzVvDagjPGCT14MvWDZf3LeAqk+SVVibEGukARCcnt7lRoTacdXhJT8Yb0Bjia47
IBDbxBR6EJphVoPvXazLa11rm4p5qVQUz/cE6+2kFoyFyv2fTPjhjpn7OpB66btoEof2mr7RTt3m
MeIPreAqyjsAYoQwlu5kxUg4wsZWT67e3oZ3Xyo3HrAY5EKmrKylevhBt3N0zQazhGiW0E1fhD5p
qrnQ2GJ5MF84XzQs5M5IMz0WG/YWxIx/tNXaC8TX/mloW4LERDZYlAyEYaB1rTh91hyDDprS5Gbt
r7C/yhbpNTi7/arfXuUVDUPG1wjHKvZ9pKzs61bbQPINXPwKT84cHm+8EDUQ/7Wa2YsHAQ7TY8SM
30+4HSWa9/WYd89glegLwuXCMkxhJLbl1sWxxf5+B0HhLfb93J06sphBuaxNH2gim5U8dLGDOmIg
08oeuBgW9gghNQzU7cE1S3FY+ZzRHwgCov+fHm7YaXoowKKS6ggw+MA1uDIABpno048LAQLYLqte
OnPQGROkjrF9+D+giW6/eud0nS58TRp5gep1oci3lIeatr3WBtQeuupRsVf5EerIykeJFdXmYNcg
c9F8D0RuU3SVbjYqHhIpdBcwX8+sy0/yj/YP7Bj52P+L0IRWaoFZacn1hq6oCKfbDfUUBNM4iJL8
iwl9gBx1GSWl2fYGq215Pi7Dv5JBmK+tgoKzXeWMZ2JNCuLBJfGJqzujlOHvKcqVd/SECLREw2Pv
AwkYmxxRcvSWVcsjo2yDDjc41oIFhy0bY5QjG2MZg4uVLeohxbqQ4sDJfl0IZETiedKc3b8pLXxh
7Vym/rA+cz1lQS4glZOspO0e7I6QAc+RyOLpyC1fHZeKHssrWiXllEZOe5xLnFftIwg4RwfcgVO/
p7so+5OFx3f62/k9LzzU7XWfW+jjeKiQp+qOqjdI13Sf2jMsdXkMwhSFpsEmKKfk59bT2gw521pd
t9tjQbh2yZnpRj2g17kY0eu51aTWiwZam186BCJaGRG4r5od0ZJbOUGizyz6PFWcFUHJUXOyrjN3
r9LZtKr6oBqCnTmAv0YMDQMVUK3+iE6hlKJcwxDk9VC8hZmeourOkW3GI+OGwcYUVieUIjw/MPTf
l5epCLaXGqMCSticIdUPe44vCe+zN1AaBhdWCcWeGXZqoeN//+oM7yNeSpvhJ1KzgxUfBGF9P3bA
vrcGCeQ/asQf65knfBJ4fH6WqB6AK2bjrNI9czyCsvwzh0v8pTNDZf0oGGFZ90jZPA/iblWX3mX4
7J5PUV0E3B8wXiEV7jM5ixRPnMYc8jyTWvLv2uTDcNwEQhJuCfPzsBLNcZHugQAVGZIb1ehrZdDt
Z4btH2YpMq+p8DQzfRtwqqAutiNL3z0A6RZy1saMRKJdXclgfUn83SHoQmHYQq/FDNs0Q8o7KBq8
1zjT6gEgKR3xVplHRW68b53TetNj+qq9ShLWrXa5ZFWwK4A6zWEj/gqAa0MFre2xx74/ey0vx0+A
/9o+cvi9NNO6Jm14Hx7Yx1G2JWe5d6YQW/Vq9wslf670z9a+CkMaIPnlRi80dUaqle+MWg+2YQvV
XSVUznvyUHbX9Hx7N6pOgsocYHIimACEKYTO8tk9mr0h7cuDBKlobFKYr5jpY/9j/u3BoV1JLbOO
X4JluigGCelhXttapV9UrXQXjMIqfSECnZgCKTWTx3Vsi9x3OfiS8cY7Jo54EXtILpkl6nSBxJ9Q
QdWuUk3zQryxDAo/ag64Nx44c6pMcw0UaKWpxbYeHR7xLYVWvHWEtmMivJr6UBugUcrm4KZVv1oB
YKr9rvUYQCZ7EckP/OTmPUPHpak+XoBe48kHzsMiplCyPNtCvovR31Vxvf0ZYOxuvJuvzF2HJmqV
pr9AzkyU0DgRVh9wfGcEE9Iesw9kdxDRUQv4IzJqXS4n1O8RZtPVGPET+j1KHUAQ7bqy+sqrKbh1
aSvQb/PA8e+xouRhsBb+5UCdv9sgmCQV3ec4XasUhPQLhD3SSl9ovuIol/8hz5dsYqFKdOo5Pe84
5epyQtDuqSnxW6VUqVD2WguSs4CZ5I4nboz5xpe0zCmxGJdjAlFOJdcpuYYJCqyXGxxMy6ujK6Q1
g48TBu8fgXMf06rTF4hIetGjCE9tL7bIRzGxxZ7jUFhs1l7cuv60XY3y70TPMKyFoSdiP3Oq56Di
3c5WXJoM/P4MeL7F2TORW1/brIjI21BlltQhOPgUkHDNQ+NtYdgq51sNMzcxdUvMu/Qvwli6hz86
8NPj3tlrzittQ9y3zwN/Ld6G5CCje15eg0teUyZr32gKd9LOcd8Iz4uxNfINwTAjFVt3G76tG2Sm
Azg1tVhqYVFlVl7fxDl3sn2Qcxdhpn8KmXhREgHcKPZxqL70dROyYcDYVFXjW3RmFubZsS74u9+o
GzXza3beQuDXmUHWutoycZxK4/EPZ8wcK3qmYtuCeN9hBT4x2mbDjixp2GfU0nSbq24BvE3KYVZm
MDJ3WE8SVst5/nzMNcJXWZJ/Qxop02uvdiFgqwnHBfpP+e/51TziZ4e8ezwlmVmWtHSTC+/J3EgI
kYzJbM3xRiyWJEvmjAB3AiXpCPGugSWZw3zEYAob7BCX4dqpRZQlDJrcQeNiTHvPYZVJwBtBYXa2
b49PLFD6LOpznXO7ACzVS+3efzB7P+HOvQ9FcR3y6r+dfmJOPwmbhPcqCWXYp4xXK0haOKGTG48S
XriV6f0vlk2P2Ruu8tPw9t5EFNVRkly19awqMUijxo6VagIgpooa0L+TrEEb1aCELXKZSe3XHKEh
hZHbDDI9a0vwbcpA2BxvKW7eNfSYUfFHgpHwoi3iSA8pnaw8CbXreofq1UwL9MN0KSik9m7u9LJy
wG5o74OYPt/Ofsp6+MpPFSf6s+WjHor8uTu+pzgMa/lKWRTC75zIyD9dXE8dJUaPF/dMUA4Qr8A+
Z/0eeSpGW2THlXYyt2uiWVLW2fUU2CrNR1CLrjkoluV6wF7vwBAmBhNXWNbNugjK9YVSpTlGLD55
Vk2oO/zcxzU7ZDPiX8QJH5fFkLJC0bZxG6h+TcRTIOR2Bvy9LoGqRR1EGvsv7INtf+UCGRxmpBbc
hf2EEQJ5Unz+y50bJgtW+XJcb2VUn+5WJxW8tTwN5RB6SFGibdjdfJL3crVeMBNcVOt4GIVFZcAU
BZTFSWpfIi2o0DqdPrYZBzFk4n3kv+Ftbgpm5fayI5DDXQbUhffZAEAMT2ntJirYI8hc2/BL1lnB
BzMj9mPynie3A8vz94nUkJwLmvSai7Qho6C/NgU0buIBXrgNRzwOJ6aXZvwJ0XgCw6zR2dqAaZFW
zKzs3aSsv+oFrSF/7mIba+xR1m51qVHrHOHj8V9hoHhOqxQ2ov/PE95Tq3fyA62VwrolXkIM7dCI
zr4nnO22FMppjhpKzoQoDPmusO27xxE39PsDnGcxg5S/Xb0Ei/EWsQFgTUyghb77DxUG6/25pSRD
+tobAJv4eWIVKW9ORvpxtvVis6ZXjMKByd87ZmoHdfTtHGPuKn1tgINWM2ZLS4B85QXSI3rihIk3
99m78n9U6DvSRLwnK373OB7oIC7xkn4vy51SAqA7Ji6yNV23y9BVgsbi8ZpLlhPZV9hbmjaAOYAd
JXsO6SPGjCfM4PNHXwV7iEzMJv1ZrD2JFjP2+vxrMrfMVyHRUg0DFis25zMbUGHAqD+zHyBMizGg
kXw9zi1gL307HE/yGIXoLdLWY3m/4I8+LFdrXeFvCfJUSkT9TgclZoxsWfMCV1NmwUBN/w0vDjSr
pFuALs0eXJQIoJrfilCgmbc0NjvIYxNjRKXbeeDAt58gweaZZwJirI6LIq9YtaUP01Bs8qHBMv/F
6w01Yv8zWreZ9LCKaQt41QCtxOBT3HZt1AOi57Hicr+RRdxsjHHFDOW1bUUyy7ej966XZniMdlSV
MgtAni0rRqauotJCzAtmdnz7ank+xPSGaAMM33AY6vUJsb8sApu/SSo9dWMT/mAxqw/lzTOh9fCn
Ka5QIiThOfezPZV1YaKLi5RBJXXrzqK0NYsdzprRnzevOaFIXQsu8D/HVTZPqWmwLcm1hVCLoKU6
M168Br6dLVLMuncC/lb8Zn6PCXZ2Ft1poyKVjHZSIVZuAnIsTQPshyIxfK6K2OCyupAF5K0jvbuK
DnJMSkdsemvYL0AnJX3GT/IKdjvUu1svsITYn/PsCrO4qEgIdzprK0VWZ1Sfx1sofaiYzD6kLTce
f33RDUL8u+tAFAD7czw2okvRse+dSWOuDHhPfy9YrzPW5gNW4co2pnxoGDcQxgfCljZoSLcuo32Z
mMED20BSHi02aocPOSk/3Ue5GQ2ecuJGsFMltoO771RaCFnlD3WRf/LxqmpMOO1mdmv0oTcflcdz
sZS4Wd8Gjrids1gjJ7xtdyyKY7WQfaZ/fdjzkzh/+Q4cb51UkQFTHsirADnikJmfGPbkntCq6zVV
kMDY8couPwNUumif/Ez1HdeijLA5gey9Nwnl91B/bJzxR1tPwdhDSL5YNX3YmvrPbyU3BW4ixoE+
QFwvVmba2JYH8J+ARqIa8ovLyhyCJEL4u+nc+TOvg4ptyuIrwfeRIH7dTiQThrg8NZSbQra2/3LC
rXIXZZ5F9MG1uc3AO4kBBKlmQaj3bE7DWlDWwQ5gwTJ8sq1YIILH9b3NdQvo/28f2f3iI1MOxyKg
bx0Dxpu0B3zcG/oen0HKEvvzR8DSTM3wnqJ1LbMpEaIbLIA8u8SxyKvA0YVxiKsI3ChbxEXBLDFd
3FUpPGcOi2supKRhsLUwiQoeWv3Ifd7q81VWST0ITaExSq9CIgfbHxkzXApfHSFO5puyarKvoNo5
IemH88P/iTxs2teEkSvp60DJmShfFadLlUXhOTBwydkr8GbVTAAaFVgUmMbgnNr3E1S+bUY0uje3
s1KJKVbgTXoMjWXN935XwUS62LyNLBd6JyH1CnS5bflUWTyd+zXspTfh3PA0nd4rxNiSOL3uDbFU
FDdszY6BM+okPxmYcQYVDfFZL0c/BfhsQhJAGZIJ5WDB8xIdlRySQ+60Xjv2HUUVJUrvJNJrXQzR
BIAqjQOBb2x/q136sMqEXDrVCDTEil5MsRAqztNcMlsmMq03d8fRFeVdVNCoh7KBYFayW7d+Qdcf
xsYUlHSb0iwOCcO3jk7BuEGljxlds/lXs5OBe0A3yDUL+RBS0jdf0rH3Mi9O6BYNuTm+h9GI4eFh
9gfDKx0wDQ1wFAArvM+3jxD0XvrNLL7SlN8P1fVzbwboqSxU2M8k0brcQhQrrI5t3Jvb/4wRmqn2
6WgtlpZBFb+J1VsTOlv5XQ4d7MiiXPcTzah7JsIp2z/DQ5EBBP9vY9POBEBxGuh8/UWWScMS/Nx+
NUm63rMOsxral0CLbkLFexzRx0ucs176eCL7eCfRWUUe35XPYdJuN4WIbtMi8sNoMUtl4iXMD7zw
ce8IKBUUzHjYtzF3zKR7rwfKOJPc9Cuc8vgFcZY6IW2SWXdQjF2WThXuTbigXd+7tMzoryB66HrO
lVl6xevHgMtAMysVnFP2TP+TLmb7QhVTRruKXz4RUjIU7lXzBdNghei5VkhNe+ZhbjfNPLywXbxK
8Aj4g1CEM01z3r9BnGY96+b3Hc2S1XiHlgCJZ3R/prCzF3Iq91BKwAq/DEwCNkfg3fh+zJIAVFi6
eaG70EHSiuHErjBz2mme7or0AtC428NxcbALEpyoZWv4q+jRUitKadMjWRq80Y5AR41o+VPRoC0Z
6flZ5d2uQTXiXGtVmHND3GJrsIHt2NQjGMHsg3j/kKsvOy5/celJDUNzwUVHnpUXFoWP6bmq9Tzg
Sx0CV2uHX70uCMFlaKkC4xcvyXnUzRhfy0r+LOn0Mp7BhnPQzoPXC9qTQHU3w8NL2ZLHZPjpLQe2
D++LZMZeNX3oEUVoiCwnF4qVx2tJFnPywox5uTBs7IN/nuwWkUlrBjihdcE2irLifwaWvPhtdpQb
p0ipxED+QEFJnmcFje7gBJpAY5jZv+mIvUo+pdZggkQ4Xop0p5se+X7DwGHTxBjjR6UAJ91+kN7x
ydQSctuGdpCDXeFAoPvlf6JzVQ88J3zpFYjkbdgHy7+ycDqIt9wuJZtHKhW5CQ6m9THoC2yG6+cR
YDtwBpXEzYaaPB3TYm6RkXh3N3bzmRiPqBR7eZKBr2YrqVSOQrp/vhVV3C8li05/VNu3whxm2br5
S9Cn0JlkHXC09/kXAPihliAMIoxirxKJKxde8S8JyFjTwaT68EJQ3YUxQ3FoyzMwT53Z5nK6pY0a
AOGuXx0F9zBaVdkX2BznjMy6v/KvZ01WGmBbFKmHRRAletIYLIMGn5cB96MLQVBFCBZoFnWeHrQQ
S5sfW29b3pe3vcXFjpX4IIJCb6b1m3ow9ZOQ9+vrvpnrJHYpRkIQP1qhYDLXpbsf8qtCoOvH8D1Q
Pz9TKOet8Fdw1ynP9BjRrV0zsUKOmu9zZoI0gzSyjwE1k80Sn+MLt92oAIFTw8zWl9DJhQpFMuVF
xVxL9oGxAyNBrix+35e15Anrm34gw5xCUQAp97oQtL2j1emdzJsr+AvWFMtX8k8NVCNqtMmpY5up
keIHVs397RM/3zBKfplryZ1vCe8wMCGLhJQIFcJ+pdNlsUzjPbtLw9hZyWAygmnCGgR2KfQnZM9c
+LkqnjSI8otI1R+iN7NqiSihEjAhZ8IH8fsIghjUK9YjyazEf8AuLf2RX/lS+DYfcv4c+efJLIt4
xconHV7UbhfL9ZXdwmVyjoMMKeoT86wWFjorZZwQSl0dvP4ZG5koeSKpvYZCHtBRUVYj9Ff7wsPU
0gE6kXMzSbqqj0F1lOmxwOQNJOcTHiLOGUxbSrGc7e9hrOk+xBAzB+T9+87BJIwi8Q4cIjhBz2qw
l65dZX0x0ajjySU1A6hpZxCr4St9aeAEkxCAsB/Bzk2fUx9QQ/6hqIlAYg+LZgYX/QAjy8miBwhq
V++ULjPR2xvdUfsVKYfXEdIBu3wee5tSJfIKhjHzQDxGOsZ+O6AaJ2y3K1X79zHtThbZvMwxU+23
as/fLyJZ7LDJnD1GLHgwzj+Vmj2rWyIi9sX79C5jlwlPGaaaEfBholSnFq5kMS+J/sKlTWcO6hLr
pUsnqfoXcqIyrQ2Aya3S84MuNMTnm0XD7BLe+sXSesyQEgkdXA9GVOqggkFPkuyk8OUxDb7ECnAs
E66ZZGit3ahHSd0FZnIi43fBhCxclejycvO0g+uV/4Ivs/iX1zS12Q46OqDg141aL2DwabHDSdaT
4ocX70MFwTAN+s6b4ad7LozhKx4XrGyq6HXvBvIqwmbnwuMVvp4cVfuSeDDTz3D/+9L6lVk9UjrA
FJjZ/bHQ7JWKV5BIJqnF/jJ0N1pMLaxx4EaNLNQWjQCtpf28ksI8ZDg6J92ElMCGKMlFe4ELp7vh
uS5YBSl3lzzF7slV1qGLLSpBG3m495DYuhITTUxFLVZFth/L46KX5L1c6+DK3pVfN3Kily61WOdY
wc6ihmp3uMpCEF/UA9QczOTEirO6vtutjDn6WyI2Jwk4aIRV9iXFPZcKLgXzTPT5BpjxLQkfD6Ex
i+1jMXQfHjob8tUgKnBcunABQ0luZc7bJc98NwTXLiz4el48wIQQPgVauC2FK1Doo2Xn5D8EMIDO
REbcZ4mA2QMTOC8CN9SoGVPNvlgemzOfMLkggjEP07KXgpSirJ30yjk8gSDqCVVwFIetWY82r9ca
ACSfWOThB0E5LAO5TG7pdfRDq3+gPgfkZFK1lwle8W2Fz9qc9JL5bMJypuCAEabAgTg7wJN6sWAV
SfBFuT6GeNAh2pVkaPknuf2kLpYTl0anAZq7fZQXtUVVyskeptZatwb8DXlxe22gHcvGJCPRmqDo
Vx94mbfQILbHi4KsEgfHsFSTOMed6azdKzUGv7M0cAmzt3PXZLgsCv8BLfvT6N6WgeRkBkQbV98y
xA6KnyyElITh3jcZH1vGVlOCMHv2a+l4eloMWLGpcfNMmOJjUT8DzS3FLHHyLfxGgiRZp6OUr2uv
ECDoHQZ9PeWxkGiA5owzhMl/FqyrBsbtWIMq9RR3PvDo02zBlk9jfzw3J1DcrdWDwzZNW3uTFjt+
xEyzn2rbniZ/idxdiZP1U8KQQqzDGrSUI1eV6WlhiDQjuPiQfDWJP5BC7gHFbyIcaSkBGKZjBTDA
an7wAskb+rdHCPJS+klXSXGGGx38eRJ9JupRMLawQE1b6dOtMHcas/1tVUXIxEENuuVwEBVanqS1
O8rmSNHXdgyBhryHkY8IFwzqKocJM72cW59N/IWhsA1Ol/wK+Tnlv/PPbIS3yNdvpmAE/3l1PZVc
89zGKzn/XPCyg2x1lc/TjloAYBjvpG9MVRGm4wxHGT3TUJ00BiJm7es8OQ8TB87yVZtgYKUtFqye
rgF/l8kR4vLoMrsf20H3cfJAxGnmym27IJDR/L4tSj5w8174+OlZ+fx9wSO+hhUIliWq8Zb73UXb
jAYcmaD43ot3DYgJWwfc2+fADlsOyBX3LN1GXD4fbcv75xj+UZkH7Tz2G/DnxVod2at1NO6Y8Zo6
PMe/g6sqrTgFA6mUrz7pbYzOhMLPjNScNenz28BrHiNoqh2Ya6054UAooEFayK1UNfqW4mB6z0m2
OLp4DCKJnaw6zV/fdxnlVeYhe19C0GmBb7pDQXLcxOQwbtxFpyNnRXfB23tC6uPE6Aozkoa9bD+J
+FO4RC0IIt88KUa3BomGKfWQxPOTRiWQQnHd7RieVFTQ3oMSy1R5T++qXs4jWRfoTtO6TAL82iBQ
TGxnDp9CYLW3WIg2a7VQu35qeszzFzL3JolxDG2y1QwZIqhwhzpMEy+j91Y4RM6kPNqqTyTXFpwx
HCU6yVocn1KgoYrrUFZBjcNzf0KZkeiKlMxxGlx2Udl9UOMyu0hMn6g/JDfO+yFrW+VYc3ObVsXr
FR3JyO7R3WppSIK5c6xxpCiDNnTYt1DnchxsmsQvjM+RrAJUVxn3EobWUFwnBoCEOubAYo2kAMpw
2K2npMrfOAlm3rrl+2kvIPu+SHNSIwuBGme2vUiz+s8aVttiUKwSfU++OzFtC+nr85WpIl/1b1TA
allPC5zERs+fWdnLLYWZk9tfrFBXwvg4g4oHVeF46dEaRed7EkbQiAVhTWaxI2tLAW3fS884xs3N
N1/M19VmIuIFpGyiduBzCtDTqUSrS4kS9ui4aeQnhbVMFDVeikv1NjL2kCDC7F8h/81Be2IijhSO
2ShTt6cXLLvxMedNBGQjIH2KOhGaNQGBcDhKr+aYEWIoYoOTzYWFJ2DZ6rVeYQuk56BF7wolSPst
U2JUet6BNhnFecJpKYHHqg04uTksuqFaQWI1vKHS3oQygVYggCm10cPn7x9UB5hkhP97Kspds+a7
e3lol5q5M/cgP+MqzYZHFWxYIUnHYR8ssYR+PiYUAkVe0tRWVk5chPyM2D/7EjaGxKsl/rkbKmxi
Ke1grPSOZy44WWlCnFDI4mm75ohJw+m5PLjS6SDNsmtFoIhMt1igoDlfP9gNORHYHtucY5QWV721
gA8vz9bJmhpKV99dsy1qJO62SipJ7qcozwRgNmRCsux7HA56z5HgdCwbmN0hKoZ/FcRmG1iKIXkT
hfOqR1kJIQ3TBkBrX7CmWgUAw4YfIlr/6cKGvxdzAHBuNQGxEAomb4c3cnUqfuAmRdYEmoGdaGLp
GdVnjEdFAT/dtm8ps1ZklTfB29GYeC+wgj9i8rlvTcYtM+Pz8XqKG2BupjHWNp8wJ8W9a0Tnzv5J
Qvojz67zghY47j0AeI1Y6jPbIrg1Wc+1MVG8BfM1qo8nk/2KZ9JkhyswzqtmsIYR3HPahRSAiFi4
qpi1PGr7Spt/werXE2vvKsqQj/DF/SfKm27rLtYPupmVAqjtmCNmxFgDfdwUgV/T3/rkbUU8N/e/
7JUcaZdtY/JV7HWS3v1wSBDVfMsKQuaVODQbfA0HRGVaEmR4+cNcyAghjpOJ9cyfTLMGRFD4axge
68XqKu7ZYDMIZ+yL0MYGu01d/fhpouWyvehTMa9tsRTqi9XiztUZmZDjkNR3CVaHXRl46FLBPctt
zhSnbzfKExY3gqkG7oOR+AVFo7NimvTejblud42TAs7Pp4Rp4KwbHPi6YyCuWDIDV2n4OK0Itsvq
3zSI/5eNqPOJva0S3Y4AbtEqQxYJJ3WkhrueO7a815l9dJ1LqGOlpRcNT8rTq5vjUNV7DWWqSDah
xHAyhGb1suybOgKsaxVVtJyR910RHz7mIiJENtp70sXgU8gQmieZU2DnGQIV8e3yJsG+UG0zasxa
0nhUr6xh/PGE7+HuBpiXyVj8rYiGZ/njTp5JYM5Duh9inTihNoazTINPQnwmf9QIlPjCWglq6WDU
+FUkGy6WWRR6tqpa4wBNFsywohUbcFkbtQBxDNeRespl+FI+EQwEw7SP42yx9ju6QHLjLEqjRYfW
b8KX7/MQF3Yi9rC+zqIGKaVDrTkePoAdZ36JH1nNvWrgzS3gzzBmtkjGBAfifwvSjvlh65WYNpN+
ULjwgTmR9tbZvu7ijFGf35QUhYhnpYyJa8zsSKEo5XMRhp7+JwxYinOZH2lAKRIXGuVOcXtABrmV
lv1ICKbmmLJHHKJKlVC8vCICKQJEn9IjzNwfoGWWfVd7T8x5Zek3cvQHnrEOga5qHpFvp3de+yIn
XYAOM9bC4piQ5OlMqU0PsgmQnjRnCmhRqQT0rWAXfW9Gp5z3/jaqD6KuFVGKA4QZ6MHMcvG1nerq
o1WhHdPfG+QrIbJm68hmipEGFLEdOxKGhPfv92r/RkqBSJ5o4t4uUwnxeEsayCikO3DqeKqTunc6
osfvcwICjdHEeVt5z/xRdQeBJCqIPJtUgkGSQUaHq9awpqysB7bHanPeM2TiXGCl3LLRMFF0o5zf
zKy9Hc8P1TvY65Z6iHEzPBAVwYFatKzEx7dKusGEKinsu20E7iYAipB174Fly2mj4iKkQFEFqTub
J60oCOdnTxyqqDw/CTXx4PzrKth2R+QMn/qmixRypXJTBtiALUDvb1xM5o0ZfJgJQtZmkXBy2CJa
TeIRaIJk8RmclstH0PZv9h85AWaWVuaKza3TdynFtMu6OiS0BgYtCTAS2j4kO91BZo2dVVt2A2+G
5AfZSsaUzkGg98HH0mMdaUkbBs0Po/4VjR3C6bKmMoxwqIxLdQ9sPnGPG/hzPllNNBEyUWfBlMsB
VdBDycbxJFg6yh4mGnO68Tv9UiQ5yw+x28xJ1LzyNqDBlxvVjrGuUmkvEPbR/nxDrboOSsudnXYc
8edosdtZZhoqjL2S76DlESU+KoJKdilFLAVGiMRvLXzhHOL9YRtHQHIOh718NslgxQkW8q+SozlY
t0kBV+sD8O4ufxdzm7OUdmCFcAhMsmuIOb2xVMV1ntXCRD5vCRDQwKpyopzWlSQQHXnZ4gcFqDYg
DJob3JlP8MubZvSibprdVatj2ZOC/q7eb2EF0igEK6xump2aFh+LXnClGRGDQPpzhgYdTb6v8yYZ
BTNdjUvvN3vexdYzrNIc6axljAKRaVoA9nH5n2FA75WG4WV6qTJFa97aNgqoBCBy+QnTjkpeTT3N
INyytum+IU728pCJ/94Vs+uWvnborZYdFrR4l4nyVgdllKSV5k6dkCMPARF5j2m4on7dtOOfMGKE
0C9F5vPrMzkfadU5P7LoqFv35/zA+VJg7G7pHQF6Z+azX8SihhJXOMyQroqLmaBEwoUKJEs1RdJ1
zE0QfcVZxg207RTbq2EmSJemAfBS8Nowa5po7ITGk9RYRPJDl1hG7AIGJXUF25nX43tY2OgwxYKR
TqifxkyLPyHb45Max5MjkGyYBdKOvoYZHC/P0Fn4rf8GNUdNGHNjDteF68/GkwxsIccWcz8rWBSw
vwIUuXj+Qx480I5HTIInACgSyk0Bxh3Qa4Urulqy4ZWP0N7hRzW983UD+/eWo/KTCYVsYXhG46Tm
cQyELTJ6o2mfQdxv6diYhnmiB6vkjijIHBukVx8jQHEO9gwpKK2ycOSgYbNkPJFonzxtcRftuMcd
+T4O3SpBUAt2yHcIGUCt1LmP3eRyrVjSsh1G03kgJxKWUjouVgP/620GM6O1GMdNMJD0ZUtcDh/5
if78pGOSxvhrJCByCYRupN9BW3VXLVEPnFoYsEe0XLxdCa2diOR6H7dyUYLsbOcBPKD4zz0Jf9HL
ts2dM1ZpK2sAdGMk6w8spC8vYL6BKiB+Tl2srLk4XW92dn9k6AWIxAMFzaQ/Q1F4K1tx8gbo4Vps
GQycXHshO4BKoPsZB6GfkPoKJwNpWCpf5s+awIsbFoVXWEaDloI6HrBMyXlICJy7xJvLdSqmGuz4
AE8Wzv+2dIGqykoYvSV8OckrTvOPdoZA0FLtKICkFi2B36Rt0gD6LOFlkVmBaUQ2QjKirXCF7IJk
BX4iJh0MIokFFHQHUhFvlY2lDYqGYNi0EIE/rHdPx8l8HcKCdZfKOf7FLPH0iKPPK7EHewwFTwJ5
Hzb4lwZ3OsOUodt14HLskRGXTP0QUTFDR7qnRaRlHFCE4/ntHF0XQcCMuUNu5cggXiv+pVSt2BM2
8Sq3PPGix6L0mGdZciKvP28fI+iRK4p7TS3NM0sxSU5LYTxWK8JakX9W0Q0/NsByP703kEgLbMsS
DLB5MTw83OjtvQGP1O05NzsYaU10FnYbN9u5zZ1O+P+jh8M37OokMBwi8yhekp/0Ubze2W9TTzS6
UsUSjL4rEoTOmqLUUZLT+5dGJybhGhbyyFMjMe3DBYqbISFmSRgMKhvf+zyBAXL1XLDoOLUesAFF
EMXth7TpFNxamGZiY7g6okTkBqG4FjB6p5QWn22YZGJtiFGY3uA/CzcQFfIq073RtkLfsO1wmapd
L/FaOSIl8Kw8wpx+wKT5XSB2l1TRMtR6/GG2Xz9qIVMoyjlTQLhEH8uMCdUMXh83uL3p697Ld6cO
qaQafPPAEbCWLUj46K8JThVEA1Nbq6ZVZ+blkgWtTrzKHCTy9Ap5E2nuFiYlLCHdcu986LNy19YS
J0e/UUaJEdpB8bbd/22YHbHu9YFID+aZw6tT+Qt13B8VjUnldWSNk4qe5vjrdxLxyjb3K2LWvyru
hOZMY8145DNUjmR9wLJ8Vni4FDhVKSb/QOgQoI8+CfNweHGaQm/DhOzldW1C6Sp/zKL8N07OjdLE
fZLsMBuSzI/k0qyViBcV7Q74UehL1IEMwGudCwQm8eVAw85r99NPql6MXlrSeYAD8N83xcqzOWU1
635OUU8CS7tSAWK4xaffsU0Muykpp1PxvMQHETV176wK2H+rMq6Ia4tn/WiQ8lPxEzXM+j9PdprA
HJhZhPWAEmXlhByejYYmmIzXXX9s04zFQIicaYQcl1paw5ut7d35we5dgBFGSvBPtDoTR6GnFFvI
LyPPBGa6cW2Akw4slsguYGnFecbvWwBRgvRsyUS+j1X/rKiHMaxKjStr80BJBCsZxmdiIue2mzRn
DyCtECjMsMMbCvCR2TLt2zs5UOo1vdjjqOuB74IRvH49j8OBEBbHvE2dyB/dMgAkfTrgekM+fw+u
nvBzSDO248IKgXzVSN4MX25ctRJtltpaTuybxct1pQ6c9g5Iowrv1FmiLD+w9+KiOT81v+K4K0rL
TO8TYXeJWnyy3ASbETR7I1nyyuYFswEfbDH4c7yCLVwZvRu+oJX34j7cbpAweHnd5oVreaTmrXDm
2MdIEQ2dZp92uZDGKJh9kakRjW+/6AO9e4YUkjXAtb6sWZfgWdySe2YrsC64rpgG5WgC1w+01VVr
0Gysz+ZvsqVxALio1lyvF3x0ErcI5HW5kGqOrrcENZ9+wylE7QDtkheKWLL2D6octIIT8KjNGJ+Z
npNwnHV8q4bQM8+zDi7hHgpd3D6q9PXheDlAYSxyt2CAgTvB10SUmP7DhPPyVNE5BnFR9hKncDm3
7NTsYM1NqefkZeA00f0IoSciQ8wiUXMpUjyxynfaQ86vTfyDb0UKVqJQFMkhFVL95zj1UMbKW1Jr
qVtPacMmiaq606r9knaMWg/uDoqIGxuIyFukoaZadiZPZHiZTIfzH8WbFZaPfQPTKPOTBOCLJZFn
S1BkhYHQtK4VJf1HM1g9ZVgGwjCl7ssmC7VNfcMga3XrsjvYAB+pHpy/PjCabRmdmyTbMNbImKX/
VB896+++Mrgbv/Xq3vGylGC82MPJ9gVTEa5/Rg8P8B0zREyECREGrIj7ARr2l95uoFdHUmd4AOl2
1EQUms+KFNU5OuZE6eXKCLebFtTwd+elOl3bCs2mlVntqAhj5A9W4QXPX7K/slOXh/9/N1fTIJ4C
B1m1YgRTLYp1Ri2zKpsLfALG/qAJazCQG80w1A82QV0fFJX4boAG4tcUfWeqoaCu1vFqExE7qQii
g0OM5c4MYXjeTXWk169gQ5JO9jWARY0C5zi82sfNmdB/SUxfWmJIvuOaACe4N8zyhrdJNlaKEDSh
u5RZ+YpuP6ZYhXMqrytBFE4mhOx89FkzMHvDEDoHgXY1Rbn28OZKVnaAJTQQcy6Gjql/1qhft3NQ
KcAphr7e5ZAWXKjogKOUvl2Ou4WB+HjGaorjstK+k88N/aDvfxutttwm1js6y1uZ/xh1dIDVFohd
Ji45kCEwrGdyRtYPPIYtu2OhffZ3f+nFcAGrIB2uXrVDERozWxJv2yhTXk6WC9mzBoZg1+MVNt9H
ZwIbqCf3mMd5XwORAyMhY7f6Lc5oUb+8N1jMmr0Nn+AUKTwImtVkA80SsDjRClsIHhVrZcrfvo3C
SfFS6vDZoX6fJv4f5EsEUvonfpyYk55Eedn0/09W0/wHim7n330kEd2uJMJDZQdSDmGIb03ptlM9
+R7UNFATb/EzASlU/IQ8fUK4QvBSxJLTPfnYIDltsDqe9wUOJe+SqHaD/Fz5Pmrzin/xDW00Vq4q
6gTUiNOtndlvYv2lT6U9DEu8kkdvPkMts3NINpD2Iowhzu3IEvsaUS2l8PMxGNHA45ur9HMetX5+
v5C8kNPPwPhnq3fFeAeIaZq90pyIHnTTgoCIdn2ZN7HvtZboiYqA9xhv7uH5s3vpXVpnbKRhh8z5
BYAI8Kr6V/3SJvo564g/999tUgkFp2km4M8okbZscfvMU7mNrPdcSkS2eYVTIBSnmAbY8oSze5at
EjOb4z5xZksRC225OaT0ZSYhJaCX7IOJMWJmNdmueBf7wKRTu5qGCagzEYVJ1Bw/UaKndlSt2f4/
4N3dAHKWulIbV3NPItC24W6i8PdxngLDLHj29igTzu9xpYHk9aJfe4DfosNrxuuEfR0dolEImFgj
L5gABkOTWsmrmKw/U1E2+TscAs5Ipv176rxJ78Qj2r0FJHbExrB1ov84s2xT/Ti4vvrc5nforSi/
utcllWbBjaD0zcDXL2hSDRLz6pjj1rOkoog6lPV4SlUUjpj966+N8Z0AjmoFWZYbR62iS+ng6MjG
Pfm7+k792PRB4tJKvQkOiW0P18ktgu3SJH850jSWyDlLd74qxgiV1yKA0YuUSFdFiHq/pkOcHIgz
RF++8NnvpuPy5gEpcvSEWLGZ4o8ScH7NeAhhvGzAVyaPalwJbF4PY6w5X+2Gg5pzp4aKatYo0+/N
uu6ifwRCHWEKZ0D8M8EvZuNph+/N0uY/+s2ccqBXdiVdnF71lf2OPDbZLfeIq1f9oNYyrAsNRRBg
LLN5qSE5flshiYMjN639Oxqrooade1EbJBEpEbrwTAYVTDP35yOW0m1Z6LPACk9ivovKq1ro8my9
6qqGEBEBL71OV3fp3oBrW5t8gYj2hVDdhRmXK/O3UOiXjYgx8P1BCUAk0psY56ckFScXB4TgKP6O
+Hz32KuArw6Mb0U3y9zFYA8osdXuz7LXb33I1MARINPBxSy5kpuI+lqX1eWtJ88FRnz6Sn4v8uZt
DlrKyGD4VUyVqW81LtS4FAAZhELj396i5BuMNaMl2po4OJbSyXoX34y4hHb8kMSPGR035vBqy6sf
qszQyKP4ulOftxVM9TZJKH7UOh2KBdMX3UY00ZuSnCXApqCLL8rnfhUYKXHfzvdp4HGgTjK+9okp
y1VZCURwUmRGYPogcyjkSW3Vt8kMK4cChRcIwDR1pmRZtfwDtwQ3XBNc5gmCBb+RdnPxZIocRKZ9
1AHJ5H0ni0DEruFA0w2lK2XUEB8enNnS5ZrTZmx9ru27hcYdLwbH4IxY25UnzrhFTtpzRrk7mR07
inVMjNj/BLhbAm0HOv9f8D9Tuh2X23fc785sMBh59HbkG1kZ29pdY2IPbFLvyJgJOLspNteqP6E0
3NVuTViPv+rbCsll5p/rGjTAbs4Un0DsFo2N49WUN9pfuy4k4iEkem5Y0mm8rXLB/4eQDOmdpWvF
dZGALX56GFIMerxAzf8M7Q2FDpeVOA5XAEAEdLkDH/n53OpLQ2idkvkzzcZsq6S25XoH27pYvCy7
+2pkTbwi85GwL+IrzWwGc2oMFD1MlXE7FXasHQugOhUYHGLv5B+6mX4ZR419b0fn81/5UY3RrppH
f251s9AanPPreNKNCDANxZfpWBVz6aJqywkqh8w7Ma9sCU4h+vbILhowXxzCxCBIYyus2oW6zl9i
3ims7hIk2ipmrhmOzDRTVJ32keuJfl3CKAfKB7j5djWN+kA9ot+eCxO+ojPe3uUqsSy5sGOcu975
tHtU9ZDQRC5WXHZ17cU/5iNs6C/JZ9Al9uBfU2OKYShXT9vsHDq/ExU8TmJfJo6Nt+4+vVyRIkIp
K0Gam2ZuHwySeNgSgz2ieERfSkxX/zbvrkkbSotC6iny48UUbzpOMh4tAO0yqBSaQJIvaf254RLH
VBt+/4ECjgIm5CLMuSbUrhceAZv3QsfHpoRRFm9E05kbSj1gBI86bl6Idk6mUUFkHGpFmQv5V4t0
vR9AlNxFejmN69OFyifPvFPSwWZDUOPAAhQPE2VSFGqJv9bfAydfpNDBC//SHSfLee0Isr3a+TrJ
dPyX/CRDz2tROoVwX75W1M16s7OKj6sh/4E1Y3k9Si60jGGA13vZUuh6uZD95YqUyuEM2UggxvIz
w5reb9H2QCM7XruQIFLxF7cj4M7O8GTeOMmWdT8r/W+aOCOg6o56T6ydpC41q588ICeyfRSJcjFI
P7wylEWGTfErm/ZN5yossaOzzVrf7eKPmqlp3KT6WfzkDUdr8DHYv8GY8Q9rhgFyUtQxLgOjONZu
5H0PMgRWicb+7yV4++Ed+wojUsG8C344YUFIjB2ASsa9Q3CEO2cz3R43bxYEwTyny+Pmj4tdl8PX
TnNc/U7dhvPzTu0et1WMZEaIEKCW+ARNfcEqzdQwpomZf0W/zEsrr+KdkQ6ibAVPQNEL3FXpr0dT
enuKfLdXzVCbC/zDtFkq63s5HyYmVhrlqsoVJLypZt0SSWge2yQkAbjoaBzrUNF5n2ElQOBMbr/A
KQQ67Vda/XJOdv1QnV+GKvsmEgScOXtfN2WqEQO6R1oIEUBBUKZXZJOVj5s5ejcvWH/NB5IHKTue
Gt2ay7LUYgmwGLCWWfQiet16whBmzLxp8JBD5RB6SebTjxZYBnEbZSnnwkYW5SxhkHmEfQ3E1l/R
IF6gpUV4fXxycas/24Q023hsvxfkLvPi82RxzIC7f0a4xzlKeaMD0eIifn6Mv+DUOhIqp2F69Na2
wyc9pXR64MK6uMUsPlHcUKCdVTnB2kSQ/WKz3xlAEHEBAu2MxX+dTr6XFiXSLADx/wsyrQPGtTdQ
BWtqAYGMPT/U4TaYzShePjpa6O/c5id+P3qt2DODsuB0GYEGSTPPhzPsr5TK9Q0HpfB0oNQHy6qt
s48LKkQKt/WVSu3r3eHWjT5U+tucDB6iEGkaiMoP1e/2blXH4J6DqfnxYtI7gtakgV9TU8u6p/IN
hTmlBq6lLsyb2Nn8IEufbs05pM8GqpDJAzVazGYSawlkyJ5wJdMerKn9Osf0keBe4ZrgvUV4+5De
SMDlcg+66idqHZ6uJrsmKLD1jKXukm31zKDcmWTCxOB/H2+P22WIfNy4Js//P7M0gFvM7FYtlw1F
elbJ5vLvpwamQ8jFboFB+r56qUPT4Y44Ex89YtCjqdWdqbT+Tq9wM4So6LeDHqr8s9UOsAkGQ3wx
Apmoo0i5dlKlZ4PP0muPd0mefxdzeRpUcGdhTkDagwSOykhKD7Q3P5lWimGsehmOm6P8pSGvRt0V
4QT4pXsuXwsAU5xtcOjW0VBvbbzXLfFttsEkBlwfZ1IS40elFkOYV3w7hACOKavPL3yaDNZd7JR0
uRpiTrdpi9Dxj3qqlkC27d2FDAF7opPk/pk3j4KtA8LpfBFDnQPYT4APf8ZekNYV0DzTGt1qDfEP
glt6tLA/mkeQASPrFNciiMHUKwDtZLA8NYIkMwp3HdZLuBGjECElIh/U0xKQGLZLO5jf4+S50y+a
ksVnqZjKXf8O9Tq0f/rREK3o0O/kqDDXRYxbTaILXETkgNGbAwTt4GYvh6PEa4MwpsqwzyOVb/wX
TDA5+LkgtfCtoLYBg+Moy774CQQZggBwE82v4JML0/N6BSOhOPX9jgULForTQbivModAIgiRR/7h
GzJxt3uQj4KhbPGEbdoBBVkCixq1dBZSaX73wD1ZJsud/f+O2e2UYbMtoqtCSIKqn1MMNbEP1RTq
JTVSKaAql8p3NRRQG7Kn2XjTHSJtU47C5bn47otTr6VNeIMEFJdyR5/v8sglhXZm1Wvqi0uu+2Pm
0osJdAITsJgu86z7pVJuYWjTfZXJkF3or6L9nFrSN1bXEJiThKCmBTmrIQRiYSjERSsquBj8H5dF
8TkmXs0s50hcZabGsc1UVfGnAiEELdMkRz8q8AYEc6AIm6EPKOC8+w7ZxmOCZLI6r+J+IRcRq9ql
4ZyeuTfqc+hLV5RXdFuC8xcUyhYVSyK372WR8i0HBvlfCs83wQDKM+ZGOi9HrbW+yYweXH4YeX8V
vWxOQSmHI4spxxLc7UgSUS6jW85rqXqQPg833XCKLP2aqjbCl7/OcEDfWSHAUWea7CQIXcVQPkBc
5DAOoVybsS1Dbfg8ewg/cgXWPr9h3igTvQGgu9JSuhKxhhtC3a7Ly7SXJZk4BJUN7M5j7qkL6Ww5
T8Wu5kTl9kh+3gi8tewOmzIT8dZAhYhDy0e5LKRVO2B44O77xilhCNZA22V68gh3oIBxn+J0RhrD
fLZWqTQ8t/y4BeZgs5G5xv/fNCfRKAUveeQxYejB43+Cz7z/AB9OSE6ywRmDuGFqrljdwcIr58WW
VlRI6JT0ZKzyAQj66iB4Qd/OuMTbhMBfQTpWV3X5NNL2rE+6Rhkffn0v/DxCm07j0ovsus93WJQv
TgNOrrXieoDnIg7abs31SbU60nRdkowKb6oiVmZSGlKAa39vSebPDsGciJ/xhCFkZN0u21Zst6XR
PkgNYVwDBzS+/2umoyLMKwy1NJKode/S7Cxp/0w650rPrN3MNNq0MuxAK2Cvet0/kTXs2HjYXMWU
38O15dGUDaQ/PILqeusUkheWoQIKN+uZUiRazUedCRHxA+tf1hzzOek8ZL4je+LPxatku/P2dD0+
zw2bA6Y1ivPTQBIL4aXnsDEcz1BBWzaSMIbL5kZkRkCVCAm5J7Glex4+k+bCq5odMAYSJ9EZ9yDJ
t26KdG8iw6tixg16HkCx3wkuVHJmnAy6acG48pbkk2dMSrw2f0n+b2te/jYWugNr4Wt4yUwtUGrR
PWi82KCujKhHDX0nGk0/QRyCf30wB4yl8ZX/J2/aG/7er9NBA7D0byb8Haxk1RNQqUTUH2QXzI1Q
g663zn9CHM3YETNDULVKfeQ1UVNKa4ieD4123N1aoMSpy1YkY1UVZ70h7VujdWhS0munDSQD10+3
yIR9+gvar9wKwQRtkcMvJZSSjj4I8xmnZ06LO9KfTfUIsUn9SlZcvNGU3XvZSnoI45T39cx+IgcK
u9T3wuBz9PqDGJtr/Sxv96Rj/tZJljwJhL0jZyGFNzW4PdUgZqULqAcdLcJz3Qm2Mu7Rtb7dCcfQ
eruE3rpK28AOsFtGNVTaBrdohA0vfsXLVKZhSmOZi7WQMu54mSbOrsX93s7QwpcPLdoYAgtVlnZ+
o39n8Xk=
`protect end_protected
