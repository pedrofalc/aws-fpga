`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
JGMSJhNSyyydOIPRsgaEozzMWuwwoChFFCDJE8oxkOCDImPEU0L97uRwBWK2lY+WnkzkiKoXzae9
Ch7LevDp/Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jwDXt+gNeq4mZF8ReUOTkKic+lMBSsrGDOHxmefSAcIkQVGzRhIIeE3QB1xOIH3/sX+yrzQY0TKS
uBvkw3QGeOX2uKDdEF0hsP7FI1shPhHnI/zyJotU5QSL2MFECXJfexptDi3w3DUoAsjpZFPKc5UG
jAZyJMqcSWUGRX19TYM=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bxth2fN2pc/HQFYI/97Ae3NaY6XzAmf5pPTZ/0FCEg6h3hpudOwl0niyd7xUjESC90UIpfkI4GyX
xsP/dtT/5Jes3sAlh3rPzpUqSw3kEuTlm1BJpAA9+j199Ysn7j3yfITq2rPPuo6v9gcJOfenqPZ1
6HlD9lTOxGFFb9V7OdU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nLgm9CGakuzkmfJi7A1Bt6KUvli4wOEdQmJPdOp9JWU7XHwb2T+jkW3d6V2UmDHzne3x/LiIisCM
pIrluZ5Ts2/RDgJOO6dLxKGN/LcoB8HilmrssJPhHlD48sktV0Zi1FdQbjRfP1gtUYw7U0fSeI1K
7UkzEvRqYQ57/yszVtQFkIBALX8IKVG2TLD/uYkDzEqAKa1/EfuOoxJLjK31gNq9lZt2lYbSJTJQ
rxQ2eJSI9BlORSYblqJq/1fb+UiXHK1VLTYCUozsPpM6Dn+56MoOEHwpJ3fuWRBCXObXd5R6ljdm
lQmu5OJ3+5KevsIaMVp4riGmTHGU3fxhRzXO5A==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QtQC2/DhmowIMslQf64mGk2G5yHtPk6bz3HSFR6VV/tcKxXizyTxUIOKpRGqFVF0BubckMLPpE8S
WbBb+CqCLwPMMZmhvEy9sV6ESwot+g0Rmt55kcNxq4jRdw56SAyqOdz0S6ZWsYjzeuBTLUe3pQ95
PtBaoWdj71xs2UyGh2mufMZ5LySM14cMBDz3EFMcAkqYC1KhtU431X7gnfRDKKqBWsg3RZMVCwUK
3Q0I63Zo/joLfgbXDBRRSbYdSldUx7mx6CI/utGOiZVQPzJ7aE6M5xeGgJVE6WdPdYAuAfDlJml1
Cpq4ZQT3XPaIdRa4kKxaocp537Ny9QYuB6abjg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NGIe1cBwuUxuMjweozusv87PtHhsNdQsxDes42AFGecyH5hM8ufaeHBnBQjo53yXsLJQYH38mdLo
PjfgJMJXdgnZVfp0tzw4qhutVLEDbhJRDsqJ1xAW0cSE3+PW0J5eyofktEBsiS0Kj1vUEcdy29W5
Ec5JrBn1pd5PJFQwsM480oR9m6zsPyoZMajeFKcUTzFAZBOBbIsOXPMQIsBOua3zbvHNM+fOzmhl
jQxjf88NZ/BZSo8Ul9GKyOY57WI+tbU7HXdRZzFRbx9Ym+pdk8xa/reaTty3FGH6xCHUwtkBb5GB
0Yli+xBmjb0mVklm9PrqvKjy4XRGlZG11ECs8Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
v1R4IzcVsFroXt0t38Au9wuGzGE5elKFDMoH9IFmjpmt1JZs3FFkqLabp1XThsKrf59a2O8zcovh
txJVl2Xi7nQhkKyi2bxrvfzMp3eODmtml8fSjuKPiGYOuIIWSQBJOSLqyAJwoE7tOHWiFgW0h5Ah
CuvH5aMHb0RY5mt4MSyySXXP4IQaCw0jPvBGa91qSXVI7UB8J1ibt1Fw6Xc1qYHXfjz8C7hKAF5k
hkP1QUe5iSGnYjT2YR02d0XHyKhzzhT9F433Ai6zUOIRMmnGYofmaKCUkE+PID8nGhTNtdH2AHsp
Ilbs6pRHT5jDhtmdvj1xye2WoCWTHAZ8giEmYxYoGnSH2nAIcO0qhc6HXIudQweWGHSxKdwbuDUz
kYpp/4CWcSiFR2oevWlXUJWavYgdok2kSTG7MWWQOf9zxpmuWANOPJW2hEHCMOlbaqfK7/j76wei
LaboHRTEszcydcJEucfN8XSi0Wz9UxyW0HUqf+Bceh/lGy0EnU0imL2pauRPS75U99mPgCBJ2grB
uK6PNjbGWryk6dwGyNFvZRU2NAou0RakUWI4/fFe+xAxwQjz5upbIVekUyUY8b3a8l58YyMs87Mj
/ZmnOcirF2LeICpno4+MPJwi+EofrtCUXCIQCsq0civqrnIDAPq/tvnVkq2ejNh5rBtAtOUa/YKS
6iE3VmnlS57zbowDLsqANqLvWJLTXp+QP3KCcB7HccVj/Z5tdcReFQM+YNnKBnGa2mOZUYOm2DVM
6pz/0cqZRbGpycmg4DWvSLGqxUXlQxSRX9WCvxljUsl8DZ83v4ECfu8IXgd/tz30mULDPvJg130n
mj2hGewTMN//Q9cIB/mrapeU67yCk3c2VhEVshdezHFyvfWAwtq/mhy3afKOOhUMLznr4HEOrSdP
RjK8/kNdJTPKjjwvb4gfftiGvug2SYdDOPQ+uL/jgyRnpqpOwtov47Gp0JSKmNV44OLyZ6bi42z4
BF/Sv3qoGZBRxvooXS9Cc5GqhiuGERGuvVrBEwkMLZUEHn31sYNXMoCP6rFPGQF1oESVz3z5SCzT
F8LYSnoqOwbU4yfmeUh0R+0mkhysBFm8fQH9bnxx8/XIiRP5atlfM5C6Ch3BgFDxHwWUUY/QfWjY
VPuelHl/lrKXCRaOMeXDcyDHrzGRXYtAcwzbILl3t/QRxARUuEX7lgPv2zyVFa1NqdlrJv3DpwHa
nUtk3JXLUYG9Gl+bU2P4nqpIehBLMBeZQ0arSmbG5+5XvRMoCU2oSrNx6/94AwxBh20ZymX8aDnY
XFyh6QHfoB0rsXDeBnnPjzJHaVMzRlx1P4T3WtZEgCAAPEn8zPFMeG3kLguX5xRoXkWAmKW/2Rw1
W5LgRcO1/aiGsa3iizEEBOLpW2DYnqmCjwaTlSqV0+FUq8uo3IhZKqoyyGbYsHYanDMSjW8htuZJ
D7iDrk599hezmIMkur35Tjc4XKS1ujh6E+fREGSFoF3pQqxDL9Yot7vJsMFjYtSKEKTskOa8zkvc
inlhmp8ls4BVz5oHbYMY4Rxo7sHuwT13+h6o41sDYV+NHVfU1ufMpwUi1EA9VEKR5v1ygdv7m398
wDB6P+HAuc+pH/uIbiN+F4YqQmYs/7IeD0FTMOdqJs4KW0iR/WFzVIKJsqiuxH7oEoJ8nsTIxHNQ
xq9h/43Hu4jZqvtYCdimuI9vHZjoduCvqBGStEb0KJEL3tEm7O9iU6pTzoPCaPDBSSTOWmu30o4I
wcQsiOYM7/VM7FPv7gwSMd6863VBK2Glo0IxaDJluuORFfZnWiVfNmUbLT6bJ0i3UfWIM+yMxr/v
j4voYBJ/th3lkLPXYY64oZ8R5UVi8WwFU27JgJ5vpBt86eTbf5nFzmalqOlydQiAXjrIyxM0XcTf
pUncgmWr5GgETpuv6C4dKc8B7Q7toW/Gox5Lxd44aNhi7AGz9Bdc/Y9Hn/rFbMomSmsCsLHXG6m2
oxywvPztn3r9ZUsOU2lvQtBsf9GBkjWuuzkaohOT6z4dN+O+zVRxL218Yu003UA+coz28/o5yYat
nUVfPiL+XF9hhjjoZOi2dOz3vdQUfPU72CoqIdmDF/9nNTFq439GqyYWaZFTZ5LevPb1dLvFkDbb
pn940OPLqLIKn5Y99L2hXwCFRgXgZr3BtnPEONu72YoV3ayQXJip4jWyOH/QZ0Pzh0R+rRXdmcTh
Os01UGBaC66AGmIsIKlwfH3ZIbGiHNGC7JIBYScmxpq/jG6QucQXWBLPYzko9BE2iqgvj/MPloAG
Df9hlNhFhxdr8NDx3cUUI/R1eeakTElcWF0L4RFgAvPQvNQj4A+D7f16yD9yogcOfO+ohbr6h2kU
xvDGNvJgD641cVkpiewLe5qiM2nTnYY2ujLjIgeBXamkXpAIsRhLDusb/0JuxJyXEUvWDba4F1/l
RITcV3r7MQz9TpjZ2ZRqJM3nZ6OJRytEZcjW+5jKnk9JFAC/V0h6RXOBj5XKRXxE2yWVHqTvEaqi
oAKgriXGvEJXRJbXBcrPhapqJuCeK/LlfB5RPrDtEHPKtKzGoIKx7gvu6ShJHhLYPYtHZBZw/E6q
HkRnHO0wNhiO4nLYyVA/dUURqWs18+zGpHRw07xF/Pe52uYw75pqX3sKiPbAJSKP53dJqKRXOJX0
7fmTCEPwLZvaCJw0yswgaE43qp3Q1qiC/XUmq0qEBSJ6UOhI9MW9PjSTb4DfA9QgOmkav1GPF5d3
zy6AkMupC40eBWh+5Zcbrky0giMdYEdTnBAMV15OneX1JdnxHAMwY+jwGiH2gcU5YHHDz7QqV3ke
f0OYZJRsoTkzs81EKP93Q6S/j8+Eg4cmXSjTP2V05DYY7mP5kR7YCs2nzp8ozKVrFW357nt663T+
ulaB/sN1aPT0jneTmv/anzcAQ6uocIWUjWSpZZJqH1kDJTCIWKiQogQ73K7BTcoleUqd2nojSg2W
YNTrykmuVmsv7W5fbm1ZsqMEqSzn6XUKGMEFLF70ots1YEOCdlmoAZzmmq2zv56cO9CbPyrK1hqE
hdW5+jNCjefyjvh/SuNU1YIGyaiolHXCM7pyDWwM2/eSiHjVDYpbnWEFBJnOvq545OiMeuUxzA+4
lRmTqP854amqVIVJ4BAII9ABX7/THZsJgAFFapnWAUJYd/JMf4Tl15u9Nhvj6R/YbRq2P+YFhNsR
WYs9VhsLn2qO8jzfCn7SqEvvMcTSHwo28aJdg/dzHBozFW26Vsj7mkcEyo+tuj2ePeQXoRxNoKlS
Tmdaa9aNgkxLs0mUh/7yBlGm/DH3eBE4oq6vm2BVBg+s/qr2nxKJWvATYnPFPTYd1SR3khoNbLhN
NskKj0YhTsbxDmjbfpeKK9bsmrTKkSpvgRsiFmgXrS8Wv2fJ3wU5xvSvE38ZeuesUaj8++bKlF7z
1P6WzY31RAFo+axl4FJcAY/hOOH7/XAovmaA0S9+3Ve0klsGXxdc7/E45x7NNWhk/9Bd+wmA+KdQ
Jh0b4IiBkZAmvxq+ckA0UYdWeUu6nKjpkxZVeT28rZCpQ71lmW2Vgurj21iXaXCSUUOX3mjSwbkz
o9vfx2GnRT2kX2mCktWwRvt4I75QEgz1Epu9cun5PItuA+ut7rQGTohFcOIi9jNM7Q1OAjBGLQM1
8ZEeK7QsgIeKtsaOvtBXp0V/TH9MrILck8ntmsxZSM3R0PaRMZC+sYhkn2STgZ+t8Mn4K8zbf2oM
E7C2T4SHzotes1kfG2TTNKtU1kdhFQN4j87nUbtKK3OnbCxqIUlP+UFTZxLqAmHFMmU6A5+AkQA3
gT174S6d8UeQRIKIU4ZbMH8L2/hSPDA+Q7riLnz7e6Hf0qnIlefI/wOazvMvfQcJb1Wzi9d/o6N7
RcYX5ckQMxj5PKRFDtA0wAwsjtWwOh+m6QHt+Ynk4aGocaXPyEZVQ/s2Dn4OpZj9sn/onIXrcJ1o
gHr5xP9QG9hqaqaeWdvmkk4VccooLasdNMJZcY8gX3LK9CQMm9mnl2K5E7tqab7aI9aOeKxlT7PT
odODYrSRsBTB7odnYiTyOgNnjMeOyNBBFfhvGN4deusxiDjbvLoGsQYs3TdwjHDu5VnvFke2zU0K
U7+COaDZkrjpGrilz6/gSkoA6SDj9s5VTARyFGM9fw9ovuGXj/fROt8dI33XtWBSns4Qqgj9kLV1
H6SPTPdd/GNh92a4mhb15NCompLsEn3CIj0AngyKYkr8dK21xU2EVEowPAPCYr1/OF1RmKmqHoC6
5TUrs+sd/EPJPb66gZ4oA32GkJFpeZyxuh7tJqlfuCKcw1krASY4cZoz+ww/hbBJX1RBTJGRKPm2
sP2f4znTMpkS0llNB4sbLYv6LVMsqTryJ8DZBL+Fau68zM/07uMA5vAL6wpM9xPtq+9M9CMyKU7U
ry/9+R6XFxroaVyn0Z2LPe0nIIackC12SMbzrn9xiph3wk7a9srGkMSmEUdkcJcm1PfDrc+lhH4C
260aiGRCkzdoRBZVAYBDHfhEiXW78uP7cjPFwIS/2ntEFDMHgAlYnx9mSJcVf7B6CN+wVRebWhYA
D+eyeB+ji66DSYMz5DPwTuvD1ax8FZfSKDE+mW8Eer+qQ/x1quFqDc1MMmL7ZXjcS6K9p6u7Da98
8uG/f5CZa7PJ8PgFUh9jEhq/lF28iwitCNDIB+Mx4LFTbSt4g8sI+VrOx4aWBeA+yqYg/1tOIqqS
BkzRJcLYP7nLnFOYtMADKvtN4mx2u0+Vi2XWQRLFlUF22avUp9PPdWdnXXg07+S9tcqMx6whi7NH
Sn2TtJES/eGxTBt9YXfXU5i+CfMPG0Sl7tsBTvl8RFjdDm3EOdkQwa1VCGF6Cyxl2qCZtXUmVEyq
VG1hJf1nrZ4FFRBOb434VNz2dPM4CdE+1vC9l3cpWvKeHqx0lsfE7T8BDFHfj6bUuCFtI+cPzS8I
Mlvf+9V/TNJqsqGpFTPFyIqPBrjvFQa5/4AGLPWawdMbAwQdVWDbswD+WjOolXbq633V6XXx4R4J
2jHG2NLaEeH2dFRiS4sn8tLDEPcn3N1wUecHBDSG/KX3tytJMjHebNPYlHMy0dvbOMRIWYG22GfX
i5kONn6+ssKvP7WgFfNtd6QjcYnm+M4ysyNaqhRFAPj3MPPQzviv6gygScBRPlgC3ZlwUDYUAtvY
pd1fte3PUrF6+TRhfxrqz0Yba518vnKksTPIi7lR6tvrSI/I/cA7sPhIR3rG8DXu/ZnlD38j3Jye
72lcnhQ+Esj86iZ9P56u7JdyUIOQid6S07dueVUyQTPmOSUX3sZXvK07tz7dR/aUs8yRm2cv+FoK
4xCSUOyy4bDczEdD+C4gfx1MeD2qn/dVNLcJav5AaoCG2qG1hZeXtLLNOYgPqj1YGgazhmYTLz/Q
3oTCjHGcN/+Hteoo8lewqvG5irq7Bqg5Molmril/YZ2UBIGgSzSDT2JypQjn0PYziyvYC4N+h4ao
vKd3B93UChqIxWSgUWc+MVV/61DGbH3RxeZXWAdgRkW8dmWAkaQokPaJgQeEhaV08u0y9BsRLPa8
aiQpxIYO/LBtGvInIcvs5zlOqiUtKg7q9s0yxZVCewDpa8Tq3vVCJsx8THjarJ6WCC+BCQAsXJgy
5ZzCaiF99CyQHYhoDfzOXAwTjHLc07oywm3VeLfY+selEZtNLQdIgzJpiCnImK4nwhHl5LvfG/jA
VDsU3AFOFT1FvvW1hbXPFCTkC2gg8qxrrsqdUfax26+nEGzx4/oCMbIV8Rp8YMK4eCrKhKQdvb4j
iEWvi628qB23XgncGC1DQcAQTA0P/PwTp7cODtJJt4PHOCxZexcPvzGcZ1YwiO20AD26+JYcR/mV
FLHfYSDZWRCWw36gS9djnxqDYEzKyN0RY4u9wvWnckYvvVw28tJUenomaJPFZoh1iyUnyJQfiGGl
WejzuUbA9KICn/klBBlgO+s469wAhKpS/AWi96HHV7o03RjU/Lcv93gbBhG7JaVGuAUDVkjJS/7P
yJxWMgNBHsb6HPU1eAXmgylw5/d1j3pNhU7nfLpKoGTOPkP7ulJFoD3JDAyeIkhAM+xpp15KEL3M
E3sMm8KGSATWbZuZvEXNOUSDjIS4QC4r/WyQBuEsskhpRgkSuNe02XJDPWfDN+cMKoanmCkVkzvx
7OJtSUM9FAN8dFxm5+IcJytamvFZd6CNC9YKOQHWrPkVH6sIvytRm3f5SfuFvmRRFfvnQu/GttJr
bSHz+P8oj0i0tgdd+/kv5Q64xmnsovK3GPlHFM7Ysk6s+KAhwX3RqjWrcC1qUCB3eLfveK3y0YbD
6L9ysIwxChh9P7i0YtYDORGd1qc41bFHavTv/7hdF5ImYPJCg35KmAg9q0rjYK7FiZax/S/aBNtn
4JTMiTAXJGjhjM07DXyHlSzbxBOJMuxLocULrxdUXDOHPnSkauYEiSvDmrjXAUrRHyjczj7ZjsOM
ANiG/NKGtAJF3FMF0wTALCsIj2VEAB7ZFHJt26zSBcphk47b5whbH7RXiW0Kp2squE31oRhjHcUX
MCt0BOab5e5mF/dWwO6nnPOzOJcW2JhCwSVKj3yEKRbxGpqRfTKy2nE/zkdNT1+7uBrCEK/sE4nP
R055XWHGQA1ILWGQUD8oV3lqVy+uuCbNjI3DRL9xjK4vB5KdeTSJAx6uifyG3HUvDGrL/Gg9farI
7I5ThFASBG03EBK5xKVkwEfIOnpEvC7AFFXrqwWH33L6D099HIa32D+vxX8vt3i6TrQ/AxWjtP7P
R48klu/Zn3V1qmd8eyeyrb/GEwW9Xlw74Y/mvRqrv6lQ8B2XZlPKAIm0kHqI8VprRBVKxyp3eyKP
oIibtlqYWWBYHjQzjvH+bLcH2AisQpVVLxK47EUENhKfb/8R3PmGkRQ+4oeaWN9nmPE469UDWBte
gZixpUCTYe8FGkdpU/Vt4Ss6vndTik31BgFvPAzplK3gTo0zqPJR1XER1oPgAAd9YtojktNvSl1H
6Kybm7hcS9NAwwI3QauaJROiZWMYU11A1cKnUW+GjrDYlQFDqaSqtbIJ6hggn9h6alziD/fwNmnC
gWSt/USCu473jfqReDINSNH/1CUJj1L2tiOlMu5wk+mbNZfEzZlUTsmE5oLyCisgi9BhZAJAB+Mb
58aC/JkquEzddOuZMvT4BXHzWHp2FT3YquOggFs0g/z3GwxyRsL9ZK1gsuYbHxR9xmlgMhKyZHvj
IWDvJvPCNT2NHZsvmcOjQV+58Qyn7bCQP6J3LCGxtwFJwr5peo7C1Z/DWdM+jrNkVGFV7Mkvt8f/
jaXCdVxqwJXuy1Kh3n3Z+LM4MUx9osV+c7ujsgsQxiZhN9VFgFBOExvXReRLvDwrD0sHo1bbNK7t
dJrztu7yd5O5X6F2bYyd2ab8c5YorxUeob4CI8uRVqT8F1GmAROeJaDRj6LYd5TcrI/tfFXPdYiH
3Tlt37Ibgp+RdxXtSFITbnkpg+0TG68lBV95zXSwQQaOrGfNFyK2tPJueBQtG0fZjwmhZ6Q0ETt1
ay0oNHk+R3km8SBFgdz99zBjkXLuEE516G9yoCUBTgmyOobWbc1JvJPTjkR4KPm5hrGiZBeY6cmn
yQy7OxseQF3201QtsvuQla/K3lE5WGqf3gx36e+CGi7zPuMBgBPnhnUBxN4T9OtZjui+FbElhpzV
0fBky21IBvI02MhpQH7+FQx4qHqDBlgVn5ybpRCvBD30URaaB9lM7XdYtmEJlBhJh/Cu7zEYV5Kt
cgESXXc+TfJeLhZcb6tjFruVkB7D5i8GzgAwp40HvVJj+Bh+aMFxqC2A4lMb5Qp0KYR2mPMqyhkZ
P8xftRlonx6ukW5BJT5EEhFSC2OVaCA6mL+1Ri+42wKxxwUe0kmCwQ48JZsGYMfmEztra+a9pxBQ
n4i3qw8/PSriTvgbiwXSv9RVpNXunBY1TFqTpGH1zlzSZd69B9rRsyboHUtncqK65BD3Y5F4WzVS
oskzIpuqHXSxp+Ted7oUNn7lKAtptFEHvvogsmCiXKxtf/00KiFHtYsDz7gxXIxFd28GTolnHo0Z
mGNoD2313VdVtVyzDcxh2e5rMAkXV7I6aqzIKLCUwijuqGV0MKWsQDvlt8N/u+CoG+W1kiUxZH4h
8rwoEGUpCC3aDw4/VuEfxSJL7qyAsLpH7a4XAGtEyN+wkpPxAXv+lRw0x1Yn3lEqFBtkjDGodBRw
UaC+Pfo6LJIyxNmnXystxf7rnGIJiZF5rr0tY4z2ocWwI3xbDzPW4mLb4Iu2v/99gy4genGAiuhf
rjcyFVoafWWWGZtxlgoxbbSZ8T6xfrwHgP4z0X8Z6592xHebFGL8z/0lC3Nh838P0kvxq02GXnkm
I9dpZ9pdfGAlKQ/1Ew72JIt/BgMH+Mijf5rUh0oQh0C6dzMDMXxeKJMHtSVm9rG+5ICb3ZU+ErzS
GqBgzRuFfRiA5RVbrZokQskqvFAo2vG9UX6PX6uyAtHMPRY7ATIQbSlCgzzCGgRxv2RCveYzVjwy
N45hmtFrRWhxi9krZLNuoYwssgCci1w17BDECuyglwlNpjLNxRXTxTEhS9AOZoe2sWQTB2e9DhcK
slPVyhPoPPUTKtva88jRxkx9rjYAgnvnujxeUvEQjuKVXpg3PWxf7Dh6we1purzaLfQgIRrYSB+a
GGfQEmA34NGMgy9xXlOlZ5liMS3431ZPz4tshoOg/T1MPwxVQsSVHViaHKZigR+LjDGaCZszeFIu
Rut1PlbP53Vq8P8OY7gzkW1i0kuqfKd9WPsv+77vWqSFBnbwgRgveKxrqUmsfH5gRUzae3D9HeRJ
Db8VI40kubR6tjfIJ16EIPmO/Jg9kr/fCK07BIrM3UtiVq6J76+3pxlzvoFGvta07U2v6s2TeiVp
WUkr/kvczuVpkSlKNSiKUPaIUU2cZJ6OAu2GRhyB1LlwEvM8fDmgcMo/yh7rlsqo0tbOV6q36ft9
k0tPisDJpkDsbosR/76A+oQSf0g3Nt+6qGzoChM1OQwAwstuTC427GnJC3kBzY+l1eBC4jS2J+eu
h7QbiLXnxtEbrUPCP0SJQBhSYW/C+t0j82WTELkL7paDhASnGwkJqX4Wk6MEsfyfbo+pee6xXTyS
CqfjrISwlHW+5VidaVuq6QoXgAHbStuFcniKajxtY5v44BTD9HNmu5BPUoSMrMmg24yGTNi7agIe
FbQ+5bCrvhqjeOifz+OkXl2tcAWoqcIgWpEXMtNOLY6B/oXnW1PaB6z/OJY67K/XEpj4wACKtvFH
5aWlXTWIIypxX7MqcUNNRgbxdo6WRTUUfr5FTSHRAzHAx6C8GytMQa0ArTPU6duvrNC48Tz+cvGs
Y2cwF73b1JtUOXAaiEgibHk3BV6xA8GboVqfZBJgfdY/NXs8FJqfUkbjOxWoFlItw/8u0EAeZOCA
j1Bhz2y0go9+q9YYdq4YACWQjVaM6S0MvfcxTSCNybB6tbYSXtnVKbK3ZCp7coigi7bwSFAeM67v
Y0jg7wCyQZlvLxua2kHjncrj1Uc4MIhTLBOGBIcmqvwowroC/RvWiWRvltUxkO0EHjEoOOE/40AE
P3mtXV7Rw6AEPU/n8rgXTyYneL/1y91Y+J5GAXzKWemD+BYhp2cidDQI1bMNjxbBZdvZh3d/UYIk
f1EHrVJALNF/k5P5lzpcKwnj6MkTa7D6CvRgpsPfpp1+G0PhX3DYA4LLb29YBodUNKhpko5EMa8z
DSZMvsilO0MK0HUZfeMgStYkJY46SImBBt9ULlWZGnmRBAocJQzgdnvoVHe3sbN28F3BVndjfGaF
hokTGrZ+BG46FdOYQ5Fqq8BZcnnfOn5ups+rJ+ol7RgJ3AEuxEbrQBYVAqJA6bWgtdjKVCV9Alfp
ojwDuNfxy9vsI8GvDbYWAn9rK+vRYB0+MGUU+4GPUSU1fcQ/qh2Q2OifsX2gENt1H6i8z9rfASMt
tCHNpYjyY0ARKK5z1MH46QQy5c3Aoagaw4rFmapS7CLZnLJIouu0uLbXem6/lOUyvXnXcXAvKKEm
cI1ziOsglTLckKL5VcGF5SHMJXwXxRZ/u4/hC91np9VXdJv/33r04YKql13Lfj005XV+G9we8EkX
WNUWzWRYzeMf3m1DmsLNPwp5pDgLuUbFr4VtUdZWduCKigr1eOvsn+9aPKeGboOy/63CE+9F0Khb
IakbGYTihgzBcGhEeIJ6nHxCx2QSa7ma1xXqIwz4uu6ZMJnExN1fhcORUH8F/8268jC4n4ZMSU9q
z6AzE8c1eVJ8yvkN1jOdwrQv/U+6KdhWbkBMuFFSGZoaZ3Pd3+mLOdYZqoPodf8XEjM/quYiJRoT
zsFFoUfsFHelzVB73sATYnfGpeexxVyCdZmBcP8z/4lUIUKqwUJeYIBpTaCk1fxJIJkeLiL1UVsf
f1K0dUBnai24eeviu1XrigA98mkSLRkjCnasRvDkAtc8hYtT5sP8QWKWypnvz5FETOPw0wITqqcC
tUsGSZZBGvXCMri6Zco6VRSyovyQL/pUzuFHElSXaBQvUnBAoH0mT9JeRmYxMTe7odWXEiQr4Rv1
vKirJaa98tY4EEwaQxKYX/VYa1J4aiho6+gRBpycNLdu+fXkI7dpIKZU301owEaSELhGAMaLL60/
aDIGBrjjamdSAPvUCUD9nZKoYrfVXW0v4HwBZ+f1puSUu8XW2tZT9NwDzh2swWY1u5C1nK1xr8Zj
oRyCJlq6bVB/mNCggFGOOPgN0Ewd3IlA2VMvfN5K2TYNKsIZ9qHP838X39xLQ1GkH3sPpNiN81VC
TQy9bpa47//ydvykKxGvkNhHDibcA6RJgNcapeK+46nIAI9nadkdOQKMFo4BL2CzHTpaV3MC9Mq6
U9jqu51V/5s9sVRl88nRUD3AyaSxw627zDX3DnAoHkpYHMbyMA93DEgnn7mpkYbbydz3lnzkNBC7
3sDVg2qUS0fTiIvsxbup0ZZ8MSoRPvLnWZDoViUXOq83ECJNj77wS//CRNlF8E8STySZN/52dnKL
0U/+qfIYJrlhYDsSvUKtMh6snp6s4o9Jek+YyO/eKGJQEwyNr303Y6NuCtj/gLYuJoA70lNk6Eiz
lUFK3ltC3fmWl1HZpnz8PkS3YWd0BFjWTpvg3K8uoPD8WrniXW3YtMbhmJzKDolN/in2qN5tkxbq
F5xMhqfGVM6nEmNkhOzOEEu6pdL+VfpZyDYwK8weFGdnZUnRPM/a4qU4YtUrG8PCrv+dHXaygD0j
PgKOb7SddOWF+yApmNcthdAEpi6ezonueGjn3X4r2HxIWXpt75yJ9gvTEOOredH9sqsDx8fOti3f
LKRNUaYyPxS39gADsNmR7Tl2M9x+kdVywUWyXG+ppJxG54yjr0i1BQRwAYTrSNjJ5Qy9j3k+0nTF
dnls0+UR29TuLx4gt/gJpBZlNtA/nfPwMVFpJ7pawKF4hZTZzhe+71EZwB0Fd5Ccu49+y5kNWJOU
Npt++tLX41qLtAxkZPphPLxjwLvw2Za2AJ0HyGgpyT6bc2uDxZIuc/YGrMENdih1LZT79kwaOC3t
4M7TQ/7srxao2y4V5a5KzHQaVtLIERUX5TYs+8MyXIQxZryCdhDbq6llSPPrQB8KVBZECHMUdXmV
RHDgy3UwTl9OQKgadSz4f3mQJJnAb8xScJg2VGPeo+ni2knGEB+9srY3tNlJrq9ReNRyIdLf5uRD
M4yibVUyzjZC0dyQeL4kvgf1CmCnxrGeGtV3qChCdQQbs32Aa1q0+ETVjwkfL87HQhHP5jEwvzhf
pJ0CxIQDBV4wirOJhRrk3ieiJ9vJDtkSyxIxcnN5/QPzDjOoSA8gpJwjeWVKE71ARI2RocgKNijy
VzuIxylgZvgAYmwIIL6O0/4WsJL5Xb9vaw5Davb+oi5fJJgHepuXEvOzD6OSsSkSDAahwPmYLguO
Pe2zUWr/LkfU3+Jgq+tni58A20mpK5niMuN56OVkeKOPZpVz7xhHyAzqxt+gcDUtNcgAhuFqs5Y9
eWt0MDHbq1ePN9jzZ3ezxzuIpB4Eb5OlEkwdlY6bftUMDtGWrEPst1v4woEWkToYK1iUThJSRFgD
ec/d2tMFqwqVCK8ACw+b+VxdVZHV7AG7XToZQpWl8yD8ie8e2kq2RoPP4UhalBjhFGm7Gv/OU6P6
Njo7LN10Nel1Pcym6olGNfip3ExWvp36qTZZ84Q+2d9Bz8w1sZgDe+yE0UX1ZlHFFwVUJinJvNCD
qe0spFdBWZI+zUnEJZz541SYykyhVCCKPUjhiY48fqG/S3jt7obVGmWeyB2hy9M1cqImwupWvFxL
slLmHwKs+a2GKdxc39KWu1wg+sx1NslCe0v2Kece4ZhQZdncKccuKDexLuE8Pe/mgQww0UBa7SwY
hvBT1AsTXOVrm5KyKnQT3ufhe0IBb3iBCrP7GJXXh4DLLzTbRYkKBbVUxHXejJb77WLOB8Cl17xG
moBa9DxJLnIbFU9bgTgqR622MDRUyltcG5LTJZX+O1NGJrhrUutpQj6gKdbnTnA2nKSIJDIeLPe3
WQKc00AGTcU0vPW9PMqqcHxiCROCvuYzPl5yKLWkNYCp1Q+ncdMokDJR4Aooi8VJfxtxm94ARUgE
1b4SiUzto/dV9nHqRWuDkuCr4EAyI2OJSabjzxMgcRxjfseiJi9P8MCDEteJzTFGa49UpXAqT42/
Gqv6z9/OIy+VORydSQDvHF2S3XDb4f8C2F9mRjkUqhoAMvgnWtKKUQL41fOnqGt2+Iscvbg2kApo
GpTLDvv9VM7tDWp5dQ/ESspxPp73OMcGEPCox37tSu0+OmmwMxEaoseLZI3ACrrNmOkXt57SfJAZ
n0FXcEUvJf1YFVKjveC+Q3JxzsUA1JB8dLK7f0GbEdJl98KAKM5p4czAfqDrzOaBZmWe6zs8jppX
ATPez8EDd1K9ZxG3VCjhhB6FOGeQ5FxvvYI7zmVaTY4SlPkqpQqEU5BGCvjeyrI5UacH0uX2wNeB
0rPMSRKnLQRFSiv/DIvLKdm8xQABfJ6W1UP7L96MjjNJHStzdaNZvL0x4YnRr0GptoTWJRUARiNV
25gbfL+GibwktMTvZlTuGVdjyrINEkxmBqObvYErA2dxQTDaq2N7N558nWE6tVcWrRY/2AZjkp3c
TrffwvKZO3bzEcnbhhHyK/Dzd5K48HshTJpCuhlymvCwrgK1Klm5WcB08tN4oaTv/YW3hW7tJzRB
AIw+O9bem6/ATIH9wq+RJvgiRJfr1cFiJ5jYla23q5amapymr/oG9efsIVFE69zEQU9ac3JCngF2
pfNubk9d2iHbKwnoyUOH0vrpKDZ5b9sI7iHoVnNLEo2vVBPUTVjeTvAed0b/nJC9+K4EI1MMU81E
yFgeEjmb3yWtORmxTZOd6FOMex+vdvi1IOT/VrWy7GP1J/AMaDwFCLrz4TLTmebrIxAEDpfvpV61
3OK6LjvB4g4g1RACPbUXE0QSnGz+94q2/ILbWVOb6vnMmnXrPwSBFVKPvu92wODNBagDbAzC1XVf
/OHiB9ZkG8remdGaqrdBjcXqSiT1/2gzgqcjyyuicAZlgsUMngRi4MiURo8DhOkrtoo8/CdpKc2v
u5c5c6Mi9L1mNYEzyNRAm5bAqrNn9iHT6IqREdLHfEfz9B+3+xXaUCOq5ig2KVf9LOf3KWXVyKQb
4eoRpg8o6jBtD/azDGsfYOO6MF1GYNuKIcwteaMfe2QHAxaUdjNtLjnACuStHDVyXFB7K3byfwvk
w+YwyL/HJdIV4LjVz3Nw3QC0MBkfrLGcxXe+AFC3RnLtg6Tgby6QONtxT2Jy8QG4WR+FHUkjhGMi
P5rduS1hjklN4VYE+mHXWr5JjlNSHMSBFuh9sZkizTiMVwS2yyj9Dou8ANGEaRMtjFr1L44+KoaC
cRnLOkfcm7vilTfWxxOwora+VXm7tqPsd2y5KVYqDIABPQQ0Ec9heywTAI9Zktx+n9ln3gW0ugmA
vFWA940gsR4GBTFJlceFzxdaNdJ05tbCTFG6F4CcUXaMyjN+GaTf8eKt5ELTdBx6PTh1hvPGG4En
1jWDF3HN5XOjNMDFi9WskoCkXUqOX3aR/FH8qO6ac688JvTkT4sObtMOhz/0IUP+s8+Rc5NSdE+H
98EAUnqDejsVv4tM2lyvw48jMyclL0IxfHaQPSXeIE0fgbx7WNPp6Hi7lf8bH10qyr32Seb4OqmO
FeitVmQOUbNnZrIkkCk3TJO08pBiainqGoKvhKeByaE5iMcyCjh2aKFy8PLxNBP6MItPCfFkSsg/
6NR4IborNXHxnjhKNse7RuFAeXQFCX4/ldL+2Eb4i9C8hIrR9oCAcYzXnfMdEC73GoP/iiwWakCk
Ogz3yEJCJLykxDj41USo9tLt/7luhWtIAEHkJU3OM/AguHqx4WcuOWAxCNKGKKmTN+g7TzWTvnQi
XpKfOdiotaBuKhQot/egJ5ytb7AEA8jZRBTe/3EmfvNv2csC1qTkbsYGay1RoJStJe2CDJbS4T5h
zKlpR3p+CyLF4tagrShaHExjYl07fnayA381pzFZxEm2gGpwPGLY2ekFkryH7O/YDNI9F5/97Zxa
gNLRnnwlqyZ2V8OrafBnOlYUDvWv29OH3pmyBIjwgj6/e7zU4Tuyu+3CDrLt2aig5UhECPfsTwSC
h1035jo/slBH9GatmLWlRAExovRV5N74K/3DIQDu9wsC4CUq9UaSYE896krFyqgd+ZZqehz1dmZZ
WsAs+UcuMTrT67ZT9K4Qph5iQbBnkKdDU4ZkZ66CZLTHtVhvvEcS8gxymfCdasQeWuCT0qijeuNu
I/6gzDECQ5LmWWZPrp+e2+vygZoM54cW/N5GF4F8RZBeW5aV8vX9memy6Fz12p9qcRUEXBsaeueZ
H1ccJShvObSfw2ek3FQufmdFC52IQisPNA7npOCgqgPT/dogPy0stUkgn2Xh6Fxq+QZm/hRs/tdp
3Cb1G3zOgfEdu1143Anfj4X6Hp6Nenmkz+T/Z1PkNtJ3cx8s5LTHktdWGJEwVwYRyyY2U+CsjZ3q
PlNVmmv9zBY0QjcF9/Qy/m52IdZFFlzY3kLk4JSEHxr0+rN7Pl9iQloPMekpXbOT/VOCG0deR7BF
HAtRL9NZAHGc1hGF+7eWIYZZyzaL7FNTF9EYCVlyHlmc1mn2jL7gQczUTiJMAosZali9wW8IPxQ9
bncKiFXjs75+Dux22RGD9vitjqhD4O4peuwsNKsgHONyTXleQ2pdCBFJ0dlHezBDbpXO0taSVXkW
oFvaeiQmi5xGH28Drauafvm4i2QtvDP4wiGQxhjd2EcZg7514sA6LQYfQImtnvA62xvJnYN3R/uv
1GzrfuA8mVYPuu1EAOTVyjPdL/i+XQo20EWSmC7Y0DEHj0NZbIHRfrd8kGRAgHyIptZZ+pv+t+Cx
OghJrKqEox9jlUINsMaZ6tsPitdFrXL0zMR1kaP8CZbMZpE0ZXxi7TErdY72fmRs+/VLOntW1dDV
EBQ8rW7DZp75BsBFlUYoz6HtZPOWobEJzAQ/JKLgH2cCuKh56FIcZT49evYD7ob54D1Hrg/6Q7Kx
WBUEqS2F6D0uUhkVMa+21Te2YSLJ3NmHgoH4t1eM0iLVpaHLdHKYf7T7gH3ZjpF/OORQuWWTmZUh
f975qHsS1hBuegEWUoQD/GdvyWhVSOMTWktBknu1leV44uVSJRE9F4LE2i0qwEewC+P+6xQcyKp+
mYdaOTMg4FbgCo9DwiAMZuZTzTi9+X+kf5V5WHN+psUcw6BgEQIEpHEF9hkLwIVdbadofpi92qSc
v/Aeb5K3tFXvE+Rwn0V1syrPWxdY6GBPWlGSD18EPoB9v+FCKd56hiQFn7KB0luA1j3bsHTr80Du
SfgzH9q+mN3t5OUBuhI2ETKo6fpJWeu+eSGi+OH0dS5YDF1s5MnXKQtBHkv2QVmWtUzfojbQhCva
LEC0TQd4t2Iviukex5zepMRsjMBP8ZWhtUxh2WFBtTojPX9dY2leMy5x5Xr4hRgwX/AL1lkYy38+
Lvmb/xzNbq7cdx2M5tzZCpB0BWVqMkPnBbwCili7NVKHBWIWOgCRiRgVS52bkPtCoMmUdT3QdYe6
V2vPLXAG3fJExzssbsU+GB2Ocyw69iQZHJtMqod3AfiNXXHIA9D/WQvdujJwN64cJmdCKS/mvgNq
RQUVhdnVjsUt1HjY4tSQi3lkD/KWQaboacFIu806bKmL6+shTA8dbKzAArBJ6wdYQajYuVL+cSF1
WJcjf9q9cL6DwsjA8XAXVmspFl9WhZelfyvjyTTFP8rPvce6bervldHl0r5VvxRk4F9XsKQOGEpR
zluLEEQJwGjzhwZiTWshKHAbshuFMHbh+2QLJRe/WCM2HBAgdgROLKIgd3gL6WMSliaZQ47h+mph
fNYqOAYerghp06K76RP6uR7Wpd38yR4+9OsmWFm9LDhpkhJbFxD7NONpIY4BW+/GyxutZ0iD3met
sCs4oBZXDW/QTw5XjHZ9NvcsxEdktSOus2zecmhgOaL+LroEhqHkdIZGYJEAjsc3sHONCf5j71uC
2/wv/Im0TatXRZ1ZVn/YleDb9TC/JrfXiV6iJ04hQWM5jxCOdrPZP3oiZBP+WDETN9GzmWD2u8BQ
ZiEV5MmAG1ZV2MtvTeKkZK5z5GDj/Yth90oZzMPxFpQV67B43iPFAR4A1OCrpWdgVLG/QK6Q9ksN
+NcNMFAnsMadhOrCFs0FbU4cl/3p8DvTybS8i8n08+P2+mvfqrVo2duBkO67cMaRbQqQ+nVQGwVz
8kGxGmoMQPNzd/hCtg/KSoQp/xpCJFQPvp5nYZvRbpa6SQETFi4UmW2QhFX7Q/wUwvitphk3Z8EP
WKflM0brg9v1SjWhohM1NfJyA2mNzd6dw456iRUYfPRhqCgjBovoOvhxq0pQ+MuM195FSELb0mTl
ApXVTPzZS4FqvHQoIo7BJO2r3hF5Z6qvGmGdKpXikDXcuxUGY31XAuDrmIhwIcgs8avVmBv7B7p3
NBjFfTtPWgfO/0/RSBmNgOsANVnwD+8goqR8BWMgbiY8hn5tzcCy0R3ZngzNrLY4aCBFOx6Xo7yP
AQl1S88AeOsqtrqbbZPqVPJs4KksQXW8Y3zsDLwP0wn6CiS3S4bcsv+p8ExBRrCErI2bSj6ArP0p
Q7LrGOwA19E5Z5naXYher8K0/aYrvS8DfRN7ket8JFYQL736IN6CRu2NejW5an9yBiPYRmjxygim
jnU4+sm69tQzbgWzCTOyRriSeeLQYC8G0u02XyMPW1dQyQraby51rxr2p5ULjCg4mUNk+oCx4kot
3AfOQBbmo4IgwfMBjRidvYLQbBscqJdw5+R3zIs59U/dO/RBM9m7fj/q/guyZr+ymKsABukGIZGt
bEv/m3yTUiF/aS/PctkUTmEsj848Ivt5/jQ5Q00WA1ZeHJMwW3j2fmFtHfITrcMnrNy0orLAj8SG
YtdMmA2qLNKTn39S11JD3zLLFXDaEYGoZd/y5jJYhGwmA7EbPZiSCmzCztmDowtN3x8hRZuaizLn
D1eLN0srAcxXj730RQkFNt6F0XyPnH/6HiUt4UvfTmyulwhR6QdeR40vIJu99eL5xLn0vju8bJl7
29Ja6kNSKRQuSgDpUrb4gmexjzlpOR8g//2jUlRDGkznGNpBkgCJ6vehIsX4bo6VuAq1L+gPbc5/
kSzvZaXxyu9TTuCRhvvJJDK8e8a7ZK5zH4pCxnKzmlEqMJIPqyMw5bdTQqXE9QhbClzUi0WxM7Ai
TVNs3yTRmYtyOS11xbicuQAV7Rojja1L8qNIdJIhqqX67a3pTYcyepm025eHtA31yqzgIDappR6a
IxuiEn4wjoOkPKHPQAhULvYI7oKz5S0DHft881+EdjuymZ3oaT2F+rQfbgcc79YSuPOKEBT2896k
i/JhhrzKPE3ShtP9dXo8YP+EhyclpvCzx2Z8AmoqcaL5wHugLRDwJlCb+DIL+3nMu0sjqINyInVW
p8n8QqAhHbGaVdk4nXzm32S8mHEYnIaeEVRB5TLnTQSwVLQkMLbUhHnBJ5Orlg68v4wLNttFCiV9
U0oGEFA+j9TWyD7dzgF/zh4KEdMXqXmsugdhIx9+UaoMRqfDaOEWthAS+7EXtyz/OoMnbI5m5gW9
H+b0qjEvVWleJE6MLObhNdx04U82S7cXaHCLidhs/q/yQMpyYnYpog0rZNIylJoafBLkjQ7v4WgS
k/hJUWQxVFeaI1XpT0HTu1YIdso0UKgEQZBj9Xp1cl+8Rnbi0ZkRQ0ulV8aRz2+pHdRF+wFXeImO
IFz80lQkfsHu/b9DdpGbCNtxjGqS5LdodxlFgVVrUdD0Fe12ixzNW0yau0W5pa6u/xPsoQuK+DrR
xSL3llMzs/rkhvaVboatE3fkGEqvuk43NL+p0vJz2IZg1MJKL3dO5WXqC/CEENfJJmTcGQC3L701
o9kg5rtcVEfe+DHfDel+xRhTcCcsPlgvCuxHnwnXlBX+V8C+/Wa0WskGkQOBE3eE3IBL+AvINwsV
o8eWWgyXvtROfB9HEgpii+ihMgHE0LkzahjR/BVSE+w5OoQExF9CZ3Not4O7AEHk1Qz6VkdIaM3X
g3FhAATaqBrBJcSGJ24BGItBtkk11QkJuMrmrfsohXnyXcMpf0ZNw3FeqYCG8V5cZHmlIOjoOQk+
llC5ySV3IUUCK+BzPUc2A5TMNaYI5+gm0RUgmpuReZK6iEesO6xwglS2MfolcF90ZNzyfnvqMCcS
xEJr5qMP7cv5KMt9SWXMI2BAxjxcIh9Cq40JVGuWGfjPtnQCwhr+SExU1jMYlAE6N+rNXB1KZBdj
lTZgjsvbN2I420KYOZbWwbFrEIwg2lVMkRvcS01zpuTNPWgDFYAQ8SREtNVm3mnMskI6tq0u1ubG
DIP2VprdsyLHS4lqybPVOXunL97GeOiFC09nyV3EhFKEUrAjleZtHiP+AYHp749MQlUMcOWmB/w3
7mbhXDXS7jWtRdTT/skicjBea45cFTZwH/6f5M8okO5c6hfeGYcirtJd92N/3+lXQFRqbsL/4k3V
QlBrRWL8LGlI9bnSKhO4xvh19LWg2UPh95mdVSA4rlSGpNUXXDzZkdCvN5gBI4t3y3ZlNb5Z5BAO
jjSShb53SQDwvVdcqrJJhL9Dj7Vb6+8GP1Mcfq+O5VZ+AwFZs4WUhHHDlXHex4r+2Ij9/rDC5Ahg
qXVTm0mdIAs6SLLcxuL8WPUEB0ANgAa9TaEdVu5Zkc9ITJLmxIBsTxos/h71r+hgtkEfC0QQoOVz
mqtDRMAzT9LnI6/2gi380hYxUajmkTSlvyr4BRVrfpgissR94JeMZFxRRYVBwuPnED5fGXWdDOxh
Lp+KAXsX45H45Q+xFJRC7RNdTROItNsoNXa4yTacI6TufkZ8OZd+wE2dRPIUqC50n7bqNMo8M0Go
1hW3iOVwH/yd1Sz8lK45k4qLog7zsnRYVWIPA3HzSIQoUlsOhtNYz9wQmBvBMZdbwLufLwXEIaOV
d+84bBZ0HFEhRlgr9+3nj+Bqu2R7VLkK2yxgy6td/cPVUg13y21l63PDSFFMeHjbaqjppAZNVd54
Cup0+jJsQ+Np+zVEwegNh6/17ce+ActHMeag08irTH2v43y0027WU5hOMgF3dlp+UOsFOGXTAfVV
uXv8kGHfLzFI7nK07WWSASU/pOj0RvJTBke3EN6AK+KdHcOTe2djHOIqI/uK3dBvQow966UJ3yfh
PM5D7DIM0BLaYkjnXY5+xyymaDvX47iU3ZHKSTIdd4Z7LgkkF6FGWLzBe2mbOfKLv8mZb+XKe2AT
KYgspv6n1bCC7vguMkgPD4USyhrS2ul/Iy2UmZ3MHXl9xZxGSNAiLaj+cslkN4iss9I+PdVMam4h
yCpXybVdQkpeq2ivByiIfVnqeHiswgltk9eG87dCN1/TKvCcTq+J1FfK+BLE6RJpYl80QskGtSed
iHNg7pz9w/h7YGQVyCwspzqvyuPxY4GoKYCOOxMkZjvQc9k5PqQePWVVSRqT3K1jsEU47zu2c1hM
KIbyEwuNq+TOofDLF2LDfYxSslLYwuQK2EMYWCWJJAJF0nYzb9ms1WFxOcbRotAOnGxYBpeSX4FB
5nmErajDcH4a8GY9+HclwegOxSRFsqhZaewMfKtSNBlzVF9muEQxJngQc6scIF4VbL7pD4uj2iBQ
oClnZl2KIxDWPRvV4HjqhebN4IaiJLrkq/xhxBAPjNUm9+4x9WR3YAoR2cwWtjB6THJoYjxChCGp
1V6RY8yQtBuiP4TAhFCZ6i00J9E/HxhbrJVfkEjB7ugNIlSFY1EymIZLIPNn32UrvdtljzfXDCqM
LRpcxvLOtSHAiI3uYFFrde/3ONYg/GCGFSm/3M9cSwxI7QXSCZwvd6ulG4wpRbe7+VNZN7w/qOKD
4KdXAlPsmHMACV0OZITX8l5o1yZWFWDnlTMHfmB870kvu/+IIg2iaTNhCkOInVjsvKEtYM0rWeFE
sS7MtU4XYik7P9yYlbmXThhp+QQhomIrX0MpIhcH3YrOOG2UjobpoBQFnCSKSUTRt6WPXKZnqt/n
BRGrHlmn2vugJhaVXy21CasRwkx8sNuV6Ft0GgWpuO0BegZn6bK8X8YISfPxHLSgU3xHqLjdulfb
mNsnqncEteCIJnvKBTBV5/NSo53FRqjQ5MJRrWak/x9qsU5RMFJiA5qPZ3YpFl+Of62j7ZF9cm4n
Xur9FGnhSs8aq/B6GuCNhbVo6rKwnsFhGJzcw0Opg0uGOPXvVh38Y2YTOI9LsJe8gxowYIA5jJt+
QxHAQH8K0d16pkt1DGv53dwzRGa+m6CtVghxJckSuAakBQLni5kqZMJjs7NgAkbRAIOgF2Q7r0fL
hqzE6M62Yehw5ra8hjKIUT5IYX4FexkqJFWbIrnoSFey0z3gDXX5XN+lmyvOfQF93R6OGug3Kv6o
waDbbcDhzDhRFRJl2+TiGhwR4yDTLoPxpau4SjZgIg77fsZZgmweLQanParpPUYrL34rMM81t3Rf
6YCxnJAg8NckCDWuDarmnXJANCNuGnasUlyE/tXLxK7YcpsGJI56arGesZ2RYxLTZSdoHu6fhV0F
t11UU8bLkqAZBviAMFQCaZ68xVRWmrLKHzxdpmn6Ok/YV8JEDrwWiknsIRkjQ5nQFwcVkki2yUMC
VxCSHUT+nqAV12NoaaSPStVS3jBLObAcXmbNwTKjJqVDl/FcNkOlPXXtax5m9bLO0ciPXIpZS92D
kNaQPoxiwuVjiL4d0pMRQxubLLjeGtIONwRUXFidMMuaIOq6kcbpX105FNmcBwGIt2sbCZlx5HIs
+rKG0nJ5yHtHzjgfl1/rBAppWkFBZQ7LMCjEPJWhDyL3+6oFjpJQb/EkJ9FPE/+Y/Scma1+ZZulx
UuubGWUhakTZL3fFA76ZPk0K0vXpKJEkAmUipC0hAD4hhazldPHLPWp65FMskebS3DIsGqctkeDG
kzZoSrtVBmBHwBFSnBIl8w272DP2BTNQzYakND4cG3vRn6mofe9ohE7mU7kd6GnEFzZpaWSjMlJP
CW0alQhefZj8M+3jMpWLmp2gWY49brqAW5+75oNLREZZai/2l6A1NG2zS4pUeeOB5IfWo0Iq+P+r
2HWhCaLde//flCisJq4h4caTKGATQ5DOP1rmMTBh1BSnZI36HNMsxX4+fr/IeFzxJZblwhwxzPGf
Tp3xGqVzXeX4fAaN5shNe3lvFGsqb+pOCt42h8ZHx8H+b2EWOlSl5te1ARay/7BiQy8sf0/QEMgx
yixkhjI9NiqSM84GpDZ3UjmtU7zpyrSynFEX6e+Rl6ifofaaZXv6dZAlM/9flWtYL5AEu6wpSxvQ
2BLZKAqmY02l5quGZKvRYJDEdpv8UmgbjLV4GK47k03KerCSRjZineeYO/ctTh5TtxaVBJk5S66l
g2PhFHlok/HEHyBqeydOfwn0ZKID5Xy2Zcot5O/MjHoYH7HNCTPWwRlO+ifTW0u4uJouio/7gjbL
y1coFAPOHWoefzUAdKxiurPEovwPM6xk8wXMFS4gaaN9RemJMTw/XWRNa76My24uIfFXZJ4Kr2US
TXjCGv4VniYZTytScxrwuTGmCUi9i13kuFv2Uw1SdkesVBkFoIJm5PGz3G1xdfbvHKxSH0qo4AcB
tHegJy/mhT8UZQyS3HDAppVuxBr1oEmEqK6LrNcPID2T/nZ/iGxYCx+2+Wr5FCchNWFQiPanO/JN
WZazWAZdqeQJi/rs5nZeiLwnbgI1MeQQPwxrodWB5Fpx57K+qbyvx3CpfEcwlqqxV8m7FUz4Xqy8
pMVaqqaGc1fbNfVx/Lu8Wf9uxbpCpdyyf24S5n8OG5OOG0o7imkcY1RqhFm4N4jsLmlSkR53uieU
J8igo1fT1I3zeunC8JRZs3jBEB3gU0bZDD5adBeUlwoS5Fz/5CmbUjtURz+J8ylYuXHdYGaPJvFI
uLrTAI5LPYghZManVyUPQ+fgwqruShN+hWH3Z4qgxj2OveSwPQ6sYCgs/xN/i1SRpaB8wcR9XWir
bshdybo47xmgkazWFPgBNGOtsE7yO9T5AlE3704RH4fZL8LMPErd4N15u51zWE/4gsTCy73x+GQp
7Qlg20CMIPFAfC+3M2OB7kv7GcJvTkMyeAtH/fAikcS3A1odrqn35KsPj96sETLMgLDObJYuXhGm
ivpoFMp9qXgSkZeuJDxC+hMyHTcUdGacYo6fLHzIeDjnQJoxgSq2rvd1w+JCEBDrsW6GvNUtD5Ql
RxQVEhpP04lGTgoS1/jk9GLr2xK/gqoZmZ6/++UDRuxtdpdSFyGk1q4iUE/3H5mnidaoylFhfMhr
AjYYCroE+KZ3pMJv+Ae6y2XPzwyDwpzbP+5Ru68nXsFYGSff/JtKlhrF9kN3CPL+K7ZcB5pFYxz4
RXUm9iD9bnj5c0uXqNP7R4rX1Q+oIAxX7dAcKy51iR2GOE+c/64gp9oBNnr16aPQbtGFB9PoszZA
xAnF7cGuMw2egWDjj6LnhE91A/PNxVNIhTlOoSyUMie+BHubxJja17sxzyz4qOwgEhl9q1ljkCk0
p0+UfARyixqckQOFvmMR57rRrjzQZdBE71iNKmvs+l/rFUKkCo3YD4fMvuI2zgPeZibegePaHG58
maNbSiumHoAoIXUbH4hhGP6z9Gbw4R0rwz9Vo6FvXMWiTBfdAEWOp+pauATm/6/Xj97q1jY6glit
fVRL/8CQjdGtvHj2/1ct91+eo2uXqUCsczmtLabvKgwMwmg+w1FxKAo69C5jRmq9jHkTXx18EiFX
E0BU4AJ+gG7vUCJsAcwBmDjP7ve0U/4smHINNkb4rBPT6YrJLl4WXlj/7lIOP0AeBEzyMUjuLWwt
TdqEi+W0nrzOeInCmAJHu7ZCGg3gMxH0zWx6Yx85xH+rGgomaVT338/M3Y7H9QqHEa5uJCcbIMxx
taH7aqMOf73tXTdFmC4oKFKnAujnRM5ZM+p8aX+Ls5oMq2vsjuesbVVRjYZWXtDboaYQLyqSihT6
fZ63lcRDASfjWXat0nEN5jCtiPyqXVz351e69h0V/iQOAyh+Y/E1re7fDaWe9TcK4L68OTgBriHS
xGg0jpTQsceaH4GYGCYLloZeMDv9aw3Cb4lA2O92X5L5jMK2PD8XokqRG4YlBoX7VDJb4NnFXxtv
9SMKgzT0Ty0ubkhP+TrtkNJJ4h0lR32YhetGc8Y6paUD7gBGKpRvY9OZIenbUcmb6+Zv6MBF2h5f
BwkKCJUDjMVh/BrKgh49fgvmNRLPya1NK2vFDq901zburx4yxj1J0icOmaXRLdIlsYKXc8f/Olod
IvA+rc06dRYI3k52BjbKz7hh7IqX8XlhJYLTyLpbispKAODm9QDXVPGr1yDkwzFyJh2BIu8kam42
VUFTET69rgaor+s7GltDev28Nr/T9Uf3IHmXWMPkPmBcRbRu6k0M50AkvXwuKiOktl8yN5wpCbhO
JM3Vm6gbQUdmdwK6AvpJaACmsG4S86MqDUg0Uxd6lZxT4Irq8J7EGNXK41ospj6mjOf4d9q2QPb5
eIwYTPAET5a2Fwh6xfWsEj2s3flKVCKKQv6DnXVHbqx2eXVe9c88Bj+7528VB1olZWr7ZWQJrc4l
j7dr7yYUBpeClrV75EaSBeZ4xj7CaGZTigz5WPthvqL5iy6+w39G6uhc/86HUnFI4pZJ2OSy2r0v
ew5BjUhSZVrdmXMe6cnZYHWbwY4MyRJAYZHekUtXRlncnWRV0YZO9zIiwHBBVqTKmD8zUt5/8q5S
By5/Uavv3Ts0hC4flBSmXmuE8GXMJQAjIAXFGZdszpL2sDcfsrEt8Kq42fQsvmVCGZLZCheyF8AG
Cw0QSO0m1TSFGJw9zuN/9ix102sfaldoN1fcsMX7Gxo3s/ZkZdbc9mL8e1xWMKgLgyAUjV6vSaVC
fppkSjafbK3Seo2yr6vclAdpJe7isUVJAO4K3C34lueDuBEVyTUMQ4F+Zgd8gIRtWX3nT50NT+ko
jI7FU+ddt3HgLLa7Os6AhGuHovwhJUbd7fxscL5BTX5X5ACjBlh7mufeZxfBIfhKQe4FjcaciJJI
QlCkZKZZxKKrri+HqkGkTkXCMAePW63ryQGPDG6LFur4eCh0uL1ZX/bnKOiSPFFwKFx89Y81xBTw
iPKj7naSBCSgzC4VZd8l9a2WkvknRH0WssAdQpF+qjEDhI/3/cDmfFDptqHD8HyRcu9zJdcGPFu1
lhkwk8i45bDBL76nq6Jgf8XFGeS1gTXXcVH4rMKyz63Y2GHhDilFShLuEkRhpxK3w8/o8AZ7cJKE
homE+uHsLpMZ50bVd/3Wun8i39GIAPMJ1q/F7vPJG0UB6GRVLn6YYmmoADD8gQCxHYzigjAC6hew
TFGZhbH+88QZllEj/hHAwQxm41SdCmVNfzAOHa/JOtRfq5wdKvtmh8fEayNWBqQa9JzjxLMWMubd
SoKxbR41wffFB/TrFBKj1KPC4YZpTGV3UPLQ+q3zcwUWaqeBcHGVyP6CTg2qRQcIfARUG0FH50qk
JOTUDg6IMqN7OAbGsjJrJDO0058wNeGuIY0HK6eItWuSJurB1Qq5cztCeG5g2czckkCdkc4XUDaR
pKh1jr8oYs3BdGw1jsYR4jK1/GIpPoEv985u8LIy7ClYsPBFF79eUGTFTjd0wh6CqOWGU5o7EMKd
v5w63i3C+VisDz9zy5PRyosVKAYb7HAGmnWg0mn/OErviKRggaMF00SjoGBR3dZHKzWsTHryvDk8
OcA8ZzV+6Eey1lt93OTLNVKLfXzsQ9NvF7daz7vwBDb/pr6ufELsx+pa7nBuQmx2kwyRZbiKNfWq
HfNm0aILLiH65enxoOGePaxntNvfGK2O8xGwGWQyRR19S/3QAwNhhfu80f3s3r3l9N673vrAD8Za
TItVDNkDCQus70ZYj5PrycdixcwixzlDRW1RRzBYlRhUlthgwdrsJmSONHeXwQx5Cvkrf0w0Ndk9
GxNRrEXJRNGvpOvybMfUSdJ7QCLqSphVfeaJaxq+EQphvfI5TjAhknpgFYCGJzAEznkmO2i1pVsr
TlmkGZdrBCZrm3OJburej3X5aulXo/ySSg6h+818KPASrq+EDDdWD7vApBQiBx4kYfZSk+5BOhQB
rvRTgIYJVpbzpYfykYYonoe7z666dD+31yct2HZm1/X0ZmLbqF0+rLotvVcH4fJM7BALJpJfJbkX
2skgIJEuHMYdIcFBqh8yA2JUHjEEIT83Z9OhbfWmGnq54SG94LN5w5yCARZgy94+XT2f4WMcT1yC
5zC/LVV1/kGEISPq7fZJuCYWZx8ElmE1zRv/1gIOniJxhOWwb7r3EKKGrEqGjkGtt+baLRMUmJAd
Ftx8DQTrOPyJ0J8JyHQxRDCApnOPDGVafr8O2VKF3iKiXDmWQEWtRdxUAd17olL00LQU6Dn/aNB0
7Lt/AngnSJ/GMoXSxqqa2u1Z9Qh26Vo7zEraWIOJRO3pp3/njF+EInYhB0df/PFMb6UUn3kXpEnX
Grq11xYqDcQ4Y1KYmuYT7wVmA0tQyIQ7sEMswqzs3q3vKYgDesaMkZDfkwQys+zRsedS1MbzDGMT
dbcu0JkpalXaOnNXu9yZKphnasr9Lu3Y1/LOkbt3v5Kgbjng/NG2YDXbkQ6nmDJNgyUlREzZHPy/
gKSj1ch+kXANcVuCad5/hsmlIc644h7GRhVkAGJFD0yaSxNmV9HPTFaxe8xuz0uUzk4tB5rnQRnU
MJdcc+EDokuxvZpvpf05UauhdOSRqX9V/a+1KlgwxSYPj8LBIl+nbTnKnF6BRNpio1XcF8n896PJ
TSetIvJHWqT72yzj0sbwxGEdGwYc6bLn4xeSts8yONXVboW75eWEyrb3wyy8f6oiK6GV73ZKisEs
7yYpbjO6FhkWO70CD1LEgmzPMTeKMXlspdYAK9vds9oDslrZUURgk6Hatf9GjC4hJJTrrxY6hhuQ
wPeTnRkRW2wegUTNfK9jCyyUW2/7MI1UrVerEwrNRqssVul6/bGgXwKQlKfsSg4zOg71MWZQf1CC
xQyDYs2BQn4IkbWnT4xNN5p+5WA40onxRAjgJTxE5iwMj1syY418IATsshxXPkYI/OsCvnS0YABM
7RkoIsnXdiKfQnkSrJQn4tMK9o5SBiOTcGqiB/5E9RtWoTx9Wb1fovLf6Y5DDiPjpivl3NBmwebc
H79oi77HYXXVfCZ3Kf7nK/llcWpFIQrkQ3uTRJT5M6ZbIl9x0X8e1Me/KBSF5TRsXDGKLO/NsVHa
gHZoLvhvZ77jo+HCoHBbZ2XaLFJ9Tv1d7aI7JR7mIvABaTvWLhcAQmERyyFIUT1G8+eaWucxeHFC
+OUrGXkHu+krxqQ4LOLHQCqfoXrDK0JBjmCLYfECgZ/gwcWNhaayKZVQmwgpHXrgsaG5C29UfZ8Y
jy5OPRehGUD9I9X1NBaRsdJZ8YdUYQTpACWZe3T5B5ls9e/dh5DQstf0MyQVv1WfV2wzriL7fl9E
JfQEXMK7Xh7ycXD7lYx1ZorN6OBqsdEsaKJegNQzYRukX4MTgA0/Xc/T5VgzS/bbiD8CveRSJUq+
g/tpZ5u1h/dkG94X+UuEcC47rFx6vBk5aswnNoIIHuIgXyvOQyHUCXlgAWRq0QCJ/XZolDfyuibd
5G4Z+jv9MKkFtMBQKCZeYhUN+rW0xJ1HHIKrVoSEP3tz34J5Ic2FXnVFPNd3ZLpfG0vJnR1xKoV8
Xzijlw+ltGlFuuKNKCP1sBZdKZaTxX129Ct+PhGAPQhpbHiAWGYf+OiDM04mrzVDg+PAauBNOQ1s
V6wajZWu0WjHLOJOaDJNQFHC47aJ1q/JTubk2paWh3DO0q/XMmdza0GU433gJMoYsNEwzIeG+xQQ
0I16E0Gt0O5PzWicEN74/MjPAHkIudYVNE8qxHd4wWmONYAW2xjkws0EtAi9QD1sZg8xahgs8bxX
wqGNmGbJcrDfNY58PZljwVGUAzsbjmeqQ5jmCpxh4cwoUnflbRsMA4id5DSdOCpsb4u1jE1cNHOj
KPcErsUXrYqGx6BmFL8ULEmVsa/KZZBzTswtLDTTV1kcQxCrn4vM9pxSe/TQ6iqPTkQC/K1XiSFj
6DBNm/ToOD3WHax6qwTuK2T1g54u/ZoZ5Sq0GYdc5N12n5Hc5g6vYtPBb012qF5Kbz2wp41Jafcc
cQf1c2ZIOkkBqFkHDJjTMdl+YESJzEXO4sj+O9IAiUU3xVP4h8r7QtrYyuKVKlg8J3Zb36mpD58O
BvexuspD2hGLM8Z+qAAVaWLQdLl9R0RurWqja1SeQ6DSlkzYr7ZvOMYlDpCoX7dlhLc9+yEmpQGq
QrdMnDAIvAhys866jq2TIyYKbov55bc3Z4fHrokNnToOtQX0gBcLQ6G65GktdQBrP4/w1yQ5/gkh
Cl4onIiOUE4+oVkAsnMgUtSTOu1eBE7oDM7hnGqxRV1cwTSVZhY6cVc5ObGOYfk7/HGfpKWK7qWL
UqZybY9iycGKpC/fSgau4qYfZw8xJVloCRrLjEi1cQ6xy17GDgAJUF4v4f5BfMKhYktxjYTA06/i
ghSqMHozzPtmEwYlLU9g7EthT2JE/TzdkAOQW4BCtnPSLIHWfjm4aEJ7g6NmJ3I24KnAgSmLBTEs
DZD1W1ioTiv8g2dQ7mj4OozhmPf1716UwwvGJSA7dvKmz5Q9yGGfzO78nUvebQLQPkG9LIWuS5tH
x/VGphF4In1XdO+FrzmbycXEZp7T7LRJG20BnZa8cR6U55852hKtKCzS90YfkVjKYx4xq1qA8ZY7
jeKTrX5fXM+vl8xA3CLUcvmWBvJoTQH/P3QGGpRoxP1Ctk3iwQVxKEAoZCAzILW+VN97aFlm4zPl
L5xQSfShcgIWxKuIEaZMKyfLUnH6ATOXBhYhkL4Lit9ois8BTPHOt0JuCt16NSxVN+FpGwlT9kro
LGC7o2+26Ma1LtIBsvjpUxv3oagN7s7QYlNgrDQe48oqB0Jm/0MJJe5I0a9lujI2CDBf3oLZOPQa
ucdDMJKF9lmi53E2TtEIhGbUwIYz6cvARPh22FaPjijxyjz1eMH0Y0yU8kDzOt6sj4btYnEnFEEn
jyYCrP31bUKlRHY6K5nfFDb/JnyqNSkUGHbrgKTHHAntdyJkCuoBNHor72wwAmw+lUW78yS3vpj5
01XUBDrxSa6UvP74BHFkQzU5Gpw0irNshnFEvrXtiR9hfQEzLTpzvZk4PhybX1a/Ek5KwpRnN829
/kg9eY8todGiYp8RfhjFVEzGYeviU/Lmjk53JhG/wWSjQ01paW6WgmRSmgTfcAa7B1N3P5IB6G83
WaRiBXkAKkL2Nzl4pN2g6aNdw6nM6DCHc+Elaey5RxeBzLeIwqiI61PNTRX0u0U3aW9YANbmkECd
Lq1fHq2aTqe6CgOqnqqMupLDsLOLiC/+fpX0XRXxil4eLCx69fd/I6Q4kl6ywtnMrRM+WP4tbhWN
/e7tzOzti8VGNIzJIGYUL6hql7LgdTfEv1ksd6wTG3FCFeRhYgoOQJA2nueyrXNnh/GJxnq14Bu9
Fp46DjQ8sugg2SJM80wjlARpk4vFmP7HdUMIv1i+R1Z1mMiUJcpgaTIoQIRrnZXRQyA3JnRULUXw
d6nBKb3kxBC3E2BoK0gsAFWHlggANz9yuvPgb9Vzvzm4iM4jiy/EmUA/JE5EP9pyjmrmgAbiTq48
d0qSUe5zbmlzwEK6p7lOgpJJjc9wk87HpeW1eFGs+SLE2y2YhCIing9urRWBdHyPXGO+0NhNErvg
nF7P3OPfSiUbWxPzRFrUbEU+Ii5AwONaF94HKW1lH3ymuQ7LP1epT4i5zJveSa8qRzvDfEQrXrGC
5ZkJbXJqIiPFusjGcLAxjBpcgQCaBIQyRGzS6uJTy14nmjccjFSLuh+u9WKdT01Hm/J3PfhslPtE
79J7DwXHdnxbAx8wWWAJqvpdHTrIy0z9GRCIUh8dl6OJZEJZxPfsZ5enKqRfUdKJx8LTueoXfx3t
5AdHfPlRfDuI6zuBZeg7V8Y/3/Sff1q2WY1cE0SqM5XRfS/nBtanTsijxi2gwAiNL/UQDFkF2v1K
bXRIA9LjyKAJLjhtR/6cHWeZgxu+eL2zhEFcqCKybqp4cyrk03SfD6W/+kQdgtBSjnfPh67L6gmK
bJth7YWbPzaDP+BVZq751Zz0T1tOVOx/xqJdgbd62huFwJWwFqIAPRNvG9daZf0y5pKyoT+UhX/b
Ol7yZev86KNdrwEUv3x04hISHEPC8kkOlSOrES6PCCPylfQ5JuzAJVHfD45OAJCYgdDOuEBeqIlG
fPwtQC+f0cKd8YhDHwrCbEihdyinn4gWnk2Vup4Jo1weadnRZoIu0mt6joOh7WyTIiYkl1bDGiw+
jeLPMpGV24rXTGayYVltvJsp3Uqr5sf7gND0YclevKqzip22Ak0jEsPwTrXCPdWwP+k23Z8Lz5F7
AJGqMkfdT2V/NofVL3tp1yGlMcMB4/s1Cn+jyAGuJFCqdvf1rvzHh7swv41pmHZETPu5YCAwBNII
YtPJrx4j/tr+NZIMjwD5tIL8GOrOTzPtZo7PDavMYcgYttqJqIFqEAGffo3N0gcGNZC5PQ06kGy+
eXRs44F++W4jcF2br2g9HXrb+Yzl1cpVM4G2We+aZuzloVAkDHHffrhcUVNY8JyWnKDYuOFHZBtp
nxyAUc0nLjiYZfNox5JCun1uGoGhQXw3lazpbdoySiGe+bKkOp5rC7kjtoe5NyZPDzZWRwZBdmjF
RzDFJ/r/HV0Lv9/7KblZk+d91G8qJlMwUhBiw+zCSWPb2xrIsbWON8db7R9Zaj7M3l2sKmJha068
UaKVoxxUIrATWhz/DszlyV55RttcBVPN1Brm0Zel3VUPOAWRksTx+5gZtv+Plzea1vkH0sETKHU6
39bL4Vx6AtSDyUkiOOa85aZhgW3E0csIb+Xg54LWOQszVF2/J/9YJvwsQwsiLftihpLyNcRPswGD
nyKBIxOrZ8UbSpLl7uKzf33BdbafaKxwrkmnAh/vDZz14wOR097suTzTW51+RNBPJJnVV2YzgoHZ
GvwrB5Zl378JLF2xkiqPtQWphKrBmiTepslEexsNDDcUycA/MfeIYH0cDYDjhIb0eQebX6KsmC5D
8fw3I/hp9cIbkt0P9uY1Y2DCbb1bVuQVqFkSjhKiQD2DBQkSfFAnj1/zcpRpyUyb5IvU9Up71PrL
U1HDuaVLVI1cFYHp1/UELj0QNAeRr5bB1nRFsUa1/GnjZX6NNRfjsIbV7T6W8M9zu/byGupvXSgx
+4yazuqbRDe7aWFZBFhT1fomGYhmXeKVFHuyYmxh9tDlJd74+nLTbH9yOgrbS3Jb0+DjNIuMpGZj
T1kNSjYjf8nAlvUveJgLlrFFnhGQET2RmdBMycW36ZpJ6AzT7pakTZaeWAma2GU2ESoVwzv7FY2/
B0a6XfFenrsEsCzNHvhbPddL6f8kYMaQWJsfUG6St53Q0GQ5H4cRZHzo/HxAp0woODE513gkcRIN
AL3PscnRq9RG6BixiDjvwXNX8XxH2af40BvnAP0Zq4wfdgQGqQoMBp6PdEKYCXc9/VSoRzqJJMpd
7Gq2WhKmYyZjE/k3+gZQfnHGqiUQOKbZSpRC5LKhzVpw53KOGZQGVPGZRviM+drtd+ZQQqfTdtz1
sU/Jsw2tFx5hoAD/0L82wlr5eQ+AA4Fzj56RyuKAKDxw27ZXFRILmLRpaKCTgZ4T+MT6KtAVibob
W9yo5KJLigUDDSo6mZ0waBtdp9ytnNHHsuGUFNHGrblEaBLwa5Go5qvIqipiwwdFiBSBzA2a4z+Y
Ximj/xHeLmVhwFICHSkWdKckL29HADTAVsje1JsQx9DxvCvY7JARpSwpu+lClvOSeum9FGvI0Scx
pLMLhi4+hwqTIAHBZC/46rn8ITv9q9jgeBoyZCnZEr3h3QaHaSOd3it1qNoM2sIgt8v4YqT+4LV0
LT7dqRXWzTHXAlxvzrqnIJhRhJSd3qMWYILnaawQ0m6GwxuWxNlvVNudqgF5t9DlcwCc81D653+y
7Od6Zzs8vtJZlR/wqEwXPF5KVqX3h4QN8Vsgb7QLYWQfF5JR1Cl9d+WnjBcK8J/ygEbof8UcalsD
t5mUOYCrXvm0rwubJPLWobUTBuB0Pl4o64sw0t6tKxK4MxJPWC5y0xFHkEpZsrBrI9yMq+OadBJR
2Mn9cE9I5rU3OMFYpW1/TLbTyY64Jxqfri7+boorENJuM52l/XdODRBu1i/7fVNNzanjct1NwQ6J
F08UkPYOMObgVu/tU7d+yDV2uQJHzpBhdv2mDQsV9JvwnHbMDvwU6UD+gDhvJd2KUgi+zU1eYMho
PIqcG9L2knHmTWbN3kovE7RALhyZMzH8egPihLN2tYjYonABGV0C7IsTYXbxN5YtXpNvPAICE4Ui
7CZN9EOAlsN8X3wMDvSqU4McA1uunbMKiRlcF6hQgUTvWzHqCoqvob6afyt6RjxLaEM46CbF8/UY
g2Sh1r7dAVerjh+uBHbaLg6+gmeULjna7KvnjKjOSoxyhPkiFvbduvOOp1kvBtx/81FWTtaIT4xn
ibGGd6pYjziSYmu7hW28+8jAB03cW95HAv6IKtydleehH8ufhlYkSxvEhLgvajRYZPHoINO3XAYt
h/BVeCiaaZH77IGKZ2dVGyY7pjlVDG8FVFb/0Ta7wOGpwWE1y+lei7xaXVXk8Jt85VW3NocOkezd
Simf+M4RlHYcjT40klL6eUx1b0XWuFEyxwLqOXIAu4qoKfV9+6IFLXCuy4rMRNA47SifncYNdKx5
YTgIjSSeAC+HGaTYBBOlLPqWFNI9miidifuocNKybNgJhPE9WK/oNvxXIt1cqsVUo9Oq4z+46V9R
YT+YbN2U/F2t6EIXZrG+YoW1TntaZVq1VYWlwtSeE8zxQf891JfvDcsEGtfUYXyK/1YlLPZkwVR0
IVhj4ctZ1EWOHEgIfKSZPmKT5vPjxqGbwx1RP3pzYjQrDPCVCcAaU/JKks5kVwe/MszYpbcZOXKv
25xgFnuoF/dBnP7xiC4avI7ZlWi60ThHa8sCy8gX76znb0c+YCG//8ooa6nbBWqIIAuTL8RxWVJK
5g/vnWXHCveOWKm70GyBC5ZHNJqQ8GHwoE2GaFrKCyyMi1Fu33k4+43z6J19/JMtbMSFuZFvaa0s
vNP/rZig/wiIazul8sZrsDT4lzwzX64MzQzdsiEp6G5NdPD4h0YpG4ZGSB78LSxh2thltoPtbnLL
gYz+zBOqVBElzCWqB6AKeASKtMStjzqUsjXrvhB9CT6BvYRe6fwuZuhNjo3R/iK8m2uKUYgBRqXL
64Qmier9DJoKCvaSNnNecbEQI8CHgtat0yACVMZoGu5PAZ0Sjt2KCS0iqtFoWIO7m7zvLcxiICsP
31yt6X2+4z7jc5e8PBgE9dbpZX7WCh0GZ2cJayQn8q2Hj4IlCjVPjz0wn3F60QBVRzro7tdnSxCN
4QLeg7o4rmlNgsAlNzfQhJL3EeF4Vr46bzdQ1rlr2YQx4RQuCMggqRi7WlMYCiDHrqchIVXA4fNH
YRlS3IMee7j313J9TWDzXMw/p3fEeTH+u1aXr8SiyycCjCoMIUJaTYP0nKJ1fAYitoDwtAjeZHV8
+U2dZYcShYo5u2yAYZeOHClnavIdOeYc6tew66oBHCkgB5qodNJan/3fv+Ba01nKAVyLzIi/HPNs
vxLcavoHEJvacOm3rsbP4DfawvrwREQcEKIZXb3odc3qT6C3ZcGZ+1wXjlnNhQlUY1gQcW7L2gIX
+2UZgnfmnn71H9zrFz4IF7vhlvkhZqvRcmV8HfTyAhIHr6tbVkHOyeODsmwBFW+HdpJJi8ZESeVB
2L/N3lN5JjTjpyU4SKTEbFyBpfFJJFJBerXngivCknNyh05gcCWWxLCfjy+SgPYkJFPF8Odg4KH0
CUa0FyTBoWGr4x+p7Fzn59J9zKBGZ3Lu10iCFomB6U7+0/pE7IOi3g4aggk3uWmPB3DI2eVjaxGX
sm0KMG3MwWGlkulev5eiWeIp419u7Dtf3wrfhRLXl+MDO9XUFWh9Id7U2NQ68CLPloYHv5V+8gqj
QJjtHjaOfE9Uf/JcPed3Wf2ZY+H57SqGHIidnzQ8BiicwPS+qY2S5G/NHdfcq12gqrzBVj9Hrrg+
RQue4uM2WeCm/kRA78q9QTy4e1ei/QTKvA5tetKxpRd46zVulsF/XtsmZQDz7NjXk/Y42YeSjG3E
45bzN6A4ZMor11uFKUQ6HXLTXBtjyBi1WXQvROclvZPVeL8HxAGBkSYgs7wDWlkWJ5wKuoUSWR3B
DkcrxdHpi8qBAqXDEr0BEwvFP1yeaRUGr5PX+k4AiWnpNikf5gWk30X2mp1H6HG0BQ1R+4uC1MKG
Jr2XpnXcc6rG47gkJ9YxCecnuRshZu5Y4FC60Zqk53ySPoagRbKcTJs0k3zGPIN6q3tQ+t0455lL
iqfdNg2ewFq2NPo6JCG2ieTkcFq4R3ltySbtYRb8k25VH4QjLZKKUVeLKOtdsavafvFXP81W1Q5s
FtRaOsb3ZMbpJE6CkhVyQIh+daDgn+OoWg11iT/lG/h9AOnS7iI8hoQoKJdusovWGnjctAK0h+At
qV9tbAOCBRZg5e3WcXiKBZEMfqnLezAFIOPKdJfRdD7CR61+UGnXIhr8g73yH1CRQ+1+9GhOGuI/
832UFUuKnzwrnK1sKuhkze+JZRFFxMAlmCD9tAsegyWP08ZQHNjuriD2/DKeQDJwoC2bXH79X0X5
iCaGn8kk8DcHdaSygRR/O+67aAdgUU8joBBN+n4lBF+1rf3R/sFmhmV62h/JmvzoawO4sv4ziTDm
QIJU/1eUqKtt4Q+eXMxjIeIf+9hr40svU518+ofLhJLsWHL0TzvxyWSxPFtZPDeL/eD2JdIj5E+Y
V7ewINOo1cjgCswEg8S8Z/rjIz+liqV2gexWlLIvE6hVNrmP7x70BBLXCTmYZ1kmyQpmS802MSR7
rZQpzPGSAA32JgRaxeIWvM9AB10Q6rBwUh/V0Qs0Cw30QPVBdOMfbiCDYHRZWCFMeKrMpzmrSAi9
9CXSS/GIHrKc5Sla22UdQKlq9+4XsCw3C25btN77QZqKlmv3u3NC5wFF3BJP2oyj5LwLeq2FWiQb
AbfPEKX5iAoXcU2BDIhvPntwU9i50IrlDpbj29wcc2yRmf7nRxy9ZWusG6ZREL2+cF9n1BM7EySv
J2IXIdA8603RGDQ9O2TQ1aDwLPcz5SEHxOSH/iR8uk8a1inP0Sx/MHY2wL4jJ6AsuzvIU44QDbAK
euBy2CkteE4rQtoy5SWiy81v7urLOr6Aek1q5ii1p06Z7TLZsxMTyzbjwGlxjuHXu+YBNChK5ZVt
hQYDDptK7ILkw4aGn/X1IGycYEbl9QV3irQF2GMHBhnd7wEqEY7ZjNDgxwtiGc93A3ybZVn96+qr
6G9Y3ViSndynkZydmAmTd/6tbgch0+fJBVh5rJvjo/mt3TabFtTbu3rvvlK/7iALPnFPljDsXE+m
KZsG9DcZoIKa3o4u7MqUbNiynLhjmID+ydFn3htVyJiaNfL5CecXDxCbEHeDQjKJd7ia/S2IoMcU
6Ek3xV4fNA/GgKVQXtfFirS/swgg/A+XljdJeg+1HeJ8hoM52FEKOD0j0L4oSt0GlTjCJwAvvx2A
9Unk7JQngCJ9czUYv1YR5p+czLB6lGIszStDApybYuhjjdV0JN0NCzYeA9gpny9RKJ2BeDPxKvMB
tNx7PfbADxZuk/mRVNH1BRdE6Xy/K4xOr+8uBqb/bkkMxQlN/GEZoAKBpCzZmRzYgbliQ5sIjNoK
ZX92Jabkb8C3nnvG5RtgCWtPn0xsAaUghARIViX8kHCm8Xfpw3ti1FCwKVuMnjtaSogbS5MJAT27
9TBP5Izkui/NCws9S/Pc150zB9dFXtiIk+GGGhjSZAhxiPugC40/ZH1o30TcKTdJMYHm/Sb8A78f
Gmchhufab0A8mTQ4mP4dEh5JdgTi6l69+N6iEV0SNhcd2Niz0DVImEDFk0doI7jcs+xaLnRCkfTS
1dFQ+70QpH1qj4opgoo+Ka+xWdTLi/ZLrNFD7f33niFYDEKp7iHX0r+/DRvSir+jrsJh954nRsnk
RlA60cl/WSNCdPn4QbeYZS7zD8h0pMkukuo+t1POaIptK3nsBBeuBNL+TaIDSQ6XIp1AOGA+i4SZ
s9JR9WgZTkRCY/FLIzA4s2y/6NRLA1HA9dZeNhrP+whokO5o6wSfMRZCuLrbpyv3sBphJjpJcqEI
w9Lu3gTLpwB0f1Nf2otEI0kVCOhEmwWWymtgGxexbzGqFS4CPAbEJ9WAnC+C4bHTKinbbDU99+jp
uBrnCq6qfO0U4xNEMxGn/kRlHhsHLeh7EB9y2gUpGc5xl6K0enBmyev7e/e2IHWWsZq+EBcFDtsK
GHuVffV6vvzAlmwbbocWLrHoIo5vJ6plkAufzPyQYQuiyyepdYpdJ6vPhYaWrce2ZPxGVNkY3i+Z
5CoXZmk46q6C4rFIuD8D/SbZOsojK9hW5m08Na6EotBSvuiz5ebfhhJFUxeeTUrX7USrDHBuuYLE
o8E8cgtNwFM1M+ubHeatKp0uQFELT/TEh20J0A3LBN1gr3lwBWRSbMh7+2cDvG7c2a/NPCPPL4zS
hEEHa4frZnixbWc1s0B1ydzVQxANNKpl/3B816TO10+wPeASU/I8SLIlA+eQDnyljekM+jj1JJ2R
TCdKjUyIs0TZfcSDWAfTSYadg+WHJXaDexxb1gIk0HLcbqpu4q/4+1M5DOERU5CqatQXfGHgThBc
Uh7+gBX08SLAWyiY4rmoMPeIomB0ARRsE2aDVy5hn/fsXCcSVYuqTPy2Xl+iwz/oFYKfOJsZRUb7
flq8QvwsWHfY8HmyWF1DClazqIrWl4mpEPZoxLId/iXqBkmBvSNiaLH8bjYGcgKwfGzb24ORZUSN
Py2pxSSoYRoLzPaoWqUrNLiBchl6PHdm0yRJCUwC4clX7d5ITppOa9gpIClyvhd9gb/M1YMawP0D
ARHBAd29BOaIFS8lki5D/2253QuYhuhSjodrJ0o0OVmEEo04iRcgd4RNM33OAPHRMgeWSzpX8uW4
MMDJR7T8qLp6pgRwZb13pkuXQrxrBnLOihO2AjQPcYJO03RxVptLBp9XYALktyIjsg4HKc7G3Gem
4ZZ6MPfhL1u0KPnkvtieEfAOKWMwn1lY5/rtZoQsrA9eCMj0qVWSOQQI/Nxulf9AB6a++zmWk42g
QR+Id7Fy5vnM/jBwVtyBEYnIDrkw9s+IHFKtSfGZU6MWacrOA2hsHnRVwUTaxbrLoYj6XUgXcox2
JEKlVJPVMVRg7Jd6ZuHLdFv6mSLXzvMB/pdJHVnV1s21MgxTL6Aaoe8I9qW+Wt4b9csrCgZ1V1Cn
Qh7dlwPfeoSTD3m4jQKzu1v9UMK2Zvt/3DqaxmjyTom26UiiaOc0MM6rbuNoupTw12IstBDxgcOR
9pxYwRj/iYNTCELBbGYnRh1r/tbLX7MKJ5vmEBls/ctJkRuD6K5xLNHKpzQQCftjX438Ta8NPwSz
KzXCKb+kzIJdavHDJZGYny30Y+C9igD5rTGolD3ar/47hXpT5RHTxH6x2p87fRHqW9aoGm800oS2
iAFgAjYvdmOhWHSS1/pqEPyF1R3bao99qrmCCt15euvXXhtSP/vub6qKNDpGAyXafFr0/y74Fsf8
dofe0Oo9BqJrIy9QwW7g03Ob7UdO4v4YRZLsv1F027U6GBpQzFi146yXc1KHfrg3qyGPukOeV5Hm
xRfZI3JraXTrgdefdKIMBalFU7XukmHnaesuiskvoLPU6l/Ll+asg+aDl87Nar4Xpnp1hshJWenl
ac5uV9VVzIwfF46GKRWf8tfZ8RsNAdC3Z4QeLHRlWAtZQVmYMz+xthAoYSc+070UJc7Ywg/KlRBx
TljrFmhAzdFoeIrmED2212cEYOjWrG/ap2RTKTNrnRTPNFV6GnE9j4jlJlrmiuv79TjQG7esxqOQ
KW8furmWoCLBIB/LBAmNkwb8Xq93Av4en/r8EGNi+EmVtUjjLQHu2RQAgm60Uwp0yS3cbN8jlBQN
ok6IcCbWLx0L0Mh7pfATjimCr5TBxht4n/N7KELCI9y1eUwZzjWpnglo6OvjHyktdQsjqvv1dN3F
6d083EG0Mr4v6epc3p6oZ2fDxZzN4fPX6URpZA4LHa38dZrbYfTVKb/w840bt3hzXKLqprzfvwzt
SC15/Z1ipMa8BgdD8dNW01WIMKlhMABfrhWCV/bmp3pgfVXTqbBPkiq8XnyGQYNg43cpZurZk1+a
iVIKKMREUkJ3/Kj6kWbPzi5w1tmgop4Gfll3WEl9BpX3q8jEtRlQt7yg2KqBo8jDylzBESt1AdOz
Ee5HwumGfgtjI5bv3ZQ2gIrZCkEyT6OHRG6TxuOiFbwekC6BKTj9it1h0/3B9WuhyfrkeAFYuXUD
TBu/zu+WRV4N8uARBo4xo4Y09R43ZSb5rtnDWBLqKYzQCtDW7Xhh2RGzulO7BbQ6Hevsri/Q5C4L
+EFnnnpiiO5brY/F6wHBsiIJOy/Y41L1z30BUk098rEy4I8aZa/umKUf7QNycDGf+YDZtth6bQrP
Y+2TArDZw8heqDwyZ1Eo8PiV6hzJ9PQ52S1E2mqA2EEA6dByDa7/3uHpR7uSvwKHDDE3Uc2Hqjpu
FE/ySpHw2PXU5s6Ngz2atNqLakJIGVfoySZVGGfaYeKFu2VrWupAAZ1KFg/h6ddgXz256p27nKvM
WAI2kXxQsJSGXjeGh/ETt6X9eqLSPkEsIIiBm764grOW5PLDjB+lLEg+vGdovtmXgGumiQbsnns2
ueRnwa2YFLQq0r6akhlAHu57Jq8r8VXzDPuJHARVNv/mrfkj3OsfQlvB9IQT87opSw0ox0vbsODK
IxCLKvICODi+5n4VA2rDpfXjRBojzmDKiH5/i3o+CfJPm4FE2MPYtGHD1FQq4jHG3lFjBv5zmOyf
VxjQNdqT7euq7QxTs77c58K4gK4I21+rgM52UxZfXml0gw4g75w4PajZevCHzRSGYmrY3xy5IJP3
UQtBAYEiEQmh6LMK1JUk3yRHYswp5D/Q8yivg17YdlBKVQSo/rUsEShPwo2ImDSw19doVJvOt4/k
Hu+vrpyA8HTOKr269GnzJJClg3j5CcA2HstSu61Lv4XB1sQAC++zxlPUhGZXZ0HjvVQX4njmmFuo
XHFbS8fkgd35TfeQBabBdF7z1wOA5uzeo+bqKbXbNaLAldoa76ilkkcsYn2YiT0BZoOdO9xAa/8K
stEGhaIx41iGnLNn3LsHZoavrFj0uocKHf51ucJ9NTnNj766ULYPW+v5/JDhjgyfh1rQK0ojqSGI
l9PQT9VTe+dSxKqWBF95ZUOIlNpo2xhG3ajROWkFMf28AvP+fU9vpU/2JYcFvQ1FeoXlivV6MwZR
6bK5TZbzebIRyv0M2RyGHqv4zZQ3QHKLS1wRCBiSrJVx9v9DqWcwxUM65tvfzmaVw6FY2+lLfVZL
IL7sBm99xSS/kdcmt+DECxRKXXSV2YLuhaXyUnWoj9xmYGKdcomY7VeFd7SwNcoXiTt2I5d4NBeH
u/U7gEN1vsX3bMiXDwPS5ZxJvTjn2e3P8m3rC5QeSw1/BJOPdWdPUbg9K5SezBOlqbxbX46MuB+s
Mj4Tnxtt0th+R08tuRkuhUrEjLFNXfr6oQbUGy96UUOaOOCxOsX557EEYlj4HC2/Z71gUm4URWNC
sT+Cbi3B1nqruePFG4dV5lihITqv1JXJV24In6Lv9CpEo3hw49xAZ9GakTmPQrOpmjpHAiZyOm+g
N8zYZsp92UztJA8Gx+R6dLBR90BAd5aFTzygelzDh7UcixzK5JkMfe4dxMNbqtvsKJCJuIbMOoWn
rjYkPZsnYFO0PEl2XJSgUnlkkyj6hFaAsoJXK6NEkwMEiytE5bzBcI9LaDbxS70lzk2feEO0qegm
Kxnhjp2RP9mZSDoRgCxy9zG75fpZdJAZdT2ORxo1nNP++2F+6XnkNYz+s9ynavOkeSw/nSFjAhEv
KZqrUVhLh4DEYGPk3G+uHfa+fMTteqm/qMkg3saUOaelBfZt1DOf1cS4vw7dK4RG8k9LYHLgw1B5
iw9/QjHWDS8XQ+sQDG1/wyWM90VTZIPUfKh/LYvBnfyBvB3SJ11S3GwGqgfuk/NuF+DxzeX+VLb4
SYtpAJZZeZYYodF7SbIaPC0iqgIeha5FViaecjrNofXcNG77FiV3jKe+BJLrAbfiSfqDp+Ru8qAE
wUA8XRQqNALJqMbpO6nU4HubtkdmfVeDgeUrF5o0K/1y5J79kjWBHNSyJiJPTLtbyJ4iWPvC5XqE
ohMGTFoC1iPLJ29oK5SKBYbq3V1UTTjpjyC12fZOyszu38dsQDRXxDl5XDkB95txBRUjAbaZVogL
q1q7+KBgq6zFktV+lr3bBLjjMpIe1Onz3QlbfBg4KOVmJxZOhfXwSjVIdrzKNmo5fQNj8tsvIhrR
faPgualFkgVqj+JdNpkV/FQFYuVKeCuFQhrxfYG6TPxbkClKQrWLgO+l+2Upap+0W+SMWPLI8xxl
66T48ZAOBsR1utTgydPD6HKbNDWEhkiJwQolZSPyHpG3bOG5ziR7LfHvBc3ZPqQqmC6o1DREaFq8
/tADo9pjwYeVXfbnMyQ1JbN1xENcaTAwpQFTufrjVcK/LW+GZoD2TTns37Js4Nq7lKZ6YADugYJA
Cv5y4XNFEOcHuK5cDeeQAjQfhBqRl94TQgjtz3qQilPL7HA/ptuCfR9miit4Fs1VVKv/ow6Qbduj
iBqFW1iwTEkXDJ0Q8lzETPYqzXDYYvhJi6bcmrEYYFwwkLVq3fv+g5NYqiviUxpuGobd6F+haeSz
8EYbh4MB5QNimM/E3MjhGGrKM3DOC5PuHr0nHwflo4rcYmW4pSje/orqmm0NUS6VkNmJBMIq3fpl
2fTSMpiJkXIyx0zEy0btbl/hvzFizw+OcLD4ptm+tyLmGgjkSYVNE9O6d8drpKisXwjx+zsz22/t
X1lKEAO2a3fM5ZmkgnTywRPbH1vMIgLQ6aMmn97+Q/DZsP0vWLWL7bg4+y3kJu5Zo8NqLjVdt+iC
5+Qpbu5tDcLgPpboi8yYnwk+Sz4MPn/ylEsgN+hTzsuCySAOWpLimSW5ZqnrYgD2SRhxdmH2bnZl
lr7ZQhz/hGUv62D8A5h5KDlg8aopI5mMAWxfX1yH9PqCd7ic3anmvZ+x0dJdK6cufcodvOMK5Lwc
WiU5tyXegvzBH3RDM2hEqI5q2/SsCQXbQdUBV+fUQuwVsLLf9uloY/HAiraOv3bNcJnQFq2ImYVP
QsYIHOxeLXZJ/VBbjV5Fant+ZqPfckBYpcrCBXtgBUwQ32HJIT9xrBMdu2RS2r15EXw58Ol7xqQh
uDtAH5mw7z8t+ANdiarnqKe1Es0ib2RweQR8OLwI3Euv7gtQtBqldOJm8liYwWpphvN/IiXil4ti
peozj0FdWX2KFZdeiQ2nbrVp+G1jcWivLMBx22JSk57374rj0IlBlzQ1hYehb3Jicm/cuvYSwXO3
YKdFq6G/RK8kwKmmy9sT7F+z2cndhucFBRjfJ4iK7SXh85OKejqIO6AhPwEOgE8k7lkmQxEijv5b
sQ0I9j5Qpk7I75RKqv6a/l9s50Za8TH8aHYk5DAS0gphgMfh+E/BceDNYzL8QIH4kLvfiPdCPEuZ
SO9NIhYrU1HcAKkEEiBh6hz+7W/27xs3K1a30mrWvC/YT3B8/Ak2MqVAwZU4UUX++V0EobARG/I5
5dBVhIfusgq8tQc5bDTndpKLzG1qSiLsN+KjEHjSa+O3gg/jZoJXoSSYmfi2vJeSWgFEdXDe3qit
etJD/ZoUziXCh1yNU9R2NpGJoiZK2E4xMw2qG5nqeeUOLDgERNid/f8oa65VxhyBkyhmzZVrNlMv
0JI/VhuR4WRTflQg2wXeTZww4ylo4mc6o9lYh+4Y8Fe5DcAziK2Df8hhh2j3XeTfPqBJlv4YaEzE
b8J/rbsPfaYSLWUpWYxMgddu1cBjMG7cOXxNObiQthBUfkSs3uLpHFFKXmC+zOMyoTCCPUPdCNzk
LLWGYALuSWrhhqduvbwJzlUWDgkRx8fIVwFEGt9Fivd7/I+S2BuRSAqQnCuht++awCk4aUQEYE++
XonUykfymQj2D3/Lno+n7lZNf4dYX4RLZZfKImPH0ciIjfXLg3Wr8DcIcfEw5GcHX2p/8/oMpyLl
1eRzBSktR22nDxi5ar1ZTAlZjfQF951ErKnQrVNe+bu5cQL2TbPJHrYM+n5a3mBJDSaPn/owSmAd
JuemG2JDBfC2/3J9Upc6SFahX7PbANFpJ9lkoPt6V6gsjfb+etNc9UzNPK2gp5jdvoGpdb6XojuG
aLa53ZOTF+rVGok2tgWSLvrJcX6/EVwbeJkVU8gwqkUhUR0OgSKywaQruDFSyeWNaYzM7TLHdhZk
TWODP0DRK1c5BTYet4f93VyxbiFwFt+Lr/0Ay5SlQHGFK4ulDfeqK/4XBBXa58nvH6WQUMiQq7/P
3wLitZhAXP1dno8xTTnhNw80XaDy8c8xd0djGrAgHU4lsBEnOdsGA+90fni/dJ/GoJSlivcp6OE7
Upw4yjIO+hjmUD/H5wLZON8uT4kpjgTdDsQdxoao5SjEG+N75YvRADrm5UvIhoIaQGG6UbLgWq9L
V3ibPhf0MvUKc56xLMlS1w57mOZCT6f31FfhWYAqu1QCLe2Akq9OjyMlGFoIrTSlbOxJBjGFbL+Y
APPyOQow+21Tx8O1Idmyxut1f5v+NMcyMpYHeRUxdB70mbdtPCy2zDWGOooG9nQOTrjbCOHknDm2
fgd8Lx/SNcEk50q7in4bTwGKN8TKvLGIxkY0t9S32Vn15Uogno/AJB5HyEAfBKII6fnZG9Gg0Wtm
C+ppygTJ0LjS3x/vh4TA2nKanwosn0yZ+DPYAlSvZMpwgulGeZB34W2sGkUvFuSd7eWDq+nxMK9n
ZX+M+t2dliC+bZ4BDl4c7KQKU4p7YFiEy6fsIvWuvnKMwO1iXJHNk1jdQjUgkBS2LYiX5FupR0ID
hw6fHPjOe19qCVmSbqUnA6klQ+2Fpscm5SynmqKQUcrq7Qw8iBmSve99+z2xg+nUKw0OvySIkfAM
eSeghIF/AgPeex2Pi7/kpVhgD8oTLyJRfGTFOXLTA8y2r9tFLd36ziVQAd1UkK9nStn1Jdx00jaD
V8/g3zglJIwI7aRcrSt4LR4mz3r3DoIxow02YpV3KEry7lBM/GKfGVEKv8a2VnIabM7BCdKkNmAP
UzOTlvkg20Hho1h7dmrknCEqpWWogxY3jpMzbpOjI/6TDcpGHYxOB/FhLTQHmfBamiCWJgZGak2l
WEd2OiWLQ87KrkNP7GA4cY1sGzfSXrx9awa4wKwdQeReXTmgvkMmZYIAKJBdvvYEvF1Pi6KS0JR+
ODe0lzJ9NdO5CExkzDPgEGQ8Q0Mk/VXG/SKYLJd2E4akeou6cFFo3WauKW6kfn7eKZPHyj3SRuGO
mTZGQRTVzP3SrimJpIVLAMvUCFf51161BCxghdkLFS4Q5iwWhIuFOITwPdIbMVKKu9UfK6RmaHxp
/MBx7FvFKVxMKYbTYN4kBa7m3zvIhUm6VqpAkUxGIP4hQk7DeE/T32LubP4ieAAkrZtYFKW6ck74
kU6YGj828mIoxgjdW8TTYLZ6EQ7Mi3UJhfmtW8ydXX7ijpsLuMA5z1u9KrAlaHopKYkSBhNGhGJT
6SKqun8kHyFx5NMwOhqHVaRrjZvpGoJM8HdDsV7v9ncmjfyhAhoH4ANVFtuC6Uhks2QVyn+zfs/v
GcHjLSMoDN/h8E6ZCsLKSz3RRDw3jdYYxspPc4uVIKu98YBHWKG5QL5iY2Dv06dnLgIfdU76Jkc1
2FSP/nfcQTleVXDvX3Kbe5/x8vLmevNejDSplxMRk8i7B2I9B5JoJ0eaGPVkm6ZhHinl9xy1tJfE
NRRcpIX2m2syC6eDCJK1bqutyGofd+AeTvu1JIImwfOtDUtQtNYsSH6e27LGjEQOMsF/gx85OySk
kKKTP1UnirDuglpOGZvJgr5MmSX/k0VftSjgTA5q1DKdz2wcqVTJdl0Mwk7aNFonIR/PnalwCnYP
UZXXecdjdCAvaVZHZW1sdS0tPQ2Q9mqyzRDgJvvx+hs6FWy23k3DdUgwUpBTnXU1V3XcEG1K3m7k
MFsDYSZGPOkNDgOLLjLo9dPKcIA4gyVqVQpJ8CL1suKiRzofxMXRXqr3DBY16+ndtA8StyXLutfV
GjP54MpHOA+OF0imX5tmP9HwexhZQ+pGojcLR7VI5tGQMhZI6pcNcFHZGJGRV2lMq12fCfRXMFER
+na0XavVhgoYmgJIm5doZDfCn39+/lEHldx0Kr6uY5nEhoxVSyJFpnpi2fsQauTJ6QjqbwIhsSXp
GC/kfUV8J80LgNgwas9xRU5NWbRQ3o2D+y6k78ar1UgCNQWDt88XjcOprZBrP2rNVwracJtJyW/h
hhZEbO6eCqzBZmS4hXCONHhmV3hKauIUeGET6YAt7Dg4qBsft374S+2I/sxXcgF9mfwekWBrpniG
1nWnEGTrEFThVrUEoy7RbHSKGqi8Xvy5jdgestg4r/cmQ7bbTFPhalAe1+iVryjSMQJCr4P7ZE6+
CXvMRLN1BbtY0OSG6kdFgggGS8miLwUm/EAssg7aaU1nxGHevhNu+k4A8JghVMRVdpumSZATspsp
XGJhYY2X7/s0zdTQeKfFk44H0zDKtcluhBLDgLu27GQAd/2bIYaQ4fHYn8q/LSWejKBgLWXu2qco
5JXW1EHdMIshDpmT/5UUAY32D69WXuegShscgHOUDKKKrOvgPf3cKYXvog0hjb+USXWgvChni1q/
H/EHSnGn6gAE3NKZXRDEh50INNMz4aPv0Clpo+AmR5a+3wGoxDSniHWl6qKNoscWINXCy9pzv8K6
umgUvvdQ2eA5fWp1TnJko1trepl3eddlJFrDc89nEz9E+2KYmBz/e/UYx+BhkknsNeIYhzIAO7ck
h+deDYPc7B3mUItXnYlpAaiuZHVoo1nnJEvic5fEEn3KfGEh4rCF3cruk7b4gDeZhjXNqQVzHmCo
bqYs9JCwze1o1Mm+vWoyySBN+JwnGxk4qjdhjnAtkoJf/EYFNovrJB7fEmERF4b80/rwQeeN/Ii+
efzWeEYfpEctm99rgOl4gQTxAfKBhaHBy7CR9zQLp+iVVS4zZOPEO+n0yOABPtlTgdA7dE+SMZ5L
tbRIwkmDmuYFg7Us9tmYsR9tVImsdhgvnPUW0FxxFw8E09aYjV+796aCL2WU3R2l7dqoPYeIsJjK
izr6YZa6GZkTpEEKZCtvx60g7vqT2enKHvMJE0h7RfNxuJCPPBqnoTpz02BGgE8svIEFVYHmnopO
aGWLGnYNK7+rDYHe77Pzey3Vvo3xC8Ckr2YzsT8cggE5PyO2nTCcfKGyWucWGjjWYotBMDZUt3R7
+wZ46p5qb5gXKxELjds31kCy7ZghXWBYRHoe7n/TGb9SLp0SLxQUA7EHYhA+WVeceaGCGdurid80
bpsYJiUgCoBzpG6vFWIZibhjtYYAvET37agDzNNRgZU5LWdh9hd5/3fKAfem2Wlf0BX9X361beCm
NXImQEXV5GgYJF/Z4TbpJ6fa0T+9B2+j8W7aoGtXHk6hho0IF7Xd0HEKzTdwPxKfIoYL6oNw6uaB
Tv487zQzLQarK6ZK1NszP9bKNl8XeKL1IyIEOtsN0W/jJpf58SRdu7I3rTKnTBEOS1Ee7lPlk5LL
lAVJhnjkVIIwrMi7v83VvlmCzgcs95VN3X5r3mqqChRsv9nT1SH1Zo8k/+n+/oIOcPOR1YiaoyV5
8vwiMov1GAcGoUe4NED7RNoFr1ohHokaMCeog3kz1IlsD863IXmpkAw2DmxvylZvVmAHG0f+wTh8
89BY6DrhnhGtMCDSGJVyYoHkB2RZXYf9Bx5Nn51PuDomown+AAtDyWu9EtL01noIDUXn6a/JZcXd
g84ryiz+mfU3xcHfJnltNBZ0pCQzNitW0yIiEkJJF2qsG5eX3ACliBEvnHpwx79rE9cuk7DA3uxN
wJBlbGmPAZI9DE8c7OAcEFkJoz3kH/BFPAlZ4czeSjE4aPhRFXzmk32o33LjiyaLJyNJux5tq6D5
4lB8I50RpDDJ6d+5EBwBlog1qTNts3Uxp7CT+sc5dkukPWSJFQiMk7ItQ4X25NPplroN1nnI6sJC
8xZTfWPp4OUH9uUlRBPULldO8cuiENn4UAe4VrLdMmQdHqsRvl9mzp9aQTF0RyLRu+khCTUYR/Z7
PTlGCXOD2qwu448Mm6zl0DjMwjYH1Pgdf1b7DwheelyzjMdsCGyYfu+DMnUp78LoBeZDl3j09+6A
j8N1MIkCkneOgwB6KbIAZupxJJkwgpZK1PGJMPbXxzZSZ/lSNcw2IxaW9UY0p0nS0uQPpc305NtR
WQsdeBnxgZjnXvP97DkYjFXqVygv4Pt2b+aJxacpxqpI0Yn2T4iLNwCQNF7rg0rotdMg54wI1Xb8
nQZpnV6pbXIYx2TCjjKePEhyBXPr1MvHwwlJC8zvNbYdGOfVORXSBEuPIGgh33Ihv4bXmPByJqDU
yiPtWN5FJIgW1QlW6dmAwxaOG3LM3trsszS+w4WdIapsQehLitQd3AG2KmjG5Q2sKSYoe41lPD+B
BiXDeWa9oIzv4Q1UXZWK83aM686Ghqw8I46/HO92+GG/fDLxccTk20i4lQmkKtZWM17Z40hgHztk
3CghdnB8/8qnlQxj1bglRLozz1vU05gdyiZofuAFX92eQCmJvNbicxx1lAXHepsT9ZUsy92W7KY7
uggdBHMZjgXxuw/ECrkQh3OzFXBoMwCxfjRp4py0SJQuNAPlendFVDoKrB4rR6oZhOJaorPsyYqf
uYZ5s9QmJlGDmkLeB/YW73T5Sn/RJY2rgM1ZDEFp3RuMbG7DTQmP4LA41/l7m2PnTmI6haQapc9V
MjqJrQjNCW2eHbfxMdk7hRoGtK7ZiaXT8Ug4B0CQ888mQzZAobrwaPx37z2SH8YR39iYytajsAEY
OT1VeFuGM006HPgBJ5ewUAx1cSaJWlfsd0MaCgklrVW7Dk7+Xk+STH2//xxgcDKDhXQTyoFGbH06
DuPLsxsRHQGDMRqElXMF7uAr98zfoxDJWipF1MTPQnvVvF4E/+Aala97W75PiNZ0zzyk0mGdoHkS
LX1qbP1fxirvntdDhKa2P0htEDohH9fTgCPP856G9Q7NTHNsZndsQfSj/RWkhHe4BuPS3LzpHVkI
2aeuXih0g2/BA7HUC6QKedqOygHzOAbvzq01YWsUR28kKaJ+DHCA/FofuKpdpda9uKudPe7jldE7
SnrBYJck441VJvKFAK4+C3yO2UiGOAyK2A1ozWrXFED83giO99V+0V47P2sp/ZyrFek3PJWnrP8O
Bzt7CavE5YskdR1d1Q0Gcs/5U1NWA7nlrFhtRBpQsNqLLIFHPoOHv0RPoutum0HDZfw0EdLeUcKH
AXyxeg3BurDX4uV2wkcUzRGFAj+I9hCKptH4mOJCCLs4SOH6KVN+pNuydbqF2JYMhAogIfOVu4OY
HaJN8KrO/RG/3D79o5AC1StWx6IZ0ns7361menKy5QNni6c5+AE7gjWom/wnMZdU6xHWwQ9zgPHl
d5pIHQkw8IQlA8FYY0MtaHqXX65mKfwMOUm70xKqebsYq8SunjuDrHTBLlyv5NWtGnXwdWAYzHS8
+VPk4DE1pCWVtENj+SA8NhEg+xZNtX2NYrcWqL2HlGN2vfbjQ1YYklnThmn+ULojbL72qAhEfBUH
qoMu8D8qwr4cKgTV/I4XipAbDTVQYqjojYfoLa26prphyWFHcc8bkqr0qrX0k5byvK0ZW4x+Tyeo
eDCu7mbPhY2Xhn66de9o46DACcg0E2oli+nBIYAc9Ow7rFxcXaJLwM6bd5alA6lBAsQS3LQAy0Ub
/8C5cossppTuNem0nNp49C34ZnZprr5dTPnUF01W3FxNLUmHKhRzGeoAfwWs7CeBpIorn3eC/KXD
f1zgmpkvVTVQgV2KhwBychIwtD2kdUe+cyh54XQwUOMs3qtIHfKLs8vmygQqA6P8Dcghfr78dbT1
PT0qlJ+BFMvwnTFooKIMXrwStN/k2SX/ra4Or4mFdlBMiQvLCXHlZkeVSvUpLwxcJnLTmU9Ft7Wi
OkG6Wur5h7cQxBq+ufYiBQ4MhaRURlUkD/P8/p4dp+GEGxSADhe0ofo6RYrTBwdZP2bygFvwOTBG
GCmyg4iLRETs5QTskexYuqswR3z823770/MAUeMSMOxAzO3rpJIQI569RJsD6XKKLLvxFr11InlD
fzAVDkAdb5mJgoAACcuKMH20H45RefbqxSJY6U8NNUU+wJvHbD7hED7E+t71ylLOhsG17qMVgo0N
fjl9pKVTMwwiIfgAfO5P+nT0wNt0LimI3aWaO/mVUrPNHEbQhVHK53CgXIQ0kKQVIoRp2NpZ+NZ4
eyn/p/WzrKjrhsQsOpO6g/OJmC81GKvqcouw5xfI5ouLTwYhgoCIuxd51wz/Z2/7yju5IAeGTPjw
bA46vCinU7W+i1XGTZzLyYBmjcP7qabe2hNPsN4qflWS1sX6qHxrT4I1iW4DwCVTwtndLURJSoES
g7OVXdwiyO0IcAhKmo+XgAnx4B8FsvrwxZHO2AhKEpvH9tKxmWJD0MmfqKEhaOfFptWwzvBFvAPq
qcCI9QJkG6AzetBeJLN/8695Tu/pXjZyc4Rm9JyQNL9TuMi3/aGTO5a2Sd+dMJGg6KN+n6GiBj61
VLPac0O22e1qRR9BfWEjFFJ5RAXA+/O58mBb8UZ2PPPIuWAUL6nmlCwyEkUE7yx9BvxJIh8cEuOZ
aog5OKo1Nea0hmANN+u00pSSBCOIkyxQSj0QIeXR2XVhhV9VLvClDvesZd11eV9m+AvwABcqeRg1
Hv1zSfZObGHmHTBXmAh+tSRiAQktJ5lY0bnha7FDVxvJBqf7Pr/d2Hye0kFrxYLHuWGq9xXMF55T
cbAi3UzH2no+sCQcD5Y2UasLkdh8HfzieFZw9SoupA39B8+Eu/QC/yf/TMP0RZ0/VPE+aw+MnEGs
VI+fAM9ZOa0cFyHZb8aktWDLuS4/PHDgsSxH+rGaOpmUuydLUU8+rZZ93pWcwZHSwu3yIei6Vz8A
xf+50WuaV0ktx2wVPtOcPMr8dTdVJAOJf77CtyJKPW17ALbHRoEwChwlOyPPr90Nk+7FaWPF5SKz
XJGqtJ3/XNcrEKV6gxgT8SftyVyRSS4Z1GnJcSzKPUCo2M51D6QNiDOIe/AEvBzsUrEr5SW6+j3i
fK1vZOuzgSIuV916OXJSUv+PZcxBg4tEtILccbmbnEk8nZHkz3orTrBNbYZlyrbJLvO9bna/ZJsf
2ygn5CXyoaxBXD2RMBpKF7l4HSEmfu7ziK8qMYz0bTAbbXaPVtrEADtt3M8Vhh3Rptrnj5YPlM/a
uhdN272/y8lCvfCG66UADcJ5ZNWHEEMJofuj6DtVlaiHIPID7yysBY9C3gNWOCn0AwG4tf+Obw3f
CICCf4L7YVjjjeiM1CE34yIVOcOZ3XPQqAXJ/aSE8cL0dtc8yJxr9bNQru4n902GOXOJezeLSsHR
KLaqNY5JTr29eZ4rYQjI3KBwSkUd58Dd2p0EwU0C2/rgQYrLa+h1k73+pPyzebRfWtfVOzQIk3C1
7ybHupCZbMQ7Q8rtEuLn+R+BwN1AniN8XSaGeWIF0X2VMUqcYMG5Tz4f60CnG2MEzwpA7yC5lnt0
3iLcZk89bwHKqZdwpU2X4YmtMrIdfSlzOxEl1S6z2Y+k6odzYBb7R8gEQUMq1PLN8MlqCUgeTsnq
T+xXD36PpyqXOjCdlltzMwErqPS7UTofdcXrG3G8jfXgQVf8qpX8DJeD1SkcJ05KfUyUAAaEWq9d
LXumVvpsZWmv0JDT9krqmBaxeQZ9cgXVZjXs736MVji7lM4TZ//N6gHryeBtaI40dcsnJFyODyPT
GeJO3l18uyBnvu+iRGcucFaQGXz4WMDst1znMhcGMA6V35jKt0Dtcz4rPHl9DrL5lcJOsK2UHz1v
5UFOzn3QkEJ0oODZqii0ay3DtB5eiFPdmhYYkT+p4xOY+o3l1nQZH+XttlkS6nFwoxJb7eNmnaWg
fKu77G194wA+0UhFLottgdVKO/aEI1Dqdyj6lElBCeXXiomgeNusOyUVrnYcmvKYO3kqXhFBzwKS
3B46hj3mbPs5bYuGOe4xKPtCAtvECDNtFuBh8wq+B+gNInogYjCRdf9ybykVMXgYq9Tez4ui6ITP
N7Ky2jiqcFu8dCuV9nMg0hcmOJmyvxvZQb2Y6w0QP5m9w+1faIb1JMkmTWQOAUtu01siw6PQRoQ2
s/ppQ/UabeRD1F/MX2fzaZimwOcNOHXWMZyfpTMQ4TRCvJ0HgivYNpl30pTVLegNXb6Siscl8oK2
tP8mhanhMw3fXuMoy+npoOuqlCziMcioPU4j1GDIJm6U3m+ZXXuYp28tI4rre8b577HJB03RRmPp
GsQNX3q54UdlqL1HYcW3gJyMAY+F2hKAgOgdVUykKy+ncQrXo4vYvKL6w1fI/wJpUCKRwfxNw3o5
PIu8BISIsASxZTbV147mSksg5Sgs6yCUf1Rl3br6i0OAQMtSlSwRCiHpvvTXm2Y1Ke40fwKNXLm5
U38hPG6CqIEPLvmAYCQa5TPCEoyLNmCVorkRjRmrAddFOxbK5g77wD0ayme1/jtvw5NP8f2RPmDs
TY+i6Wvg3JELm85HRi8E37CHfUPUXVDvst0X0oF1oXwkx5lbyJmTu7KRd5bgWVgy9tku0Oskjv8B
Fr1ZsCTgNntcw0MCWEMXafpy9tu5418lUunaJZtzC8Tv7VLAJCNRmF0uYBdBYRCIuqHECWjve9vO
9fwM30ZJyB3jNNMVsxpEvr6rYKqH4Obfd5Uyye9NKmcsT/TwRre8xcgKK6FeHost1b/Lp598cvtB
eey+6YE0cSqGWAYw/Xr0kPqLBnNdjipadXSE6VqEzXOEiL4zreXZIhM0+BQVyX1RChY3aT+dX/Dq
QDdueNhIbdRTq3YPJqqRWeQ00oayguCxUeMck/gl4YgxQtuEYHkndRc8LmPNOKmrJS+Q8ksEECIU
E5XAZWG2zq7mwHT8Ea4Kla9eCSo6UYZDOpnnW1V7aKjKUIAOdViGe7f5WIEhoGxTAOou6+9MYCx0
Xrpo+hmpILVYoKly8McWqx0nq9/+F11XmrBqxN7sWab3TJP9JOsrq5izM/bfXVhkYMf4dbeGseQO
WJkXIn4CFzXfv66OZ4/9tdd32W7WOvdUX+DFQ9UCqyt1aHhqLuy0IfeMN9HGxRKoiY2ja0cYMw3X
9fc5j9rGV5XytAuNghxtvz76/agV7jkDfMRH0kAxlp1c5WxuRph3Whdrf7nKhruUcwj7P4DqSboZ
dvQRxbyqFsnilp+1RyGBOiXns/GDWePgBwmSeTcZNhzm9mN5BKbDNdhx5OeFSTAk4AABPi1AgY0/
fUsS2Vh3tvZt1aXOyik8tMuErzFh2V2rvX8AMP5HYuTvO2lYShb70z132Gg6WsgsBK5kLitZlvzl
vSsGwFmubYtsFUiKdzMPgy9gup63rFKmanKjrXHPKY2zW2mMNyE3SunTBTMLH8bIjCLUpcSdzefN
XEwSMZfpruAmQvykRwun8cCy09CL3QkBawfhTtrcQo9sKyQK+xg7CMEWNTTk2dA32JNPCEWtUyPd
4B8yIF/eR3h4NBGdVnfwmXHYD8AxHKhRdO07of0s6hGNmok++njXwOq1bUid/NzXV6ECh0kzCLhE
Vs/eAfTsIbn62A/28cL82y0UTeKn0rZhG9WPdbC90cBsITk2FGEGhUdR6ZDKT9/Chre9j46dnQA3
fNK4HrOYSCM0gabRO7QcahYFOKgSGJoi1HhI8xuudADLcKY1AqOlYlkJfSvQ8PrIRc2T4p0v1xRs
TYXMPOqBqm2/MVJ6sHnZiyJTV+im1GLNl+ALkCLKUQgDQjEgDlQsTFvSM9ucewZuUrcposeoQqR+
3SlmCslJuAYIzSv2ZkytJlszbHW2PyecA2BAxoAAXraJs5qCUbmE2fK/eKwzma/1hbEGT1A2wGKT
N6rKBmf1YptULGPjcWxY4fHQBY7rD2wlmU9EYDFUJBCmSKOeqiVCYYWz5IpoaVsVRxA7Gv0LRFwG
O/YF21/FgmJG11KEzl1csM9Tj+YB69UkzKMDSk7e9eIKkMrV9czNIviZnbGPv322qhby+o2wgREh
UaHfMqfylYkaxavts9RsxuqOF2ONZpd97WMWGp5JFfCEO/Fs8QinjMerK6of5AgA6zskjizIK0kI
eyFFX8k1EfnRPSMuROExdG0rszh9031/WZRO1CDLaUg8tA4JgyqoJTt1EktBQ/2y+p+zqhbWEkes
BYKAZwJjYdGH1mehx/OtAsjI+2etyayx7ATj+qeclS2IWvXmJHG6sAiMq3eC3neMgQ4FZ0TWCHSU
/wsuxdbgR6sxWIhy4SteNzYZM64iXUB5H7ixN31O7xSJPs6FQMwF0iXZy6BWyR/fdUGkDZP57gYt
l3MPSBbUHlT0ywVWpQWXdDc4WKNz51MLQaHWSQBUJV8hQ6aTyMN4pK9A/nhvJTbeOeq3NHHh0B5L
QdHX0W8d2FmKNGaLvnP4McKhrpVmeh1y+jpv2poAIC5Y3SS1v33mBzoRQoo06xUZmab4+od3jY+R
Qeam6FFfKbfOiZymK4VqcC/HuJH93KiwC30wX4WiI+bcbahb6lagjwlWoCmpt1t1Ye2vn1bpeCGG
y1ZSxXToQGNKXCzEyyUMyYML45do6zsUEaXxf7KZucR85R8vhRmZdUJEXk2jNB20kG7JctKor5jh
nWEK/QXdzVa6JDnJ9OfCH5voGKoX0eC7NeN5+r1u/mG8ChcYKulb8N3cqYqlq6Z2QnfgGHdjN+bD
PJrtHrzsDp1byEZMmBzMigvmMWdS2DTlfP0bagYF0YOQOsiUCCJOi04kcHrxifTAJxlI4FbPnFpj
WpOq9+iIGuaNAp52SUVZgtFhtEC82WScZtiwtYZu9ZkcNhGvC11IHB1czAu01OGJEihJeebaZqjU
0xW2frN9j72z3aXRuBMYxhTvxFtngkoyzDMAvfskoSY7GVxwbHIWZKXDkk3JpgLcdNhT+9WDehBp
mOthfl0nHdhqdEOb9hMSIjZGl/pPNVV2LWEoLx827QbZmnLmAHC3enumiTwwx/2bTRP8jYr/uiTf
+O76jzjtEj1eJXQOHjCBaR5eOL/+3feNsPYROSW434tL9VV7pY4j1rYF1k3JeqcVujr2Zx3SJt3u
odhZ9gCGh7UwLR+m7W4vafA2VO2Jc8aAczU4TWatL68A+6Ccycz4sUc4rOpeEEw/VXaSvmo2jpzO
4EMENNWrLiIMosw0HeVuSOb6SDkZK3OgBZy/+8FzR//tgO0veLCrK8zdhtntEYqJ5BhADpi8KtPR
j8dBx8kzNuARQasiTNNj0rixOzge1eWKOfiYBmIzhAqEZMeKGN3qlFsH6+kBJX8qyGexgv+Qmzp6
5kNzEzzjbY0hWl8IqnHDOD+vwjj1CqDjPd6Y7PNlqCAN5iYBduqPThGoAdPdvrXnrORyvbcmM/a5
4GYuJPOd33dAii5CBkvEzdcq9flaaIFe47u+HKbWhfMuDDfYlqSR6zfGqQ/lrSYNrHhhdsaWeHXy
3AG0KBGEIa7RcD66DixbFHJcNAqFkm3/D3mK6mpejwywpLiet6LXTVlp34s8b4jpPDtSqGjIHBTW
43sCCZaTO6Oz7GyMDTsq5E5yhL5AMNkERHou7VW5nJCcPsP0S7RHhNNhx1JvNnJDtsVn2le+wNWW
E7oH45DgVchzHPKg3LibfFgLzWhqDmvcRnfwsDJ7yUXjTI8y68+dF66yjHXjJbMBgPO7IclbZdS9
VAV5R/ZVnZGudd9DsGh2sM26ju7/iTexhW9vKQQH9QSRVGsMRoTEsqucCsRTqDb5E9Djkcd5a7Ct
WZR+7qY3OcLMVSWseXTG3WiN+p57AstdrhFHsEeS3IkP/VsG96xcroW6WL0k+h8Py9pohTWXkqk0
FD+92X53vDt2dyswzdwkRZOhZcemYARP2cY/s+3yxT7SZM3b1rVuAU2Ziw780J2w+4HM7JDDL6lz
uEdnin3XBTFd3BoZWFli/nOPqxPwyT4cuJYDFeMd74V3+G/ET+ufoU1vN5500hm8p3XtjR6Se8rj
YmJT8eSP5VH1aFewrUQn/0DmT7VrMwjJp7AWqLzua2WsjNF9VQ3D5dBUNGOZ+xBeEC5r/G7hD6FI
Z+vDOk3HhB6NNtkSVxdu6GDtaTMczSr09updOXDfcI7pkkV8hRw9RZr9DBF4J31EhTHsM1e+1Y98
zU0QjN9HKuwgcwERYS3i9RuRARIdFJqjqei+Zjsa437d+Fktx0u7GjiHXlFS8BUEQxO98wPsJ9bz
3Zw89zOle5l5JgJF6O4svrprmhAKWtPdM1uMQo8W/XK1YiJNVKLA8KSVTkDdnRhE63pw/4FgxLur
TW3Yoc0yASzHK/OCELY9R7RFCPyrbQvzVM+dReHfQ/21Z2bbvDvAtMxtPUxAZ/JpDEoG+LkTanWP
KNw492AtcZlYZ3CVr3+cJs601HVEHFuD3eUwuW6I/h6sPwGPvsRaW+dBbqnKGaHOTcq8Myp6w3lR
CVqy28dVvIOXj4IWMv6i1E9UvFTLJ1y6EEsXdpAHqoYilfg27itapgG7A6/pzfORUfAIp0sl8zfC
HpHcdYTE47a6fSxwRAW3gLAqsCshH4K0Ve0vpkA0W9kkOVThJVFRcz7+qzelexaKlw2Vt95z7V+a
gvDgwVPuxzgSSzO6AtvbA2SUpXE5LMmp60Bhm8cnUaXM7DeqMgLf4UYKh2L2QZG6nA9T/6ang70Q
hq/p8y8O6R85Wpxn+0EoOCLOeWP3UadNs26A48bVsVRiKNK3pQSSlh6SORAfHFw6Nf4ws/6f2I0r
80Blny3y3gd8gREF4TdI0B9CaKY5ni9PQrG+HoPW4QD2AKZ+0Wr8iwys/W5me7oIUrtPUKuRpcR6
mIkIUqpRRlmvOAW1gxPIBRloCQAo0VNg6ahtGg84NBDSQWCkTK41YbsfrwPsAZy+KPOOWivsur5g
ShwiE9cK7VXNF58wkGYYts9MoWDN3kR6N/cc3i8UxhZXdAa8zfdpw+zNr7gD1RQdxast7jPlJYBn
WGFiZA+rfUEEqaSjXpS37UZt0aHLO6xwM7r6eDcxCb+S9ugID6AijpHntjRFNLMat54d2wLFyXpM
JbGhjCYd2XAAaF49WVUQ0wQV3pQjBpDH2xW3LFlKvcSqpgvn4gk0uK5G2gFSSGHctGeOwyXMY5wX
STcUB8VrzHaqZTkw05BS5lCCH9vj8S/8z3W22+1p6p1fRTqEkcNVZUrnNWsG33/OdMBnZQ5vfEkt
IkiLjYQuH7jL8r2Yc24V7k63VtIC0TcD5ZqGiiZz25rgxwgDbi5uUZigcpB43n4nnmLT2/57n2Gu
QTUvI+af4ipo9z+U5ebfWniuAMnyMp6MA0ZRqTNzlufqehuzDty7nDkpnJlDq14pKDGrcG72PgOV
6U/X45HPbFAs+810CIb2LVFn/OT6RiTWEXJsnIusdJ7f3kCCMGG4edASkCqOhrmrULil8UMB4Zdp
6DAoCFrh/VNHkx8ycXLGqW9Vebp20yAe8Jp+DQH6orvtMZsnWBmYbPTxlEsIbrdA9UBhDPgmI19O
tZaTcCdN09IDznu5aoRSPdX7YEcFPPI6aID2XsC/fLdOEaHAeupplBwjZPbyElkxAYuoWIKUP6NJ
A1O8W6xdglQzQn+OeRln9tHW7r20W9o8D20WEo2wO++tLyOw2Odkgc6MtIjE9JdcvYX8zDDQzClY
LA4tHJYKQeyCNxyoyFLPQ5kfhVxo6BXVZt/vtAhyPZUlVnPIHbNUrIaGKHeYMeEEbR+8lMjmrnt/
1AW6F7DuFDF/obd9BhnSNQxTvGJ8VkKmMQR0Lan5JwFcH2jzLnL22H7zK40IC07D403NDU8NvhaW
xyjVHEIGcxvVUTM4jul4HlRX7cJDIL810pMkcfTbaPT8XcoT947JdvFsxsJPKVgiE+ULqiDZWkHY
hDVrMaJsZSUfYORVCuKnfaGdE80ATvCHeDKDjxuQLRUcgCbvBs+eUeJVVrD1JaOepGXv5uFkyotB
oeLsUS85/sZHJrPPehIZWbAcAXb6CTi4/7xggQ2so1zv+9b6RLbPhFhEnloLjjb+7b+9lCmtZtJe
/tIp66cMru3ETDVA0WtDatcy6A2+gvOUpLsSSBW1rNqYgbXlipF61P3W/qEboVIwdo5vMwfKIEnL
FGPitUTKkB+gEz18goxPN3a+on2Wa5FE0MgkitexCFt2QcihYaLu3R8riMQdyDTYSkzcY1GLUktB
Yz2MQKSS9cIvk5L3i5GdHuvHM4zeLYHuCdPF1PGuVozj8d8JxzGrNkLFEY+cglKgje+hL/VqpPfW
rgZA0mKnYb/5yqrbgvHpkUBEmUaDItr7lNFzPIwhJUCH75CuGc1KNus4GxehcshM/8q6CWgUOCLs
CejI8+qtj83bo/l+Vr2RkX3jMJklF9ZJCOW0VZThjRm9cMPGlSkwxZd1xEW0BedZxoCmuUwUXKB+
Rik63QXd3weU/MRyeHlMlU1bXUBuEoHQsf2QrIXYvY+52EIp8wL81Bjm5OAbIDFOo8saNqBEfqrn
uYvMRp4KU6th92ttZiAgTsjySibp5myQ+wR+uWucersk9Pj59BBCNjYt3aa2ceBKJC22wpYajmXJ
h3A7i7RraYfLtgq3BHPUZLL+mGz0d1b3Ge6v2SR3FTLN+IFokIqspQnwS35+MVg/N9P7UwPjm+kS
phgHrCbxoP5N+FUmoGumwWa2zEDrl6zh9I+rJjpmzbw5HB2vcg5cbYO34ZOFmlA0M6U++Xw00Eaz
Zw5xDD4dwz4XoxgwqTq7D0Su5RhiLvhGzlUFaFmX/19z7gjMW7VRUSG4coAXc+/Ocqk6wJNyw7X8
ABEDbT34Yvk52EWpBNjovGVCfEldv83BPFppica0TuKvgXsitcEHiWofYegCpI7/hPTJLjAtmQLr
+IU7DCg9NYqM0zTUQfEjzAv1uozhI2yaPJhrr/39dw2p1lG5w6wk3qfC6aS+9LAtcGOwTJomXlch
adym6mOEVPoYub7LspD6lhg4MRGDFG3n9SDunGo6nn09+CKbjuggHs4bfvY8mffH8tOgj4LHmPdT
ZdB8L2uhc70N7+2i+gcnjTkXJQzSMU3KJXyP+loqoaVt4d+H5KGHTvtqUtoVL4FigzjBWC4cd7HE
/arTbh/qp4O8H9Tnqnaqx8XnOMZttLAu7aGfptuan4iFwLKrFpBU1BsAk+Snest02cFgnoaIzkHw
ugjJqO026G8yR3cJfA6mRlwb1tIpk5LstMILIErb6T3KVTKehUp4Ib54G7vegO4FlYWlwfTJ3A2k
2vONMHj8dtlL+O9J3nr0FuV0kHMvEZ8DHDIgbYVb45kgoW0JCFu+bx0dJ+YWvQJfw7LOuAaIFKyL
C8HKImkd/JVIiO3k+SN9ogT7pbBb4Ee+pExhb4YxaAXvcdy4MNAkrBAuPsdiLkdP54kEPCN7ZWem
WeDk+eEzd47nhy+H/qW49eAouRONBU4WD580lEv6hh8muEhsRgGo11S5zC1K9E5G6Z1dnDjzbKlZ
54i59bKvRGqYB+iO/gzQqQ17yJfoWB1E/C+ohCilestpOUKOtHlAF4qh5nPZiy6sve2HAxjmykAX
a4Msd+kDqIWgQkn2b8xI+09UXShoAoaycTJA0R0cMyrCuRnDESKMP2NU9SrmWlWZmDKumhRs43F9
12heSaotrce44BUxT7FZiuoyd7kxAmNptMZCmvZJw5o5oTNvDdopItP8h3WWFW24ZW/U0zObwhsN
5/JSFzF5qIzfQhOD51dCV9ORFLjqg2WsuIsmLSDkFmQO9ZfZpCCJ9LpZ3xGqr2/GD4P62J1b4nbx
wBsV7SPkva2GxuBqc3S3I1Q0EZaNhEn5HO0kjInZ1pPbMb9yzM8PAfpEFzJV79NnfK5nCpKTIViL
RaP8kLQDrgEDie0XO1J682v01SGAN7jAqCGoFk7ZswnHAXt7PI6jmODOdTFxxGVZQyOjpTosLMgI
wh1OK+h1URUIcS3aSMjS0684bCzm2LmYtXLA4oJyICM2Hat2vz3xvaNEHCnt/cuAJ+HBmcgMlj1O
MNKROXSNIx6lBQF3TZ8p+cVXZooChnpiHYx/Yqv02K4u3UnPfofoxqx8MsLfI2YNfsxV5VE3N8LK
CEueXHGFF3VsMvNJ7nN3IgKn4ZidAtVeiUWAuck1ln3it2Bje/m6OpeoarxMEwWn0vR6L1PLA/v4
fCzAxnc8YeVT9pJ4LYGERt46kJoKxkzl+HwRrtfHQfqvZV2A1qtQwMblep+WwVADl2MYqPHK23SK
k8WXTGN2va8qoVvusjcu+zwcOa3qahBVBTh6xqeJxMy7KBmpCqvj6kj+yUloHGDnVCOx77XexzoB
xFJM724ZQZGolrVGNWFwrBDpFkc2Wb2J+SeU+8EbFfuU3cEIBmxepgWlWHBkeKWjDPTNY7ic4pUy
GeNTxyEj66X6f3sW+/yYD6kfadOp/KIGjhIUQ72579MhnLSz8qUVaGjYcvrefo01FZpfJ1A0s4kj
8bjeJqwK1rzmGIAPmJfgYw/kx9+z3pQpcHp4jBiKKVdJE6203ClgeX0PpkTuNgGJwCksayCtZT/l
XO9ueVWNm9UYMKQIAMvepAMrO40XhEQiP/WZBbgvClIhfCzIizawkXfakKLN6qsiynp1oOXKWym8
ennl0iJwjIke8BDh4+tFBbXn0/8Cj2oilmQqptPK+h96hn/VnPa+9AuDTErT8C56c4NXQZZ/jf3M
UMPL4bIHOEgIQlrVMj6ENd8BL7cBgLCsm9tKPVlbdYYixsxk1JlvIFxVCcTJ1IZz+W7aaU1OYum6
nORDQV07zbx5WNjr0+rg7TVSL7hY+9tUl9AwQE0rxYsngKYMkl2B0Zz0LlF1kPgLQA4MkUP8foiI
QJbegDf6tBzGCXqtBU60shtZtiosvru2jKNOmrtfd4uMiGTkVdru0odrkKyE7YeUhGPuZDZ2Zdzn
W1BSG7r5I9ZANq7V5aI3t+VIjBH3dPG2/A2PON3B1I43tCzafIPccxwSVdUk3QV+JFVaC2L8nN5C
IGhxWQULi8XJsDBSiAxnXWlSBsp+uw+qCz41Q5x/4u9q0LXWstO5p7Ky+HN2MtNNVD3JCyM3z1sI
nyl7ZhosmvEnc5cy3si5k4KS+y4mw32A45BUJqqDGpLc7ItngBUBEFI2ebmX2ZrHJSDaZRbKtRAF
sFniyqdyBiw0TDs8pqqhX9F7cX4CNcP2FrIMPNhEmKFI83CsH2Akf0/1AbSjuqs7UgpIIkClFSx+
Z+edCiv0BT22mxWMi6j2HJ4NwsS7LE1256nc2Z8Rm2rjE7iIJJjiXpS+5e4j+/fDFBG/DUHLBC4Y
PhcbZVj6s+eb9hd7wA/4JE5fskaiobCDDNf9Ub90yiEnhkjqgqfU7DtCAD4GmkjdKAjvGvA7SBpy
gKyT5uEnW5VTUR5QArrGHy/wcAczqpd7tlQr66e66bjYRgVx9s+juiNGMAiUB+HueODSvpt7/iS7
rvhZif2O3OVktV0YZeQEU5LAgvuVQc9C5SxXsabnlpW+rj3Pq0abD/y8ObZmOoLqyvS1uKoNucy9
CPggfMa4S3GUhA+4RuVZNZYZp/HWt9XsFlRk0FNdIg0JvVlCT3jeP8V6f7JFUoGyZMjYHrS2rxXe
ywxiPwAYr54a6dr5dQ2IhCrVZcZKTy3dT0yaan7yLLUlZOWMCFz9IEOCEa56C6/WguwOBCOs18a6
jCtZfGIiuxQchsK2QoDo61ksWcS3jDsSNhNG3thSVN6ZOkcNBxvp2PNQZ3W1wiLNatd0EeeP/kjb
tRm2wUaZ6NG/u74UnM1Ckz3kU90Mkb8Bwn20fC6k4AgrDpWY7D3HIqCSHSHcEHopBsDzBokrFOdX
mjZpEv2EtYi6eBcZVxk9uR0k2aGamo15zO3XoWBOvuNwlw9EXQHQnISxswWcREwC+h963otbieIK
HUqunB4g+ehwdl6FnJyQNIJyphnE6bqn78OdONaiiQDj7rhB6dhs8NcZIfEzIZLJpmm20gzdYcjz
ow4mMT9Cc3CGdWUlILDRaned6guagYj481IpJbvYFTrKGjar3yrdBFETaboUBKenlPWXuC7DRvn2
C77fEWmrwzr632n0lnYlPIIbanMPBUFdzUQeuu0VtvJcNijWAhcMi4nhPtucIU7gprX9HxWI+Z17
RkisFZbdZRJ3eJ3DAIeQjxF/ZW1fn4gIHiH0yGrIbZ0OAClsz0wAQIIy8zZ+Y/wI8UvYtPnoWM3u
hgAiKMtN1BBcpQeNWwHj4NgosJmg1h7eHJcYaznr6qpS3IQYYqQ5pjMTE4rfiJkiR5P+a3JBefhj
dSmZwj6lDC0IqIc8HDxftSqvVph6N7ihbhr9ekJWbDV3b++z95Wf4z2WqSr9LQywnI2JEkYsQ9cG
vX5sUNEw6PBURGLS33WGF610E2gyUEGAh+huMoeC9+rBArcWn1nkqsXsfPQAYfrdZgKC1A/7Sst1
QbNzdY2Uwae0MyZGKn93oRI+4pimSxV9VyjEa06WPhn2aQcNHHAMrBrsbCm9Sxdr1dz1FR3IR8pX
f4m5Pt1S8h3sv51qF41dh2k0WbKEsTQFY7qDxGAHMfvDOW4klLdJpgst2M9WziNmkyueQ4nDuqUH
Cm3NoqJ9x9swk3ChWQj18kZfsKYKFCRjqsvVGEOZnvVfl3pHTrvP8CdZif84IjvwGw+KAYy3fa4X
w4KBuUD4z3RjhcoQfcqab5g5TyaLW3Kcm+vVxPNKM/zm5G/0ec1GxQylMrbprpE7GI1ChRlWkuDO
bifWC0lZ5ZPuBV1EkhnsIVTCno6x8K92y5NHd/C9VAYf0lsL3cjHSRSpDqJA4BX8L3T69zfe7WNF
4d5rPJ2Lhnulzbpz5tqdfbKup+ix1aYQUDCv3FbgyFC4XlEAdzZG1XbU7ZFijC9x3wCGkSlFn1sn
z7yv0whzctW1N2IiK8fPXm08RFi4/lCTPhT4C6FoZWaullc47USezQgibQkPIPiwDL3KNK/CA8hI
YJ7A3Mx3D0LAuiObCgX9bmgVqQ6Wnjdk/QeN9971IX7+Udkx2U0VLnXSZO+1wWqQh/K/cqxLhKCT
0cgzU1FN/kIEGf5TLp+CNYAu2+PLlaYorSUIlrpLvn6POUO7OZjTUeqBIq86FydgUHrSf1HPsSYy
1JZOy91CfBWKQfCwVJsU9fr+kTpEqHFu6GrO8ex4Vh2ol1g8pI0/Xyrg3E28bNvP0/2zVNFuy/sO
81Y1eTT8C1coJ1uR6/k0+9xmiplJauWLwpouZj/lPJfy8SKDWegm8mdvgKz1xXi9Lc0YzZTJf1Wv
rBkxunihPnl83muB5ZhgTvLgD/lqHjtKc9Dt2gOiJZVqH+lSnsubJnedv6eZGZRYR0FH4o5RXJk2
KM3/fKq1y5U6HjcttSckAkPs22OFR3hz1i/xp5jhd4pIlIq+WsdHWQXYAQeEbi560lTI/5WlEc3R
l9493hlVP6gfusW/sIJCqlItJpvxkMwoPFq2EP6bOYZkG9qOb5/2i6n7v/hLnxgzaVSeUmDP6fX+
YNx6cakXqJrsGwInKJZkfBONLv6X1e2KM647I43evhUCyr7vSuSCJ/H4pAqbZfUjMprain/z/4Hy
3f2EjyMGCBx9gjb4tb/lsBMB8RhCeDFH7swP+HGW/PyzZHHEl/gj1cXuQUJq8N+3yBMuTKqWS22L
2CvnjcvwaET2/3AfOjNlCEvlsiI13HQhGK86VioUEZgNCRfVPEyGJC+pJXQMJhGcW6jJRAiKbQ+c
dBF9+1xtq6L3LmXi2NjurYvHvm+LbRh8Wm/wpa3ZE5Ny13wE4142mps8/w2ihrgngxPz2WOsHuoa
3pDnBnV/OONiM0YoEnYdZ4wV8ViHqrC/GeKipGoKCyjJJUciWXm5zPDuyr98S/jDGt/YQKHqlR6a
udwszxWWCiS86Odr0ZsYGKKOZc/EAnKNyEBQgGI9Dg677HlJdAvmDHOBOIcXy1CbR1QDUCI6nzq2
IqC3a7OCaOf7fRi1zgkBTZcHYyXkpOhHhWNRefj3uO5wqWrnCjbBfN0PlAZh+wR6xakzZwdHtywc
iwxRqU8BgiB8bOm38kmiXb74ahCJv1OnGMHaIb7PyndhizSWluLT4Lbe26hKb1w2M3o4Dv8iN1ZS
v0kp0xMyK/SYZDT59yUUqEAj+ZtPtzMxPeNvuFvOwzc9/AqVll3YRXd/zULjyf0vLKt/svj2zDsB
HZdHN/EcB1HLSMLuR3lrytbBZiIE0AY1ysqgWcqXHCiA0YDWCyNtm157WxTP2eZBi0VLgo21/znw
aNs4fWvl75+jo7Ow8sJt8PkiWfRGIV6j6nJWryP0Cat7Lg5AKrcGoHcTFJi/dSTN687Pfb9AxPPs
zU66vknc/ZxQs2TnWVHi3sTBlijuNAPF+4puHUaidxNg1DfFv5SBd06T8/Guoka2HwBs1wqJCWo2
q+/5C8888DqYzqHz3JILjoJzSguPUwmwGv+qrUyCjKrRPPRv/oWL3pfiItLwuJn+exO4XnERhp0P
XbTAkDJeDP7nlFvclKbNpkOw3rejsk8r9tkY2YdFoiHm2WBAzZkz9x+BKNRtlIpS8iAJtf3HrsUX
T4ofXjQMh43rG11ZNIHgvk1Z26SwbBzLiNNEfOt/dB3dBKmqmVZkbktJVxk1tKfJM+B8pmQ65o3w
lltSsGm10/vuUDT078NGyTxcTdZVS/eGbKvXjsnZQXn2iWvuN8jSm7MRAXxNwv6glQP/LbnLWur/
U+80ZTuepy624992Burx0xwxvHptTh4IlZJXxZVzoHY4k9TxuuMIBxRt+aCl0V1bXoJHeDWpVBrK
rvGFf7KZ4p/Sw/xAqBSaxyOYFrub9+YgPjWSy10A2I1EMmABYxLsTlsPUkhA69XYWpJdoVQg1Tvb
XL0gaUf2/JTyBaSRAhcls2q7MC7QlejKwDEodlKaCN3RAmANx05qBhMYPOEnO2Irf5gw6tQ737sv
Wm/s8FDOPm0jeGtECnc1M8wLpK3UD+jV6geeRUp8IDyw94ZqIyo+19S14eLhwJlS7PdI9kGC+3Gq
FXTbAF5vWYfWS08002OFtDJQKkJS0Lm/mIUDn6Sgldbntc+HU1K3Y4phqnvZVTqvgLRnX8HfEspQ
Df19EV8kOGU1o+g+RLp+gNhN2ydCtwkSYPSFkz3uPSjozQxahwHLFu+6KIYJGTVXco2OGCbA0ysf
skzS/T/nXlp9FZCOXBv9T696uueZhCwHuuY8T8CW2m/Xtn5OrRoDIXti8mH+5pUGFZsKfHdRB6Ed
cxeXkhLLyg/qKm71OO16oaU7GKZix/e2TmvFkxkapWKyRJE8jiXbik7rTSfOafZXbLyuA3Y9HISy
DhL9eWYEMtOwFktZ9xMX6MlCefUsTrZ8FzVN8OtysoXg7hvkTfJAEPfMqOCk6pfjW0G9FHilHRE8
cjevYcoL0Xv6e/vsubOfp7b1JbLebWtfMthO4L17tInsQs3LGmcA10jCHKkuqWeOqcpb00/5vfb1
s9F6bTXvVUL5DatUQD0rsE4XWNGCyroj61/U6liJlmnEqGGkYPyZVusynZiH4S6HfQqIm3w7lG7S
Mc89WK/qHPv7vruC2RiWqnbWYJTbgkwngZdrt3g2USJgwrj9wSf1bfDsmEdYyCU4TUczmpbdhRQt
GwR36djAs2rzeHiwSBUe7jVTfTXU+BQxsuoQwOCzbwD5z6v/WZXO6ZyC1nrQTjapOrPfc2WY0thC
EpIxHA1GE6ZJU7YfZXpw6vRVysSHV/yLUvzGwfFviBSLWOxeo+U3747abqGryDy0njVFuCkTupZB
KHYw/X0jMPTuv76RlBH/MUPQJDiR9EjvNQjl3XxilB//yOmbeHqI8bzIRMqW3zYLjB2LVkiHjBUZ
xl2EUl416beMY8TWBkhxELB62erd4PdZvP7UkT+X0I82QWcXrNMQXuklnF15tDIZqe9cJMILyqEP
3DgnIfqgH16HSsD+2zPJKAgjFDuwb67cePjhQpq2AB//yu5NiDZm3IMSpza9jSZzOS4RpbhVt9in
p2UQDclT/t2bNxzQ0Hj3InPswGXBf7l4ZhJcITzi32ov2C7Dzudit0jbLbMrGHj1zfKgPZ7dWTtw
M4PC+OKRZLXe9a1yZZJ1HtRF8sf4Kd+1WFw0Yd5cKzwOcO0y1xeU3rKhaJbBjNC3Eh7KVANqbgTB
0YXFgEzMHDfQwfsbm07TXi2wSYrlyCyc31/5vzZvLbMMpkQDlTjqoQbzPN9Kuvb64FvOsgqyU5Ou
gigueOkIWICrwFySDbZJ6tL942/HUsYzky12qaeL2pJUgwQRaxEWse8gh4+/VKG9VKgETlXCP0Fk
3l2bO0Bx3u8jfEd+kaCJ1QqzLV7ZDiK9c6FJpR+Rm6tuXKLdHVCw7DQgyIC2/WAfUn1i18SWsWcx
gE9+yDarl75g3PkQMR1/YPBvA5j1raMJCEh+r6ZC5B2URlMTQKF2bsJJRE+fOLGGuinfmrGU8vRj
is6sWOG130FXdJgVWo/GdImZMoRP+BvvKCwW9df63s3zoX3zzhUaR6D8nndKNwEp+hdu6SkqX65u
Maft4TmcDemDTpnUjPX0+bN1XuHZnpCvy2LxV9yOBgNI5iTrtL+bwiMcaoEofMREtDWJFThzbC93
YezkJoSC2EW5cZH7kp47uEdUaSXxx6OM22pty9bnN9TVMM+jDauYS9lvrk0n6VdBHMCKUn4lHvSU
mk4PaJXQawosUT1biXjDIBBvnUcVFIgHcVuJyqdT6cKZdvRoUfQALGYsWQDeywohSIIbX4EqaOU0
xhq5/SL29n640ycqTWf3zXW5qwAnHTJi9J/lGoBK/3QgH67n4l9/3iSeDP80/LhmHt4SG24Sangb
j2KtTaJr+Qttcbcft7g2Gp3DZCb2WK0BdDd7JyLYCrdrX9QCXWFc4AwVr4QQr3mwURfstNW0tqJV
KWxKTVKQiRDOt3O/ATpbbvnNPWKp2K/C6/uOufrIikUbr8B71RVYWDZXKMsHgWC8Qy5wqfMMO6HX
83VH8faz23aTGS1v+MGV3NT2GxeScZZflhLompo82AJokQfBIn92n2dNA86yO4AHCWupUyC/emi6
zRn/Cs8DcC5oy2TNH1JPeOXqbf3wo1fOEn+0r8GarBhF+gUhGej0VTRkb0rNfbdW0ioCLFbtHrE0
aW7L1SmKjACDwRWgaq/zfHFJyZmqkk4JTkZ/JCOCwRR24OWBgFv/BzlSVd2PmejiGl2Zre+Ys2V3
93wB5ZTtHYifgjnZnMRE9vmDoZyh3iKycLlOnHwNPsssl9F+5TlyIBtCfic573lMdlxtMm6X+gOu
kbWHV9L2t73r71oaFiWAMrEEMETDowo9vUXZJXchbZfl2YKPAIVqTgMytD5LCq8Shsm/nKf4X6j+
bTFPrqH/718DkT6RV2VVw+9ilZ/Rwm63rqSeFe6ibNB+FwXrhODEOy2ecRt0dymm5NCwF7yPQjIb
2z/GSN28ZjHfSFXD/PCuuVzrInGvFoCJsd+aoaTRQ31BlbZtmPl4Yg5HOrbzdmqItrmT3/rfqAMB
7/wKKY0m+pnbYwuF3yUKPfkGfWjwZLDWBXstqYp0ZV81E05pbvSj6vyfjtKPnDHboGVRsZQbv6Xv
RFlaGLARMmA2Lc3Q+L/ZFj3LNEZm8TBhCf11dfHM7I/Q+VUGYw4rKwxH6LzbmRB/pi+HVQh0cBl5
UTHU1zAeg2dDT7gMQmKNul68Y4W336KOjEhynp/16LjWlb522tpdcrLHsN+5fXzaWuJCmntNVBQG
VW88Q0zyFhjj0VKLZYosW5CWKPERSIMAMxc5YczmZJuzDb5+yWPgxQNd54/gQPB7g2dDOGrIggtb
OfFsznNY5OfkngXkiGUGfLeQRBjNXWOnJyq8ECFY7j3N57KUq9tPdKFtFWOCNN38CrdLzif9evDZ
UUIIOgUxjF8YRdGLQ0ptvoQhFIMAkw5GVvVP/8fTkkBBWIEzvM9Hc06b1tLUruuXleKAxQPMOd8F
MXFN7gEHjpl1yk5OV3/9UBWdBFqhEWj7gUrbxcmnr88OzNsgiGXxfR7MQeIYhoACjSqv9dyGtjvC
o2BO5LcsoUwdJsL1DR69Ot9gGq0zP3u8/pTt9wms7IDIh3m7k5yOeazhUsdMGjXLtCl1IOayqtLh
vqr4FJbSvHw+GJtV4xXOLZ37pEWnwcYF34IvRIBupy30Y6PUWTbrpY/IxsbruJHUtPA9cI4BsUJK
XIocYQb1f5jnOySY12LCDddgAVWIzcNrx5ce3cPBkLy5puattI0PqRgk159Cu9Q9JZSa3GAOmIYs
68mHNbqncNi+iQErOmdmAbKxp2E2znWdpm0PRGYYosF0ESPNsdTR+sPCkdv2fbsrRcq1HUhp2hZY
++k4uaUgPa0ggtUXZeLvEDsnw0scXI/dlEQWB2imJtR0dugSXw6NUeCrx/BjwJXf/ahEVNk+q9Sl
qwxeQIH1X3Vg6GjxR5aHlxbEoGQXWAj8wfn4UpAyF1oURsapc5QBqtswnKA5m4v7SkDKF5ugsm56
CN3dLTllQkPTO4VVx2d67wstO7uGZayqMpRDxEylD3/tpQx+PmXsLj2sVFRVbNUqXWZEacF7am06
E1fkUMEWQUNAqMNxdOgKpP+/sJ61Wi7ER9ER9QnWiqiowNMhqmPnJw5Alx30t+YpOwQuFIU4rT81
Qbjs3jeMxKiUDcqKjqrPZqrn/Fl9VrOHEorY5nZsheNguFbiM1tQmH3KQz8Q5XnqMQ+czC71UVKm
2MgO551WhXpEtJKzdvB9CCr2xiWThHuNMfyOwz7jDceQm/WPd2IFdrq53sqzFvCmvXNl90R2JZPN
gjO8e8HKGLUNEO4fUTQ5IG4znT1Hthg41Vw45Fvd7rte7B1crzhKlrHexPFOjN7rQeOQopR6HjKd
LjeYxUDs4aYe5AHIMAF0VZaC9eFjK+UL6TPqw26OR2gKHxIuZkxLnuxhKESWhXHv9HnTE3PygSGl
VsczHHmB31qJnW1bPTIYGYaUv9dkj+iJ+UXfUBRRrylXbBgOfinovYeaHFu5j8riByjj1PC2FmgI
3Ko6lF94NqSKI/QQWAPI111/cy0JNMHmknt/BrMSy42D9/9+JqtkVhDqzf5pLi4np0L8e7irmJWr
D+romG/xSqQtzDq9A1NgJgM+RhU1G8yQgeK2s/n3DXApgGlIAlooRcCh4Co1QmZU12cSRAqorsox
FLnKZmrVeZdtBxqZfuvzo1F16Q1mPrrtLyjy6ZW/DYljCQDBLRUBz4dgiSpQpxAfyCgJFNYiLV0K
L79IiEQY+6CuBOZxfcOTNzgjo6Fx4xaDxWSIcVkL6j7dxHuiLQOyrJgJzl+4soBzPvCRnhSw3lL3
jfaTuWMmoFe3rNYHFoek5uOcwSiwzBqhWY3zluuCXKNXjFmqoww9v36VgvUk/udVOjcP7tXIi2VU
Y+SuX+EAl/+OV0spjrH4CWrlGVT7sm2co93j7sfotpQop5Us62xWbfINyiK/Wc5g29/6qOGvq3Xb
QB+v110vyLzekDambbsotL0ytb7fpg4L1FkKhwKL9qE8RumumokOIhP/wop+W8eIvUG6FYgumJiT
Qa5JG2L3+GRo7WOUDw8j4PkZFbEUCCD/VqhoVWA53vvm2lSPl39i+yy1PC70eCJ7V1HYAOJ2nDrE
Z3zIpDtyHJSAqDeyrkpsMAYHznj4Zv9CDFhDgjNxti6knWQ+CY9e9M3+WFNYl95T7Kh6ilGXbwxW
vYb4tJQzx8Q3JcXBIAz4m3uI/EwHfHnYZy/tZbHq+IO4+ARBE51w/TGS+vSNisbeWshp/7Wo7YUU
10eVmVCgWe2VNF/P7SZszs3XakdzRzSQbEt1JL/9sQ5t7QG/S5No6dxjF5w4622lfDOEoOcuzfMV
3zgzAbGqpUamz4JsY5TnNzvssS/4mJ4pgmkAMYC0kHqUH5VFjjuVGai2CHR+6zja+xLG9zydYKo/
Fn6DLetIR3Du33TwG3AwkOisx9EKFnteN5NNBI+jNLeDem4z7k7pFKbnvZZKpgXcxcER/HsluC2l
jZJsGyt2yYQC3GucGPNVuozEL3whL8his0QELKxzeP4EDgUF9lU0GMWncJnZ+BOLwa4t5EKlgl4N
ivhFZRfaFRvZ7GIOUY8yWZ75x9TvebEJvbAnZ3wtBHNvMQMhDifIjSO15/nC3hjf+XSUthDFEFXk
uFbMBEu+zGKK+kRoKumP9JlwS3mCy6FZjgkO/bBCg/Fc/2ywQZKVPZrHSIZiCWsjdRLyYAv7SUhz
AqaysKhPAjL1mZpYK4r4HjHXYif1h+z8/6cUa2+IpUGCdmqgVhorXDOBE7JgffUx1b2LWQgpdfdi
QKEZIk1LPHw3DUQoTEH+kiwwSj2w+kqywtHTKwuGLJALsHelwxUQSde2gyisyIiP312+xn+nZyAj
8/4+EiS5YwQF8ZyjzeR1OwrcfCxjOCcjp3Xm3hxQNihyU7+XdUfrHnCKzvWRb2O4o0CSfRgLM1Vf
q0+X08BHNpbIC6se+aVXGHggxUElCClQmxmWNAURAMpuGqRzal68rXqsQkbn4m31+i57L0DalIXq
41Ts6CL6IPSLjFGyZQ9eoAgTqJSzJupG/Z2y3e9RA10QuuIazjzC9kF4tESfqwPFCkUvZMTgwfh/
IGwVllZbgUTsIIrQki/rgld+g1ZhMEssdz6wkFpVecrEHroifmnB9dHr4PvHMIHfZw6ZsiyCS8YR
muBzlj/oWNiaqaGJRCYY/sNLuUAqzUH2oKSgt6uEA0BN22UP1ym3XyChAg/2nN0irGkTYOXu048G
6vSLqRql3R0WqlldMdZPbKUkQbmQ7jfi6WcHS1CwrbsedwlUh/3XoAiRWL5ZOmOm5tlOeBsxRQz6
aLoviAgVUvrCIaIgoxJLMI1ib5ZkACZ5x33or0ODy4YKgj3Gg0It2sQP6wJI8eMHUFdpJ5tpg3VG
JYRDN02/upmFhonv07yG7WfYo0s7/9TKh1B6xRiu1n0KF2QEjXmUhsQz6lFJzNTNgxJGVkt1vV/H
SqnHY9sqAz2QELc3VbA++Y8kh69shv1OZC23Vku2EATeAqT6tImlZkD5I+QsTFe1GkXeGP1DCOr/
dyVnzdMk2qr6PYmZXM441botN7YTRyTc6Q10c36wjlN2lfWSzeXZ17uQktUqJ0FIMH20WxaGb4gR
7rj62z5zc+BLuQyz+ZvLPJH4zvKRp+fUk7HAYY1SoNtTOohibDu9or53bw4aL4lmf7WqX+Hn7kIB
aDfyFxzFYYfXlGoK9qTBEnpGQlj1utC0UynIuxrQCm+DAhmK08cI9C22WRbP2ZuqeLXR+uVONDhA
5ub7vqa2uXLyQ5EeoQcKsDROb5Pxrh5EE46PbZsfscEPdJIpiTwIGL9iL1RxYjMouP+9qRXFiq6s
2PnbQrPyP69OM1j7sQKdR8iVMoHA0oyh+IwIHk3/NvFhICRm3yXKoBoAs1/ZUWUP4iiMp5xVpHrN
bbxLlD3PRqGljmKqPAEcRASnazy7tJEnLqPJH/wZTGBnim/mUKh/DH3hngU89ebFDehO+6f31nA0
GjIblrOa/NMIPY/hgLfirFeyEY/9fv0NDjPRahSrnG8ZSVuZiBtximnU6CIJv3T4RklS3zeeNuv8
FFM/T/pyY0Rcu5WwBThZCMdV3zyiYck1oAK2fGwxKJGXeycb386REwJm15GEjce4VXJZVmi8LFnr
oK8bPy0kGcz0bSourIaHcNjCT5NDifcSFEnPRZ1qTsp1vq/MKQiHq9Ulk/YvJE0SOW+TfeB6+mCo
z1qrDVPzOsWJcCiGNKWsPbR3gopem5Br9Wh35sE65/QMGVvuwa/e2HPZ/B5KfhQelTieJrS2m8pC
2yWGeydtuUTB0xkYgUOYWsoq3PdMXXnUG4auNUFcYi8h9m+bl+7nSc1bhVw83paOc2G9d6rdVAZk
RL1R220DbUo+gTEYHjND/dqUVHrpYqFUcFRfTbHmFqta9LNyCE0Tejn2PsapYEtPJoNmC9tR1twq
nMUicMXPkc9kBdHO5J85sRS1UbSk3NcifwfQz1IZ9FiPQCEOw6IRNVE60pIl1CVJj+ZeHGTYSbKv
Ozu9phBIbxk8oBBWr5Rv42cgZ6C8IQmnSN8lAIGRVJu5bYT9B9ua5bo8sPSTxYrtdxCd3adDVxRW
K+y82RoY7b6pnZhx2TNA2Oy5J91PkNZLQAmsSdGzNGW93sVe1doNjA0Ic6KM552J1bxKK9hvjLjA
IjgfTbO2B7Id4KBPJKtwsZcOMZtA1+kRxoRRl6IUideufihjO2SyF7xPzlpUkYSDcPevC008rICO
glGx5KBlGs74JXE01QuEA4VHRWIDZ1Eauvd14rFyJ3C+Z+gCqHlvgC4LgzqX80c/Q95n+/txhTCZ
4mE4FOXP3AuQk2O9kBzd8t18CslEqseGUXM6K13X1bJmlf514OCFhzG2klFYw49JoEigSaA1WtUl
Xpo4zEwwto08ebI2OwF0eF/yfaqvIgSIDfIKctqLcBGFcTMgRWbdT+2l+sM/4SRrgl7wYnR0uKF7
Mgvw9hIUtQoZrl8FHwlniyKXPxy4FJ4O3Gbr+Bc7ys2pvSFWBOFMv0MdbPb8TBwvzgM2Cf6b2bEi
opyViksr352e8RSncLMmyl55pGwATQA2FBDecjH4Mp3gGYFkx3pB1nTJaTpJunuS4oAjVmkHQjnt
lS/ZVHwgz0Ayp7IY70R+0S6S7NrTsKDdbOKS/Hd1voVmRWAUs8DwLIRmExwITmbmBR7Z0xTVR+UR
I2ETrJ+trh4pyp21YY+RBuwc9QdwFjC0ne8SPjOLjemCOfO8EGwExJ2A7YbiRPh5Ckn2V1ZLgGu6
HmeI3Gr5mVRM9xuiyKJIcMaLTLT8ON4UX0XTCvcpCmLSJPOLdIzyriNMpd0UcGzx4Vulp+LCvYoo
JYnir98Sa8dCXoPOkTfbqWUmZ9bch8pMchoh2ijqDEjnm/1r7laplzcfbM2wH9l+yB0jG1Y3vMJH
I18yO3k+ZtmkZ/Kz8iFc4BbcMG9pIBQkyWnT3yeodjVVEKrsgpvbssrkQTgYlwqJuiLAtXWf2ek9
CW5tm+EV+bH1tTZNOavQ08XViDWexMGYiYpy1Wdij2LoMML7xqZ6cju+hFTmfmAtq6j5demhZ1rj
Ncf286Tql1krs4DTz556OVN/84Z2iNvRPy/GKbDWez90cBVUiL4ficMA7510CKpf28bM4vhetr+7
F+G+g5cTa0+Z6Q9BQlnjzL7V7oQpbIwf5HUqJINHKXuqWlmKSFuvzIghpntyaEDSuZNNTti0f1pr
6oUuRVzlP2+ZaLbSSQ7dOUQ08JVLXok5SZVdtC6eNaqlgi+haf5Eq9bSmxzpHi2tP9axpNaU0kxo
miJZgd3HkmjaLoMz1WO1ppO0sZR+0YwN2u72ZY+0UmQmSD19015rKAi3fx0JAKahuF1Z1PQdtZ0X
pFo8Pg2uN6dzdFSqFxo08wcRydpyIMfwpY5XdbyWT7BUBkWdcYlf44v3FXnnxJPn3eP3uOmbdcWU
TGX8037GGtJQNWOf34Kkidkf1PftX6uI6+3hOlCj6fHb7AyayzoEeH4h11H917iA/xU+qSMHisei
krixZmkLK6a/CxadQaWcMzmijYcD9LxUZZgrnk/E6G/naAvKtN6J1n05q5RBaLVV/faXv3FfnQS9
ju7A+9s66N/2jWl7wBhEd7bUlCGu1K/NV4Cc3T6Dm3Oep8JVYmQZR5v9awV9KpyPRD1trN/7XBua
QsdYbvBuL8saH20mu3BjkvB0jWzvbYxr6JFrzhdfl0CUmzIX6/98fsxPHbgbokBEoQ7RtX1RGwr5
8A8CV9czf6kMvLGnlrV3UnxmFJVKvXsPO0hBFgfd8k53cVq/Pz1B8Ivxc9Qcegpat8awYyNWbXh6
i+Ts5/ialo9yiq86XTac9udVq48Dzb/tAJfslKwWP0P/XVM60vw4jJROGg7vLKmKTmV0nsu+/0HD
vytlR3krr1nphuWuqKIRYQGBXGq24Y70md4TZh+qlU2MvNIF+vbhsWGsDOj19dtnkb1I6eas/gp5
VjeYwPFpasCqBrdjt2MPNtwIXV+v5JmpdPsvMlJKn7wZlGdRkIy8K+ZfNlf7Pl6GchBtu0L0ngZ7
8FfccdqKqSd1vbIGnzIMKSKIal8kYZzJ1In+11ooEWfGFIx75fJAU8h3csUhr2l74C1DbitrH7si
ztUiZkUKVHMSC/U1CRZGAHhwA806H87qeO6d42khQJBJMbwcYLS42Dvdbl+HoR5WKW6KNozEQnM+
s78BixC5v0Pp6pJhA+DfqtRItyAkzYfDnOgdFFeRSxIX8/oJx3T7cmX27gF5VWsnUnOkQHQKSswO
P325fRwrMmZ36QrNhagyW9A5rOZyRkzfoSg/SlR55OuhlW3hsUcze6SWWPitOINMwQqkX03xHHMa
9cJGLZmA16zeZMIrqqusMEhQSnRsKiT5irduArQrimYwwmjFgD8WEbbfUgR/gu8kFzRuNEF8MALQ
qYNVa3DomRvlSoxPEqyo0f3SOrdiWwjSlHFHNEe9XIovZ8ItaMUxvoXREL12h69J1W6nrpP5DvYE
8gFwyEfUIA3GRyhxIMbxGXSuGvHgQGyjE9POtrzlKK84KTHNUzgYG+8tzQ4s2x7bhGF+W98SAvmM
pK/3Ubw5yTkxrrw1zAme/Y4GkfW71EmzIHtILpMGkZDm/BzjYo7hvqVXGz6WfepVShLnNvIA1kjs
u2rx9lWSettWwcje/Es4TlPEC6Kxy6UbHCxPNIgQSIQ+OOHiyzOqrjwdgmwZry6hluRgbPlQ3Mpl
RF0Qx7vB1jQEjfWTuF0AqNRnVkGS76zR3RKn1dW4n1Xjgeh0umzq7pWCJ1JYlD1X2UlEyvXOxacp
qI34x544nPf/m9F20y0OTmmxtBYoQOK6kQvZUELuXtE/xidwoBVrKC0hFgA90OOCZUDn+ZtwWf85
hjeRt8u971e4jaZIboUPRktu0u2rQd8mDntmGWSFdhPu/fMqoszg2ii9gFiYehk8IRqbtZVxGx9g
mRRLAU6Caeacznmz5Z7hlnRzbvh3IavqEq1DFc7z4Ath7VBKC+aLtHbZRbwRzDWnPyVYAJ7jRZKx
zXIz9e0Z/thJkbS4M6j2Q+kRqyccVMgiHIJazJyvp1aDAuBjxEUJup7AZPop9dIJGjwhFAr+6n4e
S4Y5uRdQYSN9Hp/4Z4J6LrxXJyOm60+sao3KJAkD2Y/JxEKEehKmzJdh1C4S/xkTS8Z6xPl3Bsoq
33tDgD9Vgh02/u0UQSCJv8nwBj8SW8XhChrV2PtmuEsC3O70Sh9stU1ymxELD+ij443Ek/rxV0MO
i8uU5UoGmDfyHULQdWHaB+yEbhFjwPphf9vM0rHWcC7+qHDOM8GOdVZ9p4SVRLczjKLSecoFjDMt
r4QwHJb0/pz0pAJyF6iGtKCAbv5cej12qa2pN4jA8FS0Zt9WcXJByVwlH0UdBlQad5MJ8KflZJV+
4d/tOj7XPwc9mZgn58weVaokn1IEU+dMwUt7MWJhUmst7Ane028h73FgEYyl89gKkykrJNaHe0NW
wD8UtFiQtcSE/sWoWIXLfROwizBUeUzlbpNQkM5xDK7uMznjwXYPQOyhCGP2osrpFmCzAmrBgUBX
AF7zjIB9aYkPDE/7O47p7TGzfiY0uJMDvzl3C8X2/6VNyA3Zdvbv1RYmFuRM/rdugyQimkczAovI
s724ixyZirX86z3LPxeb5FYi0yv2cRmpcRp3GN0aVCBmMBA85Qrgh0H/s4dG2VtBfwFJAZfT2aQE
PQ7iCZWmtYRj0VUdVAP5hiAgwyfcAlS9MzFzUQ9IOWklaXoqVylAYCc+w4rdx6unvvMQq1occh5N
A28IzqKKlGNbhnTdC3znjROgWJ9LMqCQiDkQ7H+aMlu3DhCO18ob2c4jwTKXC6XmZg2E3f7BJ+hN
5Fs/ztNxp+DBVqCirH9Vh0Of3YBIH8TQouI+1PdWDOlZVaKLjyfGouL1l89yBXASf0LxGq3wDz4a
M96PbmquJxIT08kfyLcnphc7+AqXn03wPEMYnmouAT62sMpKCsODpvpo0mV66oNOEe05SSE2ZqBP
QfUK1sCHbjL3jUCKRHyAWm2Ti7A4HllBB8nX7AgnL1jTEzWNiBO1wPMD7MUnl1B2ayu/ulLNhIDH
4i2EuepX/tvO+paNlZ/sFRB3gLTuslQS/avwx7eZ5mHEnOxmfQ9mXJ29C8x3CWI2tDmH5LlV9Flv
8t6p1LuB+epKNg+XUNyz0VmOTvt7ihd0jkm0ST/FsqirXBa6fkcZyVh6LjZzn7xltqIKcpSjkci7
/aO4IaTGNSbmf820nS4uprdGCG/8nHjeQJ3yEaW7/zYT6DpEJeJsgAsyN4aCgI047szQNaAlELwk
LUJKAL9WeK8POLdA9pG8QU5dmbWFPBMEb6D2DU4zs8tYdFufA/0HuJFrrleHC+65y69GcZWmgJiE
DRlO0B5iL4gxoNI6Ppp8MIoHdUC53BCR0+EyozgQiNYMitcIRUUGVoTYtcwy/vuqIqbtz9NTTQEA
XppbXydxp4IoVbdYGtoDbLhxqYY8dAwMEhM3Y2lPtZ003vP5+EvfOhN6Umn4rYUTT4ksctTOlwID
3bhTgqlN8e4rgA2bGFWfECgsDv3L9AfLZeypx/lPMUdY6hyVjbg7esVtl1liODfyXCOyvKRXpPMH
SmmJGKpsfs7gGkj41xxMQzlCs9Z0onxK9juOH+qZ5qo6zn1qf1E1G7ycUkjoa5DLt0VYKqYuji02
dVElvmDZGY+wKInTgGvVjdnu5KPki7AUqRBsC4JC/NuRfIT6yzoRR99Ex/VkQbWl9/4HZgN4g5cq
v8YOx6KD3dE40SzU6aCgqRB/DYqH5oFA3B0dmI+vT/z50aDiFOMiNHpVLcoM0A5cuP742Jv5cyHk
FvLuZT7zpvsU/kYiCgMXFUePG2DLxIS+AfXlqUf8APeNF23SbhKMm7dM4cfQOKyqIS51FTuW/l/S
3FRrHsF0fcSIWq9uUj6SvPPKuLHmTCEd7JTv3Hxf41aRIHnERfCdls/fkdYe3duu8dAqPPv94YDT
X9fgRFuqWlrcr8sb9CtpMiRc4fKt1JkavqR5LuuTT8Acgr09vVC5JNNkqi8tC13HZY90Kapd3uv7
K0aANSovfL1T+HXpMrxiibhiiT8BtwNgfkGI7oP6ifVb6BJVXvszNAHf5PvubJejjCgN8oSJaf++
aTntaUT7BcODaXM568xXA+8RIPagIIcYE7Nb2T+jomztOgAx6gZDEEORKVUdb865sMxzImw/gPor
lPTAePhfi0FeT9G+GuVgsrdssTPSpvQ0up3+pYJTXkwOeOSMNBrXwPLqzN7ZErHsqMwsPqcZlriX
vAMSFj0Djtv/beEEZ3Ii4mxLL1uVjjP3PFNK1GaJQBeApvxUvzUdm35D4tiTF9isED47uUbAP7xd
MEc887ysvecf85AkWmmSLxvtogqi6VlK5RDoDuAMsULxwFsqQYMhL/QikwXgTknnC15YasHDP721
ikG758A+RUFXFqj9U67IKG1I46d7/HdGS6tAwB4yrj7yomhKUWLHfBz90lE4RiswjCKdPNdKDqO3
M/3ailrnzJ6FOM5hNQlGwYFM1dJg+mQAB/vrRv+ozItjGeedheP0ucWf+dH9Lx2cljIvogg8HBq4
aT8pZTf6KEwjH2iKc6m+kJTP+Vii0ZIU3h5BvSSUirLLXtSqMBTLc+1XvGCl2i6ZgzOHHxtOVoxu
DyqMhbEG0aQISYLreMk/qcBICJiFQfWxM8hXC+Tlqv/Y9id8jt2OeFlZf8LliMHO9GQfqG+dUktV
TL8hsyt5k2F4wjpVLVq9nZMM4ofj78X8cfPgn+rocwWDsDgrB0WTA/jD5wFdNHx5va2n/Jw8iAfm
zbK/Tb4hOH3Wmti1ZJGr/gxrsgt391hdqg8jjkDOKxbGIq5qS7MYsQAI3yhQxhegRZCo9IbvQtuU
moQEVb1z8EbegcyaRR3REir9acyqjvA/zR/d/ifQDXPXBSSenMyh2jI9zkaCkBv9TRPLM+YaVXQD
/W07WjpuC4rvkVAFdTpXrXRBJ0lbTtRch6l8we6ODoGtpcvll+5sK9/txJXW7Jyq8ttRzNRwpksR
QANyoYlxFCmA1itenFjI6mmtXpI1JNhyQpJ05bvNmJG/mdZxf2giOm/7KxM04fyS5m7ejy5HnijI
m/iA0wNd+hTm3R8gYsLttlpYAMuMtSIcrscyHyTi1gnm+PdjGt4ewXb4NvVs6FRN9D1fQQjR+WC3
eO6U9GZDGF6421gKBfC6yD32n/YxQQsustvJkrJqDsuVtXxqbrdBAcpCq++3Abvw9zHwfKjXL2Nl
GQAY0cF4mcb8oUwZy918NeU0Eej6r7ET5gk3jJ8MSrGA/HqjX8WpPf4AayrOKmYNY8VQosPhIb64
g2ChkIt08PSNNz5KHeINt9poSwY51R5sXuyUeKhpJLKaISH86tkBjhi9gWBWQD+ylxPnJGOmEIzf
3bC+X5JkBUwocPWBkU8a+bNYo+zuEPulgp7UQChWy3iBbb7ybmRyulfuDYbZ9WWjNJcjn7+sYSC1
ObfUcvWpk/FpFk7VqvTapay/8ygSyWJiMIp2r02/NfOK8aK+ysM4J8JLH5aG+CC4mzc00IdFKEqb
yYZrPu6YwRJ34pSK9O+QtkXlE6Afn+M9sPwAkeTIaPxN4ICdWqdktD3EPg+OW9CRQtn3OKVgDOOP
HKZnObH8aVTLmknRxiR/Ozc6uAeUc21m79LpYNdyF+ZygTjw56jzMGdmLf/kwEQ4yj0tVJTxXHFv
uSK2IsgMC3c2uY5y7Ieq9FXmrOcQvDmOOLHsHf/jyQ9IOAnyNCY6/ARgR5FtRBMxiDPmrPlgWuTO
s6gqgvCH5lsJrnDlvnwXKVhpoa1NLo7KMmuB7urewMLrhRNTP3ygQ62aSfhFqYk2OSKiDARYxfAs
tOy/rJv0e6dEHQQt7vFFWXHeeY/5hPqyPknmLxQ1LCZ3+XpqTjjWw15C0eOgsHUaS6G1yz3F/YRt
/otQ5vgATHubb9AzAXfCxcgdQuB1MjTw1a8IEwdsJk49Lczr07zQGWfWLM79ZpWjW3phg6ERepgh
MF0VW695XrHZaSVhhkSilrL52wd9fgVel9kRtVOXwMjujyp58PQK6U7m2E1fmwMPCB8zHl24QEkG
b3Q0c3d9QOfPCJYpUK8rZCBj7iLG6sFaxg6m/gU2OD76xLgFU2RyOObzMPGZBLGu+MLbR2keUpOF
eu7wokhJnl0A7Xf6dTCpOjPNIbJAQubz4fECYIouU/xXZ73nFFnyDyy4RfJ+jrl4idef0cKDJMop
hxTkoUNf3GpyrJQtjEfrs7RAnskZD3RKngvIlvaC3W+Xl3bPkxCSVRLKzXWYc/uuvi0PcHQqXV3s
5ajDPQGVPvjTkJjNK6XKLpBua/1yNvLBjmdoBRzJRUGjT4oThIWKP2J/AHzwBR9JhFCkPzRByF2Q
3oA1LWDLHjYYrOnOvmVOsYogNwmSmj/bOdQeZ3hSFVQI9AlcmqznWj2BT9c0/hHL90jsx++U69W4
womLftPwpUCQeCC7W8QcV+VEiOyyUVJcZVBKHoGE1zzRImanRQ18CVxVU6/SDWwj0i8RRc1r3+jT
UhB5HuS0utzK0OBqUseUfbZoWJ1NyD4vzk8Eczpo7pxOEbg7+0oqHYPCoSsBymQQY1jNHIi0xcr/
3Uh6xgAqP/pd8NeQ8jf3+VkjexRAZKTwb+WpHzSFmtk3sQal790RwkxzccV3JPGlIY64iSRoVvnn
AObMsR3ifXgyp8AQWCikpHBR2wGzq7vNL17SRE/VlfdUD4ViC3uehh6fouVjQGHfwVUN+hWWW2tW
q1QHTHZUiVgjnriMpFqEuTUaY5yYobQyaUymX6Q5LKlfsvTtGUiXdlN0yJgwB0x33Xv92PHXh0Qe
TlB0EwGsMH8F7D+Ukor2RzlcXqOsgY0HJ2CJKKIHZWKcqIJzSm5dYQa/2EHrKH7hWBZOqmmOmGg1
nMriGdIDquBeEa3IJO+haLhA7BkgI3P146KClpcdG+c1gggEF+RwRY3pyqctKLt3BTm5yXwj4AW1
y4aXMxj4T4B0aJ2UKLC3FG8X8b+JYBb0sVsO+D7TU57XgcLQnWSCtTc7tNdZ2chWIypASYuPuD7F
4yl3DgwYzY/JjC7tQEeWPZFiberq18qpoecNWQ3mggHW09rrFyz838Q8cykzJ0NxSaF2vvyoBaO2
sxsBdicpkOYk51rlCQY83uG6V5mHiufHUYHkvfj32YNsET4RoTETAz5Dt31+5pVvPLWk3ORT8VHv
easHHO86FqmYvJVErkqXhuQRep+c04Duxaky0jhVy3L/AlbsgoGNHcCzlUe0j6VWt3iCyfiTSQXV
0s6CnpAl8qupgedkA3NBKhBiG0eTLoERHVowGBMQQhCvIoRzKzf1ay00Nww+qIVjpLP3wFVhor3r
ljOSklEHi/BSgz8VI4yf04nRAKsz3OIY3m4Jmwy8fxN+IxziwUqE2JYg92/hqZqd7VBOaLK42lUd
pewsxXgn2fLOOpQzydWRwc0qjZHmtNfU3haJovYxAZTOZXCew2CndB7cUFfMsLci79/o9UBQPB5O
8or+fskYr+LzWYYvH30LQrMNn6hghTL4Oz/PI8Vvazv1Ktgj/kAIjkObN2HLLFyk0O8J3glfwJsu
rmQLUjQ8TjtfxWmW8d/M1omRRCLg0CoNAdtMJ52HPkYoOWrTJqY8o1DQaAuXJYzGmkgkUb2Kyylx
0VrPPZe1Km0NMMowLh1MrBbrG4VXQpSe4LrpcyhBCiAWnGZ1+yjTFcsTXtMeMp4zH30uUPn7ZCMs
fCeiRe+EhHGTMXxYw8BdZeSe9Ddvu2Qvh5x58/rypo03yo1m/nEtiqmaQ3ePU4MTkNVSnDrLRBvc
Q+r9lZ0scEdgpMyXS/8QZ1oewJziwbc7zi7OjalufCUSDbr8FA4y3XdkT48YFP/GvxwKGh/gdYi3
873FQokXnBjn+pAbEb1xCKglsG5/fjuDFdYyScWetw97zSuhtkFwe7HfhoWlnbQCAyR/BVR4WfMw
7Xv6JiKFMMuswZkwCtY/QZ0khi4Q7x3N47OfEL6jp7PMePbCqjUnKhTngq4Cn3Cktq1/QU0q56q8
22KvpnJiQKJujsz+Cz47ZC5Tl+BJ4RtXMJW5u+3I7iqLDgMY3xupJP+z9hDTrJpLPzIi/tvkh5k5
7wLiXo8g9Zo7ZyGdPan78On7tWakEldXKeY098oVkH8W4LKJDC6Z/JQtLEVLKV7kxG8uMwnJmpqf
1/jFrvKkN24NLNofDPQhjqnslQC6LogY9qI35pvgBTlq68WII5NzV9O0Vx6W6n5NYrdJDuAAKmyb
EyN13nWrfUCC55dq0c/CfzR5FSrElirZmvrnC1Zl4RWv5tGn6050Z0742rTc6ElfJzM1WK2LoigN
85UnJSX1B+VolfyL4kDbbvat/ImJDCaiLm0gIQuMOV7U260zDD/LcAflod4LoVtEe58U8N8imGXW
n8VHGER8LZoLMMpLppLd73vaaXCG1ONxg4HiXUS/8LlWEIy9fu9n5tMq5isFr4vVvdVMOx3tSp2M
KoFRW7hKrc6fQtBfjB4c72V5q6jgNXmj8pxiMmLo2zHyacO0zU/9ZLSNCg7MT6T4MTCuyt0E805e
xttiz/2ONPo6g+BG+LqfruXS3Z9FDwKj4LAWBxFphgpM9h2f4axEXdR9yeWKcubO47NXVsvt/aY0
/AwMZ5RrUutARAIAsyZBwI+56hPFld3VYK3wjfmdpaSZsUOzYPUKGQ/m91P6EaaxrCLHez1+ea5i
Xp11HUvDcVAijoT6ZCpIoFF6kjBireVYRMVg16zRJkKbiIIyCsrPfaOqZcjOKMrIBuPqJjxazufG
J8OZy0YFU5CkD8EI0oXIR/nRywLY4xBScZyOQ1kZcn3JYhsliFbY5Jr7geiNdVL+SFuKGyrvFRyo
6OZq9VZWmeFhyC10D4MVDGuuPLMd6oWCcpMjFFv9yEGMrtzOOyRE99rQTx6i1ooEHXl8k2SZIFcT
i1QQe+aviTFbpq6ccR5+SBWJ2+GHqfTMrMbNpb6iWzupH2TWu5FvWszI8DqIIPtZNiRABSydaAII
OJNpBZ9O61A8jJjhUoXGUUgBQ2q5hJ2Wto6e9QjnrFHEAFdGCNiyms1DtL7RD2eUHpyfuXLysTBM
UafFjHpglHPfNryMN4O56z5zMrRLWeF+uSE6zFXRd4IZgii4YYtsotLYe7tZTcf2XMVDCU6Cq0Z0
E2Kx54jfFC4oRA1eOkvaqvoxibS9oZSARnSAFa0OnNT5tIDaPB36vVUOySP1N4n8NG9pSMOZUSSU
V/ap1tHcZJrp3aZm6k8p53f/tNy77tf7NVQ+BvJ87KXOx6HJxrRpCQSiz63+W7tpafpfS1JC+SBr
W7g3J9GpTDQjDSEkcu1nZ1rmALUgdCZjiQlV2klq2jOg6Z0f/bcyeIAPYpj/ILuwdpc9i6Gk2IV0
3z5vrmyELgPFyROUDm54gaJqGghXR+PLgDOIfnQq4yKbHf7Rj/zuUb6upPzDTHrQVQfSoyi5yGCB
ViZ9MoMDoGBiQVutPbGLC/Kc5g4G6sq4UBSTTrESyAAuiFZCasLSACSzIRbaoFrcL32eWZCb8KkT
jsaogG0xpYkA+GQb/pM2QNXqA0qFNCwDF+urWwWOf/cfWlqPFrbTERknNMDy7GgSTyg6SDgfmMNG
j1vRQq+MimEkQJJ0niHSCIujuMU0iYRTJ2uoJrtwPJHUu3E4Y8tJE5i3cEe9hwHiHzg5uPm1rD7f
/SiZ+C6msfBY3FEQJYw3hvXwpiH+WPDidNCyX++vkt7RtA24QD3Hyc9lJml3JGjtTShLVblR2R/H
XpactbVTPURcUDxmwYWVSE2DvPvaqgzJvyR+e6z1UoHSoTh3XPJ8TiPqYl7dcadgftnHumdAsnY2
3tRX97CdxZsyeSaZoohletDAo7g/Y/AaSJywuK91bm9AYTiWxNhOPKJoD8H0ijyErcQh6b0Eff/z
nvNhnMjkCQCg5QIKw9n9pBQBIZatdYgAmUKoKexAs9mdzYOPP+19KnjLIdVo7p4rxbAUJc4UpuNP
fxF0oK9yAw8VVaTOFJx4trF8BxYS0qr2H6gnmczRDN+kCEddvPmIQ702F2lrZWbQ3U3mZ2snvrL5
24d/FP0AQ8kbAAlB+VeqtaIf+Y6aCMvhFb3xHJgJWZZohWDfog5n8Km1tr859wbH6HuqhDLYG+3D
tRbYK1CpXbj2CYisHi3z90twmuh6S8zdUzskMJcQ4t8wmm45MRdaH1SNkhbNsZbr/AW00MLZomD9
Ks0R0F8FFE7r6ZiqOY3Tog6xrykTNQdmgywI0hrwCm7x5qn2zU9x5hpITW84xB34X33XN5DjEGOg
sUz/sktMEBvLvKf95Guh3tdiMj4KBqQe1hvAWrkNFYS+D30B7bz6vNrKEhVTElo1VAlXgCzy0Ub0
MjYR6PAcpORoqa34unZCvCL2qDfIdqIjgQWzy36C5PcOf5fndzu8w09yPr6s1QtF8zo/k5c3BNZo
gzb8wwc4FNn9ptIGP2RS6fN6Jqum9TKA4P6fWisCH+u7aFbBWgdvcV2fKCPyG9dfdXo7W2XavX3n
EJ3yuryb292oQ6+6FKvw4X3bvtZJTZBVuzy5gQKzpkcwEizcB4paR+gK1CC0c9XwNIzbaFmO4mb1
bx6x/ihiq1VSx+1VxHyGomq+qmU5A/3T4jXichCa+XLQ2o/uiypmIWNqdqyeF7nX4rsFgqaZVgSt
iE1sHVgW4KyWJHqh599It+jDQeEWZYtUge9nllNRJXzd/gATPNts3GhQLlzJAa3iS3g1WuvMD7oz
HK8yI26VHc9NUfnJX+ox8Pjlh589333Ru80H6munXRMbt2/Kw/1n9QXiLRlrgFGu6ZpnGA+Zehtl
y70cezMg40eYg5VRVPlQUaZNJzMeanSMCkxwnoyHQZa0/SQmqNRVKGcQtoeAd7vDFwFz+LAwCeWK
29GJr4Mbxj+7oF91eT9jD5nStW8CuU4Fv4BYQolrGjgLgA8JNrE41SeTvljfdHlGegoPggMD8d0h
UYUVD4BS1wOArn7v+9B1mpBaCxKKyaW6M2EXa+xVUaYXYdLoViap4vxg9OrXpQA//T4sttx99m2u
vuvEdAO9NKdv7hvNJnhfVR1oPG7ArsvIWZoKi1TtouzAgDudxO9GIK4/067q/du8y8r5LNE1Jsu2
xT7yurxrGFDJP3SxqDDP3jLK3iTpkkYJpGR4VFxWdlixtTBOiaJ33qtnIVyxYgka7FVBw2RHooGL
kTdzctwmaPLIgj/gxanLGo+PUdrl3KyvethsYskuUAJM/vDCL3IlMoCgobSeYIbUWBhM8ioZ876+
oKOUy2NHMUJev3jV92rGxyu27WwcpYXZHfWHSjZFGoyQULtI4S2B+nAonJDApJ2AWaLGG+A7mnBt
/s52poNDs4uWAH5XHsTzL15oIIm40pYBAm0PS60hJIQZRdwFB90vR+VXlaVpxZU5ZRj5U2LF0DZX
6HMggqsCo/AUZGFSDk4681uyCe2jLY+CqYoRh/RJg5PvA6ySlrWFh7Wh387FenRE9rBtwG5bdYdG
1L3st+suz56CZU2r9Hs38EnAsdSy+9wCe5vgVVSJoRnz1K341czshuXRYSsqyI2JyMfWA0tgfL+7
DkSKkOrCnICvMD5uz6ILouyU9L+0kwxQZ582RliYAqTQsJBrKC0RHujHbo/JCkdqJl/RFLVU13iI
J4CIXmhTmUx/vlIC52vpI9pzRxUXxey/bm/v7mr+/hbV8LmIZy/lJFJHBt6zQ/7fbNGVN1/EM31P
avDwM2vboH9lmKUSQ81B91coW/uIx9ST5WjRy0HeC09K7b9QGhTEyP73vFRAbmrlfNYckANSEzWv
TIGt9dgtAiSDMHis/Jeir1OFmChZtJieopDx9ffQHTs8Tl4Xl59dwfgFAlTqKqVmhvuECBjRc/1v
aaOhn2T/EzuKCMoWGTvmfmH16CjsVVaOLNb3T/goBDIE2i4ZYUZczUyf5ZsfxYA3dHM0DvNqo4QH
xTrI8VhembZCPn4N6gLWX9ugvJZBMK6j6YQs1J2JqCV8+/jCOZx8Jo2+12cWd9G5hHOwZqO8/ZQ5
pxQD2BFCu4DcUv8i3JjQRv/HKtrSPDW+eLYcthKCZRR0bfDtNHuMhVegv9vmYENLWT/lY9AJWNb1
P7hmBEANFnr5bNglGhMnP9UWWofJztn5SK5wbAA62ciox3GmOkd5WOWSX6cGy6LkgDQWRVbKDvS1
B0q06eFi7uSCVc/9Wulkbdep1NMUmqswD3Qy/ciF/u0+AQT4sNFfmKFvC1E3UyJLdms3wZJHM6Ds
Pgl5BCjCkU/z2qAqwe1lbMM66y+BXbB5LP/cOz8wX9DwyCfvrCqOZiANA9Wf/uFFU5mTK2BYRPBg
80d1iThPqUkk8AOuGSfM8x18pcWd3OUph8RIWpnXgpzgDxxiah8/Og0oqmBClYG+csMpcsqizt7E
uokPbvHfPF3EbVTuT+Zi1gmpN81s+hlfV34d4t8RMF6r4aW8V5sDHDaOeKjrBd6VdnRgrA+jcGRE
nD2u5lEfJ7KE5kPq1NYENXCujZ8tcvqM+gnS3j+9PjS1lIkL6OyLnDmnQsDGs8xZShKVisf+hGYQ
7AnhVr+HhGPyz0Yi4z9zUcLEdAopgvge8oggsNMTZO4q9CRbrG/EpsnmhxnVasEBO1DU7TycwUMT
TsMN50XMMjlaq8cJMJ+uIIJ4klThUK3SmU7Fe2xmwHBTEEfBqekGVnjpd/bCkLzCIhGSEVZxL9XS
sHbe7MlsGaBjOx+qos/LobmLRoKGDpwZi01LJiBg48wU+B3a+g9vGnXMCeiMDmj9GvZNZQ5YXdku
DtWq8VNJPdnF1wuRfOEwgVZR8ia9YARX281uHcKsdjxH8/c9VLteOhiuHjEsQonJ0TY0GaniU2/X
xLAtW8GSjD81dTDEyD3AVVkAVPl84gKKlaStAbbhBb6Rmtbs2WVQVLS0UToP+zRUSmr6R48TKFB/
KtkHlzFCPTQZ0m+hJjszT/hwoiO7I7/SfLmqhlHf6uWM1Enj/HhZNC9m9/Thake1KLMYVEdpoYtw
8go0/ydTQ7pA5AQKOs5bzRpINAFVbp2Lu1Lhri0GYxZcxX85E7u9ByiSUkH83GucOWRrvAUrfpn8
Z3uYGkEhlfNNjYM1u04tV7B9iLIm6WGOBzQ5Yd8Uvn+ffOmkKVlnbIrS2+F5kMDlENEpdealnuam
iflq4poAuc8KkARXas9FO1RNepFQcENf0z/SQeft+ZfSSxj87qty5yLcB8fXt3CT/ygUuP02paRs
mCnOZy6YvsrghsCVmnpCzgPT5qjcecTyl+Nm4JgkXk8G8sKIsYawR6GoZwgXvMEauMCRtLa/DTk1
sb8XDusmHSQ/+w3J0TtR5QsezzdolA4sUpvqrlTnV0ARHmA+7+DmPXyo63s1+biJnL8NwdufK1mt
VGR/0jzMDWaPwTczputiI9npjwptojcYB4HbxD7OcrfjrqehU7HCb5jnP7AIzeJ+o8JCxU3jFjIB
SbeteZP6FEwpP1JLsUP5eOyrYIAMCo6nHrreAL0XXnRISB4TOdboo35OTdC7B0E3JUYcOMKFGBzn
yOR+XplaPgp3Prmiw6IpwKhcQ63th+GyjRF6uPJyuRN3RnlkwETN/5zG2P1qO6AuEpSbELPkHjOg
cehwtBRMvERGxuvrtFk46GVWOpuZ+khORmPMlShbaa22eM+N2HLyJ5lqFfFe1Kd+l+9Hd3TWihah
fzZChTvJ0p98AafCeKpH/DXIX51ttbt3NQdXHDrcU2QGftYTCex/5h6F0y4G6LXxqyO5RcmR79z0
x7Y+uEoNi+kmTlH3z9Am2oWvP1H2LNwZDJM/jwI7GxbDJwjgzQwSDAPP+1QMJh9npJqRWI6NnnCZ
1CL12qfHBcYmUH0IjtigG8+PEJWNJIW7VFufUzW2SP5JHFpDZajwBSKselQXcwiSPuACOWX3aScZ
/qdmY42sYxf/3keshf6ErHWJhhe5CiGpENzitPRhaWWACAbodM3qCczTF/Ldjbe1BtmJL5ZHQytc
mzvT/rBq9mK5VkcBri25SdyCvXTyHEeFnS6dG8ZXRdQIvqcOXnTb5xgrTYab7jTfYLw2hoTG7zWv
jAkQZR7xYpijasIQViHsCLoe2GbeYwMkWwY/laWpkUt757OdPxdGzGrpc24/yr3nODawLDWvhMmp
DbuH+hvFdUkAXbm+jOIshA98AHs5KHyvvy7yLFx+tMaB2Vn3Oj/iLg7tmhfSsNhc4eS0utEv20av
dXtr7SQdKyzN5qi73fXkZphRbj2vIBM5p9TB8lRNM5X/0nkhlX2TUq2PUAbDhViGyhud946Fzeiq
pxDdaJlQIQG23gjbHp0/PqPPCswbygmWWtJDM7/VHAcq5QY1Ve+EPT4Y6DvYttPMl6on2OHsJhaW
pBBaStVF0C7bZ44GE6Dp/Wh8+CnJ4nbLfx945w9XhI0YE6SRt243U95iBsA49wVP+RrAtGKdg1gb
1czyC0Q+VoG7OhZnXZi9zQSr4x/JjCCS/wswM49ikgJtrcb0yklIUjLK2Ljm3IHR7TZ9G03/f61l
M0EvY5mfmFYDD5xfW/BquNBq+RNPARk1f87NHxAhe19qHMQf/sJDOI9kVCcHHxGys6qndDjGTR5A
EEiN0S5dT+TrV+NutTUAyayJq0qVBK84cZxH+P7r9B3MWjIwDnuwQT7CG8t3akvMpEQv3udWSHzX
njtda3MJCfczld+DR6oQCXeqYcFSPm/oOu/qKkQAHytqwKAqmHeNiN7xmHyME2YAb/8w1ZTZCMZG
dcV/JDlqyulLd//zefiMnZ1QhSDQc9Ob76Prb4C4PokBKf1HZt1A4YhVAl7jX74BaqbZoK76ItFJ
oX6UMXmatFXdps4ON+eqKT0S5WklNB9LRdpSDoRIS1NoPN7xUEa+BEFgyz+dV8AhSw/nM+efsluq
genjDC77FNhaEal4mak0ErMVKgJznucgEE6nmi5ByWJzettVrIT8dIOE/gy4hF8z6F5ahkyjyiXK
wymhEkkbDYcZYHYyTJeRPd7zmeZDQ/EV+2xQvDrrnwrygnmAvBezi6uS2CVFnK1ISvWZW5yMOTCm
rUEkDSJPc4ob093JuOuA32iFQfM7nz9KifmBa2oBRCFcm5UCv6OBkkee9vQ4SvQT10QQExkZYt+p
gEfmdZN+j0IYwQNsyaSLCu+OfyMzBTjX/Li51imLTJZ850GC13I4RXZnOLHp7fC1Wh7kV4hQjWWk
M0SRRglGf4iNPxX+kGTwNHwHjgFjG7ZW8os0b3Qzb7zuxgKeRcRpI3fVQww9gph43NVW2C1eD/yc
ubOAgp7lomxsMHqYeeyz3GmcRz5BQbkFgLtvDVWVlmq0relXwqNDTyCAx2c5cluBj3xe5ukn2SUY
Pyw86taaFF+1Ussfl+b60urQL13EgRLDX3ZJ4fSItatSql9D+ynrrmtpdjl6xXWx1615CXMdbL0A
rArnLl8EarhnOr4mP2jNdG+JZ4WkQViiEI17+L9wZrFPf5NL4GMK0CmQV1E9HjoS2Ym/yk54ZUVy
rFgi4hck2Fl2P8kBItUekIL5s4eSCtZOEQy6MS2Tn6zc8tNGHDcgAvKYtReqg5+dbK1rxvZ+vh62
qI0anDlZWyJQTvCOXF8/Bit//FU3THnUmgqzjmQ5kkngUJWr9R7Ukp/LZcR/2sfFfv90G/95NV2r
vqIH7KXy+4mPwDOdqdW2ooTzWUX3dB/VTT05Ensvs+/1K0kW0PpJI9zIraHccLmujVvkGkzeZ76+
v9Ywcp1sl0ddl61o26TewVwRmhTNERx0Pxuijv9arr1lpg+Uc/V1QFJQMOLFkJkBLDMOZWRydHIn
awRZhmjViw2D5Vsq2J3jWbaMGAiQEbAyUsqopz+irLWVK30BXQH41dnWUrV2i+c/6qZvXh69rrUT
WNtEsejkEeoIa7sAE8vElc8+XcxEP9IiNPXdMJrbplD5WL479YLfjsEPuoImT5SARzG3wtdJpZwc
OHbJI587PFs5YYeMvd32s1suScVNLTIAtkP2RfdHEd+Vcxp0dyiG+O5di+KixbN8dV/q4M+OVQHZ
rqB7lnh5RqFwCxGtq+3Xn/rUhmrGKLzvie3V3DwPEDAN3X8OHflC4nVHu5zdi81LeX6+kZBdzMFU
V/2MAKo78Fi7O3UUuyBX/39O938oTC85L0yQuxxHfj06MPZvRXuAIVTSYPHfBNNUMKIwTvt70LLv
hZSgvJ6OL28avqKx34p3KotAPsRdw1V1ufnpIBVdH/4JcwmwlcUcQoBYF3B6PKT8H5662IjjPqYm
WwUgZFt6zpe3fEdCdTLVBq2MUVUqpkN0SskR4I/OMLsVpzAsJLttaFzHBZNk6gbTpB2F/a79lnlx
wtPfLaQTgrkIQjUSYvhvMokLEjiZqL1QqbvbnIoAreW5YMk6PZtLeOWuXtrAAIAPEZAOQL0KwyKx
TlFMQVVGab9SdunEwnb3PGk3oOcy79fHSvvoVfNODnBTz0NEzGuILV37WMXCXGH7JC2MJl7fTGiO
IdnUo6YdS5XtQT3cJqvAgJmj9WJGCsD3StpybxtP6na8D9pKCqCUF1APwmT9A6dKkAdVEitir9yl
Sb5aZ4XrDy9qYGCTI0KgnkC5+n5NFNx6nk4wkxizRwvaf6tM8j98KX8QyNQKz92Mvc4BP4FetMsv
5xUXpPhLGnzPUg7BSPdeUYxr/GYTPjPiMJdofkbjGi6di93w3ylYCR+oHghSP+jHOQUu4NFHwxzs
SRHi7Mjte4KqTyTZGnFGSBQyhv6VFLOzNXIkOS13p7J96NcvGXOngty6BFwkDcDzQcRDzLQPWQa9
hehdQQpnLceJrG4v6unR7OOGYIExySjFe3qRKQ4teoKGwiQpRE5o0XC4pjsz4zPN7SkKLJCi6YDg
45dU2BWJbDcgGsP+yWzc4h09tfg1XDIkjacxUDsDfpTNVvcKcsA0Df+5Q2BgbSZLweuKv8fCf9gx
vOYWUYtyVOtiZFB0wtgC1YJaRBgxz24/ZZDcxPcdFRQaEiYmAmaEK59yihCUTJDvUeL701Bs7sK9
bQigPQM66aUVkp8eErH9J82Y1hBc0hofO2w8jbqXWKg2hF6KMhavqogwM93lUkjDpt7IPaa7Lyd3
Z10LvU6o9nlwpQbPeIXCJAOjhJFjmKygN6MJ2PVl63BdKv2fqx2xG6ZZPgnJ3u149ULa2J9+TvWS
L3sY4VJIZzCpGN90NN42kzqOzrpBuMfTn6FroHN1/5dbA1Rg83vmIuGo01jPd7AQWFJvSwkjsjUZ
QW7eoy0iRdcIGETuC0kg8gPzEwtnzKg7l+xsqm/26fKyb2c5jiyXH8l7TgHctLPXWn3mexeVRbpB
pOjbA5FwzaVGw1zyqLtstZH4785B9O9d884gZ2GHl5ii7KTlAXR1f7zHsm3xwGtY5eybBMiz5/zz
VxHK/Jrg+ZgXRSDb3jSgbEjmTiWqVC/kAXRW2Kr62URUZ3cEUwqJDYP4TIrnVwW53WADzfqpKLi9
Idg4CXLduTOffnGaLt79kJSsgZZUeIb+mCGN95oJMY5YiZ4KtIGy+wuPPvW5qSmSx82vYimy2c4E
JkZOcLeHeaf7qofikTWSkyGm9HQrSjmhwOvBb69EILRMTGgn1LXyNlZudoN4A+b1HRkq25eJzn99
fvK1Q557LjwgZsih/A4GIo831M90TwtNq+hRyhgc6ebkxzu0utfn24+I689lawt5gHOgu0bVOxJG
2kjsSJDD36mrakAyadggTQ+f3YSYA/6wf3o6/yQA/aB6LiHh7o33HazSHzP1g2cjNBNOOt35XFeA
JsQSkh8wLmhbM9nReAqOucGeizPUrgmZxfeIIakjaFgeJ45KROtSBHXPZDgqjzJZjQRM1Hv+NTKE
fbn35UOX9L7xnW4vFiJWyGbJ1MTgxs4L7pr5VKUrqx8K/HZ0s0Ef9q6h2vVH33HiCtAdt1aTqJXu
HFXzXhPeoMo5b3vA05Z2p2WRb2KRxojlDYxchWilLPekv4Lm26ZA41q3YJJ7ih+5gMWNPa/EvMjt
02oXhzP+JCswWkMu/AV5VYa+C8f4l6aro/uT0XTF3Y3kMspYOq2O1aFarOhlvdJKwCtLRJ3xeEb4
0D6tY4EovB91UNyFJX5+aVrSHzetNVxcd6MBI6t9ZaBIJVRRCe+YBAKb5J7PNgNilg7NQAtbyhOJ
ZVM37c/HqvjCMdB6k/tDz/LkExyproKIPSoelWjZZtwaVuCbKEQpIMKeth4TgLnpDPHmT4E0wfjK
MYnyinFslpoCNrYTGUSN0glmn2R6dj7vq23zN4Cm7Wcc+8X5IlIhQ3Vc0fgjQ60/WkjLYKVWAbJt
k67hGg6OxLL/0JD1dx76G0pMEJfO3GT/IoHUZ2r+5Eq2lA0gClwu9LafhhpoDrTgk+rGeEcixf8L
1X9VT4ntb0HbIgwYLUo7j4zj9fNZIalrt+WdDidVFaw/4WB9IUK62X1k6DxljQkywALmu5Mnm9Hk
TlWp2v/wc6GBwavoLnnm/2tUTLeAajM9Zwu5zQUdqDqFECapy98xsFniv7HY21pHdKL/lb0pE5CU
FFQrCWQWYbzMKmY515zwfpPgDHiUItngsSURxdXqoQxK//oCpyJxKFhNHujXNQ8KptjKVNDxygQp
+IE9NoiED8SyRAzyYAF3J+oeKV1rzH2O6r0G5NiPzTd9J3Ofoke8HGDHyX7biXEbpMdvp+b/zF7+
oaDtB17YUOHot3JBi4CGZG7zeelToP/f+YjNb87kONFisXHrU3VHGiKCbblqeEeMTGy4zuZ9u1Yp
6kEBRYhcQKEUR6ndzd+hL2Bp30OOjuY8qQYhi+WpnUXjzuNdE336l523IcoibBOIodXlhCoGJN1T
gDhhS//u4OPig3H9MwxWt7ze73Z5Of98cUg9t340X51KQ2uwG81rpT/kO5oQMgANu6nrIKpzBsbz
m3WZ5xXgaDd1byIGUzBEBkcxl8z9/2PD1+giWFcvCcFh9vgkIMICqDlIOm1Vbn0B/SDP6yAp5r7D
pRpq2hYKNypdcQdY/DM2d3sS+Nkq2gbmHkb5MfrRP9sCnT/ztOsIaLf89xtB9BoUoz7Jxi2yO+Jk
ML8ucywFJV3N6j+ifTDLlbcaJB6BnZySgdUUav4o5Bt2oKjUb22RAMhqJzFgva5JzIJFa6ceMiQ2
A717yX8wGWLaFAKg+fLhM+nt5pmsLjFOIyMkRVgGDmZQKoFSQMGkCa+u+/Jkq6Io4oZJSSH9vnA7
w0xnNISgFV6oLWDrvcKa49DvM8q1hqZcI59QVjLODFCkQvK5nEEJn2JSZahR/N7dglfIfI90MVd8
DCJ/EU2KVN4DceqCr9gt55Y1XywEBdT1287IpjctYRKDo5Fgjg1Kl3s6u+Gj3AGAB6hU4YGrtyFT
HoWFCt8YZMvTkBvdlKrPU08cMxao4V0D6YnJP91GTifRPok+9+elt1h1M4WFOv2KgnwPt2IN1Tjp
qLJU6KOz8lO6i5S0SzkvnMaj9r8fsC/cKH7alV5ZOiALPX//HEEsntHquvvDiPEmvzlS92LAMjsN
5Yk3/W38Fpj1IjNPmSWPjkk4Se7GBJsooot4h4t+N/xNSTEYWtC5U5lCprVcbrmfuRM7JISbRjOx
7EgR5OaRN4vcSJhqLNP2R0T8GnFIrvgyOD17n6gNvykywHx+EQR75mua19v5Xld+WX2P619zMOai
HEN5m/7u9mLvD2fX2W4RZlaNYRlCM+MG9y115G+9iBWu5r3z7D9bv4JBfUEw8LS7wIy1wEORYbOU
12AiNM8Fwla/5mQv92pXPgBqGfCz9OHLURnaYfS0SDIVHCxj4P6bzUEwSLjkHMKSPU+sHp3tgBRa
zSv0RpV6NSbwmKRkyiuJU39V41u2azMSB14IMNEB1Z9zVoyBOD7WzLJ3Ft9ZYzhM/aS2gyJP8tkM
u1YLTfTn5OyrYjB4+enTdRqZ6neSZQ/FcpZua2VF4J+GB+XBuU+A3zISrGg9sHlYuDaaNlJAP/yM
52Cg5+PUHwW5eXA9LXO+0taJXab4Aq3Hskm6Qs1dDv2v++gphw1Q0NVPaU5/O/3JeSb2DGvYNiqH
HGNiZ5p3iumpCbcgMkpcU6ZUEcspY9cg1kr8PdaRCD5rtWwn6gk0yFDK467aFW9zKJoovfZjLNke
gJybLru0HnZldq4HxSQ7VtTfONBYixqXNMEhLLO6HFvvLwA8xn3jKb6GDvFaWLKCp9hwUmlI9JPD
FBUhIOmZOUE80Dphv+BcfvxauC7feeDFuNWpse/GVNc6/Hx9wR7/7O4wwtK993zi+qUomXsgI7Na
CW6dbOPpgPrSbbxe42+9XUNKJimmIDP3Hprzx+IqBqrIpWisiewrnnoXaim9uTJ4EhJxenxiCYXv
UKm0vu8YxA31DkK1psNsmN/iVaPU5gqmVF1x7ZXh28eiWpX+YFNY4KTaxOLtvzOCXKO+rb/7zAo4
9FJnGctkthEW6Ge3FvYKYg5PfXdBwwTtC5Fo5Dp1UMYvRUsy2u8d72j2BA8m6FVfoVPyfYXhL/UD
Cvir2Ykr0iy+tkQbjBrgL4j8wZg+GJ8/YTA8/zIr+7MOVUBAnTZkxn6mkLQLxQ8EjUPtf/BNey1j
AjACnsA76pPK4kUvvHG/8sxOnePsSDXl1n+utsb2cbahj/nLCsygDNQw13dxUZEM22GQoFwIpoY6
3hI/Hp8qqjey3p0PuvcDXO+q2TD8M2VIZ4tU4gY1cnt5HZ2/UUiTY3dPJvHaHPkGJeIu7V8X/Ya/
+RWhZhKwYdP5+Xh4vnvOXH20ZY8c/rydS+cRS+yF1He8iz8mt0yxymQVKP/7scf8iSUlGoyiE17B
QLO9F+s8Jm1lbHtHJ0MaXXUstnG6KJp3nXWv8kKaS3rZUjDtQ8FPVpY+DF8a1GaBFgRKkvpd2jlm
fXuOXNJmXV8m50vOJi/cLA77AXe/lQJ/zSIQijnuNYv0pn40aVvWTsRLugUzoAEE/pFX2ThIOR5Y
rX4I9NPmtOWfKARIKIjPQCpIGBihhhP9+1Qw3R8FgAft1Y+zz88ww9PInf/YHe/hTz6V57aROyrS
VjOUgEVPEI7Z/EEA810BjbQlanHzUpYAvaZKkB3ttYY2i7jdODFnOVbdfwS3KV32XGW1j4u/Vqmr
PiP/rhIly7pvg7LVGVx32jLA5B0RTnipDkT5vxd/EJ9Vu68CG7V6SVZ9b8ODlAu5JHeU0ARVZlKZ
Tk7oVg6XglW/LQlABJBS/N1XkyFPXHNsP7bQv8CjCUDRfiMY8RQOonY83UklHto0vBJ+xCsIvHuN
WNOz6oGoRXS1m7Y+fxCnS7qDuXHZcWUorLcv2fULQ3vkXcfyVieRnqmTABXllB5q3xkdAIFPFnd5
jvy1rK5kAc8E2lxj3aJbkIrLQ+7Gy3N0+JJWZQ7eTYzBEn/SqNZDoSEQAp4c9kTX1O2JcUA3YoAe
cwI2tVCsqqc56Y+yuglZ6dNDY1zPh01PxS5IPJmG61CyuR7PEN0x1hpQhDIhiJJ9CxzEN/fD3VwO
3YqtYqdEJYqUGZkupPsUJLX81naXJ8xDBWKTyd89gccnrnIuy5vkDeRrI44lnuSe8C7LdqhO/uYq
R7L+M00l67LdAn3EXqQ1++t7qX8Q6FiUPWgj94UrAWR6Cn2ykcyg3BoW5IPr39AOlvKipjTx7Mbv
fr5lkAkGpT1LIjqwqfnFGG+hWbfa99kjCBQb6h+dK4UNrTgumejp8WxPSTn3wnth5c5UfxUHDJnD
BjmQoDWMDLhn0rf9EmKuHYKICTcK8swtHp2D+jgE6tW5ZOGFX6EzuPeIjHZmd2IaCkvJC70KsNq8
mKbZloZ8SMoP0OEXMbMnr9mt/35UDxGgwfhIywtcj3PQrqljA9f/2WcpcGxRokewNZIOmepUSPcv
i1AzELbJy4PpOkkprGUXXpKeE/QXDuDBqbd0n0ahX++vPzLCNnKk3qoiAlEnmk39TnPZiVYUTBpS
abaOXWDr5nVHnOHh4M2ZWHdlndzGXu8niJ2nwcqorNLsAWYbIi9Jte/PVuW10B6y5idaQiJzg4ss
Fx2m3P7V6oAmZ3Pn6eMUk3Rgd62qRFz7jq294HWyTEAjjQPRR85kM3sS0lLVsFooz+nW1YQCTXNq
jZCu5gqT2Ole+LBGKPmzX2tFy4s+HSU2zSn+WDFbjU64OyF/oZzLURsC0dJ45hv3ITINnLadou7n
uduU+wfPRBzbnpPs2LcTAAXHelhohlCEMIGEkEC7910r7w1ZOlzsTBHCA2I0zPBn51UI8Dt/IXSI
TCR/h58irry/oY+vzEl07AWI0DERqOdqzwQaRQdIJEtKu5MtB/x2iYysZhdtl92YnvTkEeXjs3N6
cs1d6QArqAfBBxFnCKJHgQKYVW+6OpoRNUN2YgLtX5Ug6uQq2ySzLZIbOIwHwkVPCR78hKyXF5cg
RylgD0Xo9pQqWTfHqpRQ5y2eEx7EDFCE5gqYMYmczCKFyVd/8YdPZoGD+BZOOpHiLDHu6L9ytrtF
O5qd351SZYpq04fd4nynJ1TMYe3OkTEvyG65J9Ra+cgw/ME+06JgDMxUCX1EpJktHKANDeomTfTW
xTkYTnz2X6e/IF+9dvgkqVGiudnOopMse/Dpk4Uouw94aO11RzNv5ddxcw1uSKELA+0rMIOCscWp
IG1vKPDQTNS/dtY84tyDmwv25r8n5bmL4xkZ1OUH5MNB+Ct7CdLy/oqxp2eUtz6tnvVUCpqVLXWe
Qfy4DAqV5fimO2T5t1afroQ/9ZAzpFMx7UPn8vxThDM6JWnNHHZLpeqYnRH3XJ4i/F7oOScwiCgh
ncaD+S6wS813tLoTd/k8Lrjgo3hi/EUxFroBxqG6SILS9T++rIa3Czo/qa29cg0286LsT6nxycQ3
KnxQ5cCd9tDTv85/DbeTQ8sqJclyro/bhbV3gmrehQ7EhHrm0uo4VZXG3/LlXzmXI278waoQJ9So
MXbxl9izF99zMaIIwpkOyYM0N4w49IrXxtHLqQ3Axdh4b4fp0SJPHQ1M6fOpiZrUXqFFD4ocHw7n
DYQCh+N9q2dXbwRHVoU7qqGeJqqjiYeYdXyaja7kzrdlGOq5geS6CLmh14XNnpQDFBFAQJGkys+E
Y+NN54wiAZ5jr+5iG5yybCzzFYneu/4swuGLbernh4bDVdvLQNYHwRAfzsqxo4HBlKnqFMXmH2PJ
giBnmB7ypal3sAdBpxkf8Vl4gnxe+zbDzq4oOmqWCoVG+CLZ9RvBn/k2ke/cQyn/Md5tpDlQwxuY
iTphLUJ/dlPwjwhkTtysZXnyo3CJB0TbTA20bvGgfRfTtsSufbfoG7oZS27joop30vBzj20Rb+yJ
SWzoYbW9bAJdC9TijS9zekKltWyQn4FWvBx6lppzBSdyTCft5UZwKVyTs2zwMya6lSAsrMx3O3gb
ynYifFkiR42fZOJJnE54OK317PSbdnxceBoCZxhJ2Evv3Vy4R1/QGq8Wr1FcjTY4vttBOcMsTX2A
Sq5SPSaY/HyqJmsreqVsIl1R1LwOAW/KpuBx2gWkbnx/4Xj28dejciPaRT9DzCjxGxTXNi8ulCkK
Nm33wEn/EEgB8Mp5mYFu1MFZUHZQoe6QyTtiURVQBbioOKKHpTGl2CYcsw2EavZgyruFt9S5Mpnq
0lLZxgGkvNSBDD9QbkCAAdoSXg7WKWh2XjsKxeWY3ZzKjgNTrAI9uOxI4bDtsoX23S84JoUFtnJk
L0q68GahOoOC4UXtdzcXEk5yNeJXU7XBy15lJF36/bLIhcntgWiwXudZxJ6zCuAEfY5aeP9ron+J
SnFHfVJ/x/TXsDuQt0TiMb6eyY3nAPyCE2oZVciMUIkYNNXkPEpq2YFjCCM28l7Z6IaQ0loIQzB5
8zefhEtRX33F/QzlohKlc373ZiZnSdtokyK2U8QfMGNdMbfCxkvxvH3B+iZhepjFAmvIEijUc2Qq
TwnxMwOp3BNe45JJrKwkoUaFT08EyDOROTTmosQc5UfIOEyIzYtLKF5i8ywCYWUb9edRX4U1TnKD
CKkJ/i6GNnD6wL5Uk1COeQhuN5OFe7aBI30QtcSnIFcjSPTTWPV2yCWvw2ycD8SfBar7FkYtl/zr
cA08yDFRks2z3Hyi0o/otRVxbEFyOY6NIQGzFp6njV3kxoHpUNyOxC0a9nLd/yG6o9HUCSZZAaVK
2DlqyNWztoxWmFwJIteNoJ4vRBYULndfk4mpJ5fAduH1gkaFXAuRlZ2KRFcH1WrTl2sCI/pn6qGh
NH25lklzKl+ACI1RgFQsNX+CVYNUTnarjl6iPAOEBXCyLUSzmv+BubAaS7dXX3JMQpIUj7nEOwUx
SRBDa3qrTp0pASF7zVzg9PgvXe5OVH48sD8OASme/+pA/kd0nKdGOS26IQHsm+cwloSw73l3jzWJ
25x7iby5rtxXXv4rzK95/gyxbX8856f94yWakTctFpZzEB99YMGijyacw7GHXkIwbzEb8+wHpqFT
6GjVqNKIUKWm+FM+hIGGpupYahF5Qz9V0+dIaGEvHmWxA2XiBPYHcoPwpEE555Ml7E7eLGDbV6AU
Jj/bt7tHS/42/YcVD+fXxTtdnuHj+HSOhZuKBYx8AkxvMhxycO/vyFsKOg8gxi8oyz5Jf7VxTTdV
+IMT13PqfzP7XpvmNr1Btjk3O5HJL12hFen8OPO5iPm8x80qcRHx/Erw/Ne3pgGxBUu/h5vjyMeM
dl2Jano39ZM+eKQPtKRq5qE6aYzGZ3oHiFJPTbJv/39tXzh95PiWwxEV/EdgdKhynbOG4KDGGb5t
J6tqO7f/BByiptDFp/CVOQGNneRp9EuSbBBn7FpEDdZ073kW4p9/xQ8iKMKJwNd5UapXGoOO5SVg
OTtMAMXeIqtBKZmARf/yFrjwbXgbYEOK91NKLMbeGQTWDpAAV/W1K2DQKRuWo9M7cR7QLXAjOY1f
Z7ZfKSZ8MT0EZPqqkje8zVlfmbNmDKaKcZQSnRyLMltkskE3oOb1P3vGPue/a/yle1zVq5CbWtAl
gjBn0vhLdSGvErEQjz1HAH7Li1dONxz1epPW2UcJv2uun0GUDbn7nKuc8yB6lqb/1T7ICZRCOoYy
RbWUgBOdCgczCapEOVSw5iRgkPIMB2HK8WAY69tb3CJO7h57ekx71CoXH9Bz9ElHF/yjxn19XeoK
7O/0y1sDDsy4MV/kLVh5+ycAcfpZ1/Op6OkAPGAaVVSaUbVBKdpb8LnQEVCH1W/s7Cw+065GNE0A
HxYeIH9zToqmdbGbRSngNkcI6yHSi58TGsgEEP3BzcIOwhWzV0loyaTqPe5zucpxkP+do2U1uJYo
ulnSackUjZGhRDGScoUJIGYhJX/ZwoImvOLu7xR+veODQ4+MuJv/H6chfOZQHaB+crzMSIaagsOk
04BnXUY0Sizk6RboqgfhBbOpQkK9QCCdDRrgfCA7b9nNRNuA4mBHJpZJjk9q3e98O+ru4eYVd2SI
F/nJsgntcF1bgPT+JX8nZ8K5O0z5xA2Hlo/i/Y2kRUNbZvni0IMk3y1hpf3pH1vZ8vRFT8PYLx7n
8EK0e/tJ6DI1Rsc6Fq6yNd0Oyz1qNHlva/y57uDyS3OH1tbJngiTt5Gt8hpWQEQLM+l5Zlzfscal
7fOlyCl5FR8WRqxks7oobzDM7v21Wg2IQZZQkI9wjElR2jvDYGCJktm7lzO/4/W2fkDwJ4m2kZrd
5c25hiHEE+Kpf4RJoQAdmncuEfcK60NMTlaNBy/7fB71nEP+JTNKoewd6/sRJnYpB10ULV7V0Fxq
9alYYITKh2OwYmzf/47KNr6h9tYj5By+uhZz5thMywO4GlSNyOOsiA5ZaTzgnGDODB3Azkam6pM5
aX3JHpyYwerEqyp55QNBq1K1cZqElykp66POhkN06LtP5Xdm2w9OEBo1QMCJq+FhgM9//r29yLDo
V83kzJiXsm+zAMqL7/erRlvnpQQ0To/QNqbgFbogn7oiHiP71g96CISorYAestDS51ysGY6CYB4P
qRz3GEBQh9Tgo45cZ4sOuHPHlPz/0OGqhXRAQ+9a6gS1lgN9DTkBTi9I3uAoaRozkoUsF0A3T5AN
SXUS644in84/bnxLrEdKpLylXPZd7jCj2YrSrhXtp0U67r+KoY02zpfTozBUnMeiRsh/4779YXrL
IPxZECzxZVtG9JD5MYDlqqkDEf7uBZnqxFfdrY2LlrzwCVRPPjAN1boWaRdq9r7EJ0Pvx+Ctv1uO
ZqphMCRD9xsBkTWApWbppBPBmCyLdooa8L1PhQGBWkMn1YaGr9VjKJ7Bl/Q67fB3Azx9VEkf8E2T
3uGmFliqEjryWEGqNFY0Pn/tvy5wcHS9MItL7hmiZtW5wFLTJBfxZUyGK+kw4Z/Gm0MS/WtTqwHH
7NpdmV4zTzC0rU4fTAvMJPvT57N6wH69C4INhZ5Lwm58HIc08iyYNf/Mol/Tm8mrsAoHWh17bc9p
Gfa3y+VHBvSvmLLHfiwNzn63d1h7U1NozWWD6DrWOAxdaiVqsEIj3o1LND9fI4zkeFnaZa9th7US
BIcAAUbGPgE+Y949w2x0JyL0hybcddjaXvexUacKW5G3Hx/iVP4NfOrNH569rMGh3R4Bw+1UqSdS
rcLFan4+B3zJU9XtLAaqBEuWQJJugfvSiCg+fEVnOPE3fCr0IBsgc69u/xo+yvnBXi6aMelIdx1Q
1ynKnekhxheCi0iGA3fLW49RXd0qo2m/jwdvfPQSwfG9p1mTvErMROlhzClz0Q0nhvuFOFssBGO+
IW+5WFsGC3LMzgeag/312vyqrQ34RXgrjAOHRZu0ohSt9GH2jlSgpFk1nwHFQXJQOPL4IQ4hmGRc
J3zv+PrLVtwlAjQ+A3Y2crHZLgKS0LX273dLv3EQXNaiccQo4I/KVfelbvdRGY+x186BRiBvUmIj
o0U/L5gD+XxJbhuiPK2ugcIR329eKWYkLpN57QCSRJcemTudI/ClvUtMM/xmaVAL3PmlAOxe7bbW
2gRslqgLWgpTbkGHHKD/AP/E5fpF3v8h8+oIccVa3kuzEXVD+87oLBV1udHODU9QIaNvn48ffikn
wqwZjkM3loMDGjRbTtJ5RtmfsasdxTsanvs2g4e3CoQ5vhwEwB0lGeZyg1dzSU0SOcBH3iDyA8gF
y0oAl01I5egiUNUkvWCYKwHj5s8CkXUD9rMlhKoQnXNQW8KJG3r3i2EXV367k9xvL118nZDwyIxK
Rc3TGpuy5uxFAXwvi51c8fUYKLmI3IxajitDx1/g5LhIPes6ZqHHbemSNuDy6XnvLxuny8jF8tPr
Zlz4FjErEh3qQvdcXUAwQLmnbB42kThQUZzWI9L8WYLMfDmlU51Au0IpIj/QcxanmTaJ0jHeBqnS
DlmbJqMGUkXwEME4sFfkW6vufaQ1uTA7l4sFbxVj7jxymWYp5x57b553slqwUGTZ3tmeOMm3ZrTA
7FmREFJMjxImQpzphZYjJmV88dLqK0BSUnIGCbUp1M07KnzRXPUu2DaJynkZH4AAnYyeZ3jsvYGp
N/XAz1UpHSbVQHEBtzj7ghSFoOkpurtuft2Ry2kjG/Wo7g9dZVud+OXqrJhrvfBPVb+6HsuFMgfP
pSLflbnRNsHX4fDIdJ7gzf8WVFFcBVRW3mGEJvn2KR1DxlWy0lnBeLtFlLbFeHX+YungJLd2UZPJ
GwWg3/bVflpqzWC5YkbxVp6n5i/Vlh5faGIxNv30NbuHMTjL6JU3lpgAQDeaX1tWSA1Cm6sQnMhw
wQQW2USKrA5Amg==
`protect end_protected
